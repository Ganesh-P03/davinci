module ROM (                    //Instruction Memory
    input [16:0] addr,
    input clock,
    output [31:0] Inst
    );
    wire [14:0] address;
    
    (* ram_style="block" *)
    reg [31:0] ROM[32767:0];

    initial
        begin
            //$readmemb("inst.mem", ROM, 0, 3);
ROM[0] <= 32'b00000000000000000010011100110111;
ROM[1] <= 32'b01011000000001110000011100010011;
ROM[2] <= 32'b00000000000000100010011010110111;
ROM[3] <= 32'b01011000000001101000011010010011;
ROM[4] <= 32'b00010000000001101000000100010011;
ROM[5] <= 32'b00000000000000010000000110010011;
ROM[6] <= 32'b00000000000001101000011000010011;
ROM[7] <= 32'b00000000000000010010000000100011;
ROM[8] <= 32'b00000000010000010000000100010011;
ROM[9] <= 32'b00000000101000000000001110010011;
ROM[10] <= 32'b00000000011100010010000000100011;
ROM[11] <= 32'b00000000010000010000000100010011;
ROM[12] <= 32'b00000000000000000000001110110111;
ROM[13] <= 32'b00000111110000111000001110010011;
ROM[14] <= 32'b00000000111000111000001110110011;
ROM[15] <= 32'b00000000011100010010000000100011;
ROM[16] <= 32'b00000000010000010000000100010011;
ROM[17] <= 32'b00000000001100010010000000100011;
ROM[18] <= 32'b00000000010000010000000100010011;
ROM[19] <= 32'b00000000010000010010000000100011;
ROM[20] <= 32'b00000000010000010000000100010011;
ROM[21] <= 32'b00000000010100010010000000100011;
ROM[22] <= 32'b00000000010000010000000100010011;
ROM[23] <= 32'b00000000011000010010000000100011;
ROM[24] <= 32'b00000000010000010000000100010011;
ROM[25] <= 32'b00000001010000000000001110010011;
ROM[26] <= 32'b00000000010000111000001110010011;
ROM[27] <= 32'b01000000011100010000001110110011;
ROM[28] <= 32'b00000000011100000000001000110011;
ROM[29] <= 32'b00000000001000000000000110110011;
ROM[30] <= 32'b00000001010000000000000011101111;
ROM[31] <= 32'b11111111110000010000000100010011;
ROM[32] <= 32'b00000000000000010010001110000011;
ROM[33] <= 32'b00000000011100011010000000100011;
ROM[34] <= 32'b00010011010000000000000011101111;
ROM[35] <= 32'b00000000000000010010000000100011;
ROM[36] <= 32'b00000000010000010000000100010011;
ROM[37] <= 32'b00000000000000010010000000100011;
ROM[38] <= 32'b00000000010000010000000100010011;
ROM[39] <= 32'b00000000000000010010000000100011;
ROM[40] <= 32'b00000000010000010000000100010011;
ROM[41] <= 32'b00000000000000000000001110010011;
ROM[42] <= 32'b00000000011100010010000000100011;
ROM[43] <= 32'b00000000010000010000000100010011;
ROM[44] <= 32'b11111111110000010000000100010011;
ROM[45] <= 32'b00000000000000010010001110000011;
ROM[46] <= 32'b00000000011100011010010000100011;
ROM[47] <= 32'b00000000000100000000001110010011;
ROM[48] <= 32'b00000000011100010010000000100011;
ROM[49] <= 32'b00000000010000010000000100010011;
ROM[50] <= 32'b11111111110000010000000100010011;
ROM[51] <= 32'b00000000000000010010001110000011;
ROM[52] <= 32'b00000000011100011010000000100011;
ROM[53] <= 32'b00000000100000011010001110000011;
ROM[54] <= 32'b00000000011100010010000000100011;
ROM[55] <= 32'b00000000010000010000000100010011;
ROM[56] <= 32'b00000000000000100010001110000011;
ROM[57] <= 32'b00000000011100010010000000100011;
ROM[58] <= 32'b00000000010000010000000100010011;
ROM[59] <= 32'b11111111110000010000000100010011;
ROM[60] <= 32'b00000000000000010010001110000011;
ROM[61] <= 32'b11111111110000010000000100010011;
ROM[62] <= 32'b00000000000000010010010000000011;
ROM[63] <= 32'b00000000100000111010001110110011;
ROM[64] <= 32'b00000000011100010010000000100011;
ROM[65] <= 32'b00000000010000010000000100010011;
ROM[66] <= 32'b11111111110000010000000100010011;
ROM[67] <= 32'b00000000000000010010001110000011;
ROM[68] <= 32'b01000000011100000000001110110011;
ROM[69] <= 32'b11111111111100111000001110010011;
ROM[70] <= 32'b00000000011100010010000000100011;
ROM[71] <= 32'b00000000010000010000000100010011;
ROM[72] <= 32'b11111111110000010000000100010011;
ROM[73] <= 32'b00000000000000010010001110000011;
ROM[74] <= 32'b00000000000000111000101001100011;
ROM[75] <= 32'b00000000000000000000001110110111;
ROM[76] <= 32'b00011000000000111000001110010011;
ROM[77] <= 32'b00000000111000111000001110110011;
ROM[78] <= 32'b00000000000000111000000011100111;
ROM[79] <= 32'b00000000000000011010001110000011;
ROM[80] <= 32'b00000000011100010010000000100011;
ROM[81] <= 32'b00000000010000010000000100010011;
ROM[82] <= 32'b00000000000100000000001110010011;
ROM[83] <= 32'b00000000011100010010000000100011;
ROM[84] <= 32'b00000000010000010000000100010011;
ROM[85] <= 32'b11111111110000010000000100010011;
ROM[86] <= 32'b00000000000000010010001110000011;
ROM[87] <= 32'b11111111110000010000000100010011;
ROM[88] <= 32'b00000000000000010010010000000011;
ROM[89] <= 32'b00000000100000111000001110110011;
ROM[90] <= 32'b00000000011100010010000000100011;
ROM[91] <= 32'b00000000010000010000000100010011;
ROM[92] <= 32'b11111111110000010000000100010011;
ROM[93] <= 32'b00000000000000010010001110000011;
ROM[94] <= 32'b00000000011100011010000000100011;
ROM[95] <= 32'b11110101100111111111000011101111;
ROM[96] <= 32'b00000000000000011010001110000011;
ROM[97] <= 32'b00000000011100010010000000100011;
ROM[98] <= 32'b00000000010000010000000100010011;
ROM[99] <= 32'b11111111110000010000000100010011;
ROM[100] <= 32'b00000000000000010010001110000011;
ROM[101] <= 32'b00000000011100100010000000100011;
ROM[102] <= 32'b00000000010000100000000100010011;
ROM[103] <= 32'b00000001010000000000001110010011;
ROM[104] <= 32'b01000000011100011000001110110011;
ROM[105] <= 32'b00000000000000111010000010000011;
ROM[106] <= 32'b00000000010000111010000110000011;
ROM[107] <= 32'b00000000100000111010001000000011;
ROM[108] <= 32'b00000000110000111010001010000011;
ROM[109] <= 32'b00000001000000111010001100000011;
ROM[110] <= 32'b00000000000000001000000011100111;
ROM[111] <= 32'b00000000000000111000000010010011;

        end
    assign address = addr[16:2];
    assign Inst = ROM[address];
        
endmodule


						
						

// module ROM ( //Instruction Memory
//     input [15:0] address,
//     input clock,
//     input IRWrite,
//     output reg [31:0] IR
//     );
    
//     (* ram_style="block" *)
//     reg [31:0] ROM[16383:0];

//     initial
//         begin
//             $readmemb("os.mem", ROM, 0, 16383);
//             IR <= 32'd15;
//         end
    
//     always @(posedge clock)
//         begin
//             if( IRWrite )
//                 IR <= ROM[address];
//         end
        
// endmodule

						
						


						
						
