module ROM (                    //Instruction Memory
    input [16:0] addr,
    input clock,
    output [31:0] Inst
    );
    wire [14:0] address;
    
    (* ram_style="block" *)
    reg [31:0] ROM[32767:0];

    initial
        begin
ROM[0] <= 32'b00000000000000000010011100110111;
ROM[1] <= 32'b01011000000001110000011100010011;
ROM[2] <= 32'b00000000000000100010011010110111;
ROM[3] <= 32'b01011000000001101000011010010011;
ROM[4] <= 32'b00000000000001101010011110100011;
ROM[5] <= 32'b00000000000001101010100000100011;
ROM[6] <= 32'b00000000000001101010100010100011;
ROM[7] <= 32'b00000000000001101010100100100011;
ROM[8] <= 32'b00000000000001101010100110100011;
ROM[9] <= 32'b00000000000001101010101000100011;
ROM[10] <= 32'b00000000000001101010101010100011;
ROM[11] <= 32'b00000000000001101010101100100011;
ROM[12] <= 32'b00000000000001101010101110100011;
ROM[13] <= 32'b00000000000001101010110000100011;
ROM[14] <= 32'b00000000000001101010110010100011;
ROM[15] <= 32'b00000000000001101010110100100011;
ROM[16] <= 32'b00000000000001101010110110100011;
ROM[17] <= 32'b00000000000001101010111000100011;
ROM[18] <= 32'b00000000000001101010111010100011;
ROM[19] <= 32'b00000000000001101010111100100011;
ROM[20] <= 32'b00000000000001101010111110100011;
ROM[21] <= 32'b00000010000001101010000000100011;
ROM[22] <= 32'b00000010000001101010000010100011;
ROM[23] <= 32'b00000010000001101010000100100011;
ROM[24] <= 32'b00000010000001101010000110100011;
ROM[25] <= 32'b00000010000001101010001000100011;
ROM[26] <= 32'b00000010000001101010001010100011;
ROM[27] <= 32'b00000010000001101010001100100011;
ROM[28] <= 32'b00000010000001101010001110100011;
ROM[29] <= 32'b00000010000001101010010000100011;
ROM[30] <= 32'b00000010000001101010010010100011;
ROM[31] <= 32'b00000010000001101010010100100011;
ROM[32] <= 32'b00000010000001101010010110100011;
ROM[33] <= 32'b00000010000001101010011000100011;
ROM[34] <= 32'b00000010000001101010011010100011;
ROM[35] <= 32'b00000010000001101010011100100011;
ROM[36] <= 32'b00000010000001101010011110100011;
ROM[37] <= 32'b00000010000001101010100000100011;
ROM[38] <= 32'b00000010000001101010100010100011;
ROM[39] <= 32'b00000010000001101010100100100011;
ROM[40] <= 32'b00000010000001101010100110100011;
ROM[41] <= 32'b00000010000001101010101000100011;
ROM[42] <= 32'b00000010000001101010101010100011;
ROM[43] <= 32'b00000010000001101010101100100011;
ROM[44] <= 32'b00000010000001101010101110100011;
ROM[45] <= 32'b00000010000001101010110000100011;
ROM[46] <= 32'b00000010000001101010110010100011;
ROM[47] <= 32'b00000010000001101010110100100011;
ROM[48] <= 32'b00000010000001101010110110100011;
ROM[49] <= 32'b00000010000001101010111000100011;
ROM[50] <= 32'b00000010000001101010111010100011;
ROM[51] <= 32'b00000010000001101010111100100011;
ROM[52] <= 32'b00000010000001101010111110100011;
ROM[53] <= 32'b00000100000001101010000000100011;
ROM[54] <= 32'b00000100000001101010000010100011;
ROM[55] <= 32'b00000100000001101010000100100011;
ROM[56] <= 32'b00000100000001101010000110100011;
ROM[57] <= 32'b00000100000001101010001000100011;
ROM[58] <= 32'b00000100000001101010001010100011;
ROM[59] <= 32'b00000100000001101010001100100011;
ROM[60] <= 32'b00000100000001101010001110100011;
ROM[61] <= 32'b00000100000001101010010000100011;
ROM[62] <= 32'b00000100000001101010010010100011;
ROM[63] <= 32'b00000100000001101010010100100011;
ROM[64] <= 32'b00000100000001101010010110100011;
ROM[65] <= 32'b00000100000001101010011000100011;
ROM[66] <= 32'b00000100000001101010011010100011;
ROM[67] <= 32'b00000100000001101010011100100011;
ROM[68] <= 32'b00000100000001101010011110100011;
ROM[69] <= 32'b00000100000001101010100000100011;
ROM[70] <= 32'b00000100000001101010100010100011;
ROM[71] <= 32'b00000100000001101010100100100011;
ROM[72] <= 32'b00000100000001101010100110100011;
ROM[73] <= 32'b00000100000001101010101000100011;
ROM[74] <= 32'b00000100000001101010101010100011;
ROM[75] <= 32'b00000100000001101010101100100011;
ROM[76] <= 32'b00000100000001101010101110100011;
ROM[77] <= 32'b00000100000001101010110000100011;
ROM[78] <= 32'b00000100000001101010110010100011;
ROM[79] <= 32'b00000100000001101010110100100011;
ROM[80] <= 32'b00000100000001101010110110100011;
ROM[81] <= 32'b00000100000001101010111000100011;
ROM[82] <= 32'b00000100000001101010111010100011;
ROM[83] <= 32'b00000100000001101010111100100011;
ROM[84] <= 32'b00000100000001101010111110100011;
ROM[85] <= 32'b00000110000001101010000000100011;
ROM[86] <= 32'b00000110000001101010000010100011;
ROM[87] <= 32'b00000110000001101010000100100011;
ROM[88] <= 32'b00000110000001101010000110100011;
ROM[89] <= 32'b00000110000001101010001000100011;
ROM[90] <= 32'b00000110000001101010001010100011;
ROM[91] <= 32'b00000110000001101010001100100011;
ROM[92] <= 32'b00000110000001101010001110100011;
ROM[93] <= 32'b00000110000001101010010000100011;
ROM[94] <= 32'b00000110000001101010010010100011;
ROM[95] <= 32'b00000110000001101010010100100011;
ROM[96] <= 32'b00000110000001101010010110100011;
ROM[97] <= 32'b00000110000001101010011000100011;
ROM[98] <= 32'b00000110000001101010011010100011;
ROM[99] <= 32'b00000110000001101010011100100011;
ROM[100] <= 32'b00000110000001101010011110100011;
ROM[101] <= 32'b00000110000001101010100000100011;
ROM[102] <= 32'b00000110000001101010100010100011;
ROM[103] <= 32'b00000110000001101010100100100011;
ROM[104] <= 32'b00000110000001101010100110100011;
ROM[105] <= 32'b00000110000001101010101000100011;
ROM[106] <= 32'b00000110000001101010101010100011;
ROM[107] <= 32'b00000110000001101010101100100011;
ROM[108] <= 32'b00000110000001101010101110100011;
ROM[109] <= 32'b00000110000001101010110000100011;
ROM[110] <= 32'b00000110000001101010110010100011;
ROM[111] <= 32'b00000110000001101010110100100011;
ROM[112] <= 32'b00000110000001101010110110100011;
ROM[113] <= 32'b00000110000001101010111000100011;
ROM[114] <= 32'b00000110000001101010111010100011;
ROM[115] <= 32'b00000110000001101010111100100011;
ROM[116] <= 32'b00000110000001101010111110100011;
ROM[117] <= 32'b00001000000001101010000000100011;
ROM[118] <= 32'b00001000000001101010000010100011;
ROM[119] <= 32'b00001000000001101010000100100011;
ROM[120] <= 32'b00001000000001101010000110100011;
ROM[121] <= 32'b00001000000001101010001000100011;
ROM[122] <= 32'b00001000000001101010001010100011;
ROM[123] <= 32'b00001000000001101010001100100011;
ROM[124] <= 32'b00001000000001101010001110100011;
ROM[125] <= 32'b00001000000001101010010000100011;
ROM[126] <= 32'b00001000000001101010010010100011;
ROM[127] <= 32'b00001000000001101010010100100011;
ROM[128] <= 32'b00001000000001101010010110100011;
ROM[129] <= 32'b00001000000001101010011000100011;
ROM[130] <= 32'b00001000000001101010011010100011;
ROM[131] <= 32'b00001000000001101010011100100011;
ROM[132] <= 32'b00001000000001101010011110100011;
ROM[133] <= 32'b00001000000001101010100000100011;
ROM[134] <= 32'b00001000000001101010100010100011;
ROM[135] <= 32'b00001000000001101010100100100011;
ROM[136] <= 32'b00001000000001101010100110100011;
ROM[137] <= 32'b00001000000001101010101000100011;
ROM[138] <= 32'b00001000000001101010101010100011;
ROM[139] <= 32'b00001000000001101010101100100011;
ROM[140] <= 32'b00001000000001101010101110100011;
ROM[141] <= 32'b00001000000001101010110000100011;
ROM[142] <= 32'b00001000000001101010110010100011;
ROM[143] <= 32'b00001000000001101010110100100011;
ROM[144] <= 32'b00001000000001101010110110100011;
ROM[145] <= 32'b00001000000001101010111000100011;
ROM[146] <= 32'b00001000000001101010111010100011;
ROM[147] <= 32'b00001000000001101010111100100011;
ROM[148] <= 32'b00001000000001101010111110100011;
ROM[149] <= 32'b00001010000001101010000000100011;
ROM[150] <= 32'b00001010000001101010000010100011;
ROM[151] <= 32'b00001010000001101010000100100011;
ROM[152] <= 32'b00001010000001101010000110100011;
ROM[153] <= 32'b00001010000001101010001000100011;
ROM[154] <= 32'b00001010000001101010001010100011;
ROM[155] <= 32'b00001010000001101010001100100011;
ROM[156] <= 32'b00001010000001101010001110100011;
ROM[157] <= 32'b00001010000001101010010000100011;
ROM[158] <= 32'b00001010000001101010010010100011;
ROM[159] <= 32'b00001010000001101010010100100011;
ROM[160] <= 32'b00001010000001101010010110100011;
ROM[161] <= 32'b00001010000001101010011000100011;
ROM[162] <= 32'b00001010000001101010011010100011;
ROM[163] <= 32'b00001010000001101010011100100011;
ROM[164] <= 32'b00001010000001101010011110100011;
ROM[165] <= 32'b00001010000001101010100000100011;
ROM[166] <= 32'b00001010000001101010100010100011;
ROM[167] <= 32'b00001010000001101010100100100011;
ROM[168] <= 32'b00001010000001101010100110100011;
ROM[169] <= 32'b00001010000001101010101000100011;
ROM[170] <= 32'b00001010000001101010101010100011;
ROM[171] <= 32'b00001010000001101010101100100011;
ROM[172] <= 32'b00001010000001101010101110100011;
ROM[173] <= 32'b00001010000001101010110000100011;
ROM[174] <= 32'b00001010000001101010110010100011;
ROM[175] <= 32'b00001010000001101010110100100011;
ROM[176] <= 32'b00001010000001101010110110100011;
ROM[177] <= 32'b00001010000001101010111000100011;
ROM[178] <= 32'b00001010000001101010111010100011;
ROM[179] <= 32'b00001010000001101010111100100011;
ROM[180] <= 32'b00001010000001101010111110100011;
ROM[181] <= 32'b00001100000001101010000000100011;
ROM[182] <= 32'b00001100000001101010000010100011;
ROM[183] <= 32'b00001100000001101010000100100011;
ROM[184] <= 32'b00001100000001101010000110100011;
ROM[185] <= 32'b00001100000001101010001000100011;
ROM[186] <= 32'b00001100000001101010001010100011;
ROM[187] <= 32'b00001100000001101010001100100011;
ROM[188] <= 32'b00001100000001101010001110100011;
ROM[189] <= 32'b00001100000001101010010000100011;
ROM[190] <= 32'b00001100000001101010010010100011;
ROM[191] <= 32'b00001100000001101010010100100011;
ROM[192] <= 32'b00001100000001101010010110100011;
ROM[193] <= 32'b00001100000001101010011000100011;
ROM[194] <= 32'b00001100000001101010011010100011;
ROM[195] <= 32'b00001100000001101010011100100011;
ROM[196] <= 32'b00001100000001101010011110100011;
ROM[197] <= 32'b00001100000001101010100000100011;
ROM[198] <= 32'b00001100000001101010100010100011;
ROM[199] <= 32'b00001100000001101010100100100011;
ROM[200] <= 32'b00001100000001101010100110100011;
ROM[201] <= 32'b00001100000001101010101000100011;
ROM[202] <= 32'b00001100000001101010101010100011;
ROM[203] <= 32'b00001100000001101010101100100011;
ROM[204] <= 32'b00001100000001101010101110100011;
ROM[205] <= 32'b00001100000001101010110000100011;
ROM[206] <= 32'b00001100000001101010110010100011;
ROM[207] <= 32'b00001100000001101010110100100011;
ROM[208] <= 32'b00001100000001101010110110100011;
ROM[209] <= 32'b00001100000001101010111000100011;
ROM[210] <= 32'b00001100000001101010111010100011;
ROM[211] <= 32'b00001100000001101010111100100011;
ROM[212] <= 32'b00001100000001101010111110100011;
ROM[213] <= 32'b00001110000001101010000000100011;
ROM[214] <= 32'b00001110000001101010000010100011;
ROM[215] <= 32'b00001110000001101010000100100011;
ROM[216] <= 32'b00001110000001101010000110100011;
ROM[217] <= 32'b00001110000001101010001000100011;
ROM[218] <= 32'b00001110000001101010001010100011;
ROM[219] <= 32'b00001110000001101010001100100011;
ROM[220] <= 32'b00001110000001101010001110100011;
ROM[221] <= 32'b00001110000001101010010000100011;
ROM[222] <= 32'b00001110000001101010010010100011;
ROM[223] <= 32'b00001110000001101010010100100011;
ROM[224] <= 32'b00001110000001101010010110100011;
ROM[225] <= 32'b00001110000001101010011000100011;
ROM[226] <= 32'b00001110000001101010011010100011;
ROM[227] <= 32'b00001110000001101010011100100011;
ROM[228] <= 32'b00001110000001101010011110100011;
ROM[229] <= 32'b00001110000001101010100000100011;
ROM[230] <= 32'b00001110000001101010100010100011;
ROM[231] <= 32'b00001110000001101010100100100011;
ROM[232] <= 32'b00001110000001101010100110100011;
ROM[233] <= 32'b00001110000001101010101000100011;
ROM[234] <= 32'b00001110000001101010101010100011;
ROM[235] <= 32'b00001110000001101010101100100011;
ROM[236] <= 32'b00001110000001101010101110100011;
ROM[237] <= 32'b00001110000001101010110000100011;
ROM[238] <= 32'b00001110000001101010110010100011;
ROM[239] <= 32'b00001110000001101010110100100011;
ROM[240] <= 32'b00001110000001101010110110100011;
ROM[241] <= 32'b00001110000001101010111000100011;
ROM[242] <= 32'b00001110000001101010111010100011;
ROM[243] <= 32'b00001110000001101010111100100011;
ROM[244] <= 32'b00001110000001101010111110100011;
ROM[245] <= 32'b00010000000001101000000100010011;
ROM[246] <= 32'b00000000000000010000000110010011;
ROM[247] <= 32'b00000000000001101000011000010011;
ROM[248] <= 32'b00000000000000010010000000100011;
ROM[249] <= 32'b00000000010000010000000100010011;
ROM[250] <= 32'b00000000101000000000001110010011;
ROM[251] <= 32'b00000000011100010010000000100011;
ROM[252] <= 32'b00000000010000010000000100010011;
ROM[253] <= 32'b00000000000000000000001110110111;
ROM[254] <= 32'b01000100000000111000001110010011;
ROM[255] <= 32'b00000000111000111000001110110011;
ROM[256] <= 32'b00000000011100010010000000100011;
ROM[257] <= 32'b00000000010000010000000100010011;
ROM[258] <= 32'b00000000001100010010000000100011;
ROM[259] <= 32'b00000000010000010000000100010011;
ROM[260] <= 32'b00000000010000010010000000100011;
ROM[261] <= 32'b00000000010000010000000100010011;
ROM[262] <= 32'b00000000010100010010000000100011;
ROM[263] <= 32'b00000000010000010000000100010011;
ROM[264] <= 32'b00000000011000010010000000100011;
ROM[265] <= 32'b00000000010000010000000100010011;
ROM[266] <= 32'b00000001010000000000001110010011;
ROM[267] <= 32'b00000000010000111000001110010011;
ROM[268] <= 32'b01000000011100010000001110110011;
ROM[269] <= 32'b00000000011100000000001000110011;
ROM[270] <= 32'b00000000001000000000000110110011;
ROM[271] <= 32'b00000001010000000000000011101111;
ROM[272] <= 32'b11111111110000010000000100010011;
ROM[273] <= 32'b00000000000000010010001110000011;
ROM[274] <= 32'b00000000011100011010000000100011;
ROM[275] <= 32'b00100010110100000001000011101111;
ROM[276] <= 32'b00000000000000010010000000100011;
ROM[277] <= 32'b00000000010000010000000100010011;
ROM[278] <= 32'b00000000010100000000001110010011;
ROM[279] <= 32'b00000000011100010010000000100011;
ROM[280] <= 32'b00000000010000010000000100010011;
ROM[281] <= 32'b00000000000000000000001110110111;
ROM[282] <= 32'b01001011000000111000001110010011;
ROM[283] <= 32'b00000000111000111000001110110011;
ROM[284] <= 32'b00000000011100010010000000100011;
ROM[285] <= 32'b00000000010000010000000100010011;
ROM[286] <= 32'b00000000001100010010000000100011;
ROM[287] <= 32'b00000000010000010000000100010011;
ROM[288] <= 32'b00000000010000010010000000100011;
ROM[289] <= 32'b00000000010000010000000100010011;
ROM[290] <= 32'b00000000010100010010000000100011;
ROM[291] <= 32'b00000000010000010000000100010011;
ROM[292] <= 32'b00000000011000010010000000100011;
ROM[293] <= 32'b00000000010000010000000100010011;
ROM[294] <= 32'b00000001010000000000001110010011;
ROM[295] <= 32'b00000000010000111000001110010011;
ROM[296] <= 32'b01000000011100010000001110110011;
ROM[297] <= 32'b00000000011100000000001000110011;
ROM[298] <= 32'b00000000001000000000000110110011;
ROM[299] <= 32'b00001110010000000000000011101111;
ROM[300] <= 32'b11111111110000010000000100010011;
ROM[301] <= 32'b00000000000000010010001110000011;
ROM[302] <= 32'b00000000011100011010000000100011;
ROM[303] <= 32'b00000000000000100010001110000011;
ROM[304] <= 32'b00000000011100010010000000100011;
ROM[305] <= 32'b00000000010000010000000100010011;
ROM[306] <= 32'b00000000000000011010001110000011;
ROM[307] <= 32'b00000000011100010010000000100011;
ROM[308] <= 32'b00000000010000010000000100010011;
ROM[309] <= 32'b00000000001000000000001110010011;
ROM[310] <= 32'b00000000011100010010000000100011;
ROM[311] <= 32'b00000000010000010000000100010011;
ROM[312] <= 32'b11111111110000010000000100010011;
ROM[313] <= 32'b00000000000000010010001110000011;
ROM[314] <= 32'b11111111110000010000000100010011;
ROM[315] <= 32'b00000000000000010010010000000011;
ROM[316] <= 32'b00000000100000111000001110110011;
ROM[317] <= 32'b00000000011100010010000000100011;
ROM[318] <= 32'b00000000010000010000000100010011;
ROM[319] <= 32'b11111111110000010000000100010011;
ROM[320] <= 32'b00000000000000010010001110000011;
ROM[321] <= 32'b00000000011100110010001000100011;
ROM[322] <= 32'b11111111110000010000000100010011;
ROM[323] <= 32'b00000000000000010010001110000011;
ROM[324] <= 32'b00000000011100110010000000100011;
ROM[325] <= 32'b00000000000000011010001110000011;
ROM[326] <= 32'b00000000011100010010000000100011;
ROM[327] <= 32'b00000000010000010000000100010011;
ROM[328] <= 32'b00000000001000000000001110010011;
ROM[329] <= 32'b00000000011100010010000000100011;
ROM[330] <= 32'b00000000010000010000000100010011;
ROM[331] <= 32'b11111111110000010000000100010011;
ROM[332] <= 32'b00000000000000010010001110000011;
ROM[333] <= 32'b11111111110000010000000100010011;
ROM[334] <= 32'b00000000000000010010010000000011;
ROM[335] <= 32'b00000000100000111000001110110011;
ROM[336] <= 32'b00000000011100010010000000100011;
ROM[337] <= 32'b00000000010000010000000100010011;
ROM[338] <= 32'b11111111110000010000000100010011;
ROM[339] <= 32'b00000000000000010010001110000011;
ROM[340] <= 32'b00000000011100110010001000100011;
ROM[341] <= 32'b00000000000000110010001110000011;
ROM[342] <= 32'b00000000011100010010000000100011;
ROM[343] <= 32'b00000000010000010000000100010011;
ROM[344] <= 32'b11111111110000010000000100010011;
ROM[345] <= 32'b00000000000000010010001110000011;
ROM[346] <= 32'b00000000011100100010000000100011;
ROM[347] <= 32'b00000000010000100000000100010011;
ROM[348] <= 32'b00000001010000000000001110010011;
ROM[349] <= 32'b01000000011100011000001110110011;
ROM[350] <= 32'b00000000000000111010000010000011;
ROM[351] <= 32'b00000000010000111010000110000011;
ROM[352] <= 32'b00000000100000111010001000000011;
ROM[353] <= 32'b00000000110000111010001010000011;
ROM[354] <= 32'b00000001000000111010001100000011;
ROM[355] <= 32'b00000000000000001000000011100111;
ROM[356] <= 32'b00000000000000100010001110000011;
ROM[357] <= 32'b00000000011100010010000000100011;
ROM[358] <= 32'b00000000010000010000000100010011;
ROM[359] <= 32'b00000000000000000000001110110111;
ROM[360] <= 32'b01011110100000111000001110010011;
ROM[361] <= 32'b00000000111000111000001110110011;
ROM[362] <= 32'b00000000011100010010000000100011;
ROM[363] <= 32'b00000000010000010000000100010011;
ROM[364] <= 32'b00000000001100010010000000100011;
ROM[365] <= 32'b00000000010000010000000100010011;
ROM[366] <= 32'b00000000010000010010000000100011;
ROM[367] <= 32'b00000000010000010000000100010011;
ROM[368] <= 32'b00000000010100010010000000100011;
ROM[369] <= 32'b00000000010000010000000100010011;
ROM[370] <= 32'b00000000011000010010000000100011;
ROM[371] <= 32'b00000000010000010000000100010011;
ROM[372] <= 32'b00000001010000000000001110010011;
ROM[373] <= 32'b00000000010000111000001110010011;
ROM[374] <= 32'b01000000011100010000001110110011;
ROM[375] <= 32'b00000000011100000000001000110011;
ROM[376] <= 32'b00000000001000000000000110110011;
ROM[377] <= 32'b01111101000000000000000011101111;
ROM[378] <= 32'b11111111110000010000000100010011;
ROM[379] <= 32'b00000000000000010010001110000011;
ROM[380] <= 32'b00000000011100100010000000100011;
ROM[381] <= 32'b00000000010000100000000100010011;
ROM[382] <= 32'b00000001010000000000001110010011;
ROM[383] <= 32'b01000000011100011000001110110011;
ROM[384] <= 32'b00000000000000111010000010000011;
ROM[385] <= 32'b00000000010000111010000110000011;
ROM[386] <= 32'b00000000100000111010001000000011;
ROM[387] <= 32'b00000000110000111010001010000011;
ROM[388] <= 32'b00000001000000111010001100000011;
ROM[389] <= 32'b00000000000000001000000011100111;
ROM[390] <= 32'b00000000000000100010001110000011;
ROM[391] <= 32'b00000000011100010010000000100011;
ROM[392] <= 32'b00000000010000010000000100010011;
ROM[393] <= 32'b11111111110000010000000100010011;
ROM[394] <= 32'b00000000000000010010001110000011;
ROM[395] <= 32'b00000000011100101010000000100011;
ROM[396] <= 32'b00000000000000101010001110000011;
ROM[397] <= 32'b00000000011100010010000000100011;
ROM[398] <= 32'b00000000010000010000000100010011;
ROM[399] <= 32'b00000000000000000000001110110111;
ROM[400] <= 32'b01101000100000111000001110010011;
ROM[401] <= 32'b00000000111000111000001110110011;
ROM[402] <= 32'b00000000011100010010000000100011;
ROM[403] <= 32'b00000000010000010000000100010011;
ROM[404] <= 32'b00000000001100010010000000100011;
ROM[405] <= 32'b00000000010000010000000100010011;
ROM[406] <= 32'b00000000010000010010000000100011;
ROM[407] <= 32'b00000000010000010000000100010011;
ROM[408] <= 32'b00000000010100010010000000100011;
ROM[409] <= 32'b00000000010000010000000100010011;
ROM[410] <= 32'b00000000011000010010000000100011;
ROM[411] <= 32'b00000000010000010000000100010011;
ROM[412] <= 32'b00000001010000000000001110010011;
ROM[413] <= 32'b00000000010000111000001110010011;
ROM[414] <= 32'b01000000011100010000001110110011;
ROM[415] <= 32'b00000000011100000000001000110011;
ROM[416] <= 32'b00000000001000000000000110110011;
ROM[417] <= 32'b01001110100100000000000011101111;
ROM[418] <= 32'b11111111110000010000000100010011;
ROM[419] <= 32'b00000000000000010010001110000011;
ROM[420] <= 32'b00000000011101100010000000100011;
ROM[421] <= 32'b00000000000000000000001110010011;
ROM[422] <= 32'b00000000011100010010000000100011;
ROM[423] <= 32'b00000000010000010000000100010011;
ROM[424] <= 32'b11111111110000010000000100010011;
ROM[425] <= 32'b00000000000000010010001110000011;
ROM[426] <= 32'b00000000011100100010000000100011;
ROM[427] <= 32'b00000000010000100000000100010011;
ROM[428] <= 32'b00000001010000000000001110010011;
ROM[429] <= 32'b01000000011100011000001110110011;
ROM[430] <= 32'b00000000000000111010000010000011;
ROM[431] <= 32'b00000000010000111010000110000011;
ROM[432] <= 32'b00000000100000111010001000000011;
ROM[433] <= 32'b00000000110000111010001010000011;
ROM[434] <= 32'b00000001000000111010001100000011;
ROM[435] <= 32'b00000000000000001000000011100111;
ROM[436] <= 32'b00000000000000000100001110110111;
ROM[437] <= 32'b00000000011100010010000000100011;
ROM[438] <= 32'b00000000010000010000000100010011;
ROM[439] <= 32'b11111111110000010000000100010011;
ROM[440] <= 32'b00000000000000010010001110000011;
ROM[441] <= 32'b00000000011101101010011110100011;
ROM[442] <= 32'b10000000000000000000001110010011;
ROM[443] <= 32'b00000000011100010010000000100011;
ROM[444] <= 32'b00000000010000010000000100010011;
ROM[445] <= 32'b11111111110000010000000100010011;
ROM[446] <= 32'b00000000000000010010001110000011;
ROM[447] <= 32'b00000000011101101010100000100011;
ROM[448] <= 32'b00000000000000000000001110010011;
ROM[449] <= 32'b00000000011100010010000000100011;
ROM[450] <= 32'b00000000010000010000000100010011;
ROM[451] <= 32'b11111111110000010000000100010011;
ROM[452] <= 32'b00000000000000010010001110000011;
ROM[453] <= 32'b00000000011101101010100010100011;
ROM[454] <= 32'b00000000111101101010001110000011;
ROM[455] <= 32'b00000000011100010010000000100011;
ROM[456] <= 32'b00000000010000010000000100010011;
ROM[457] <= 32'b11111111110000010000000100010011;
ROM[458] <= 32'b00000000000000010010001110000011;
ROM[459] <= 32'b00000000011101101010100100100011;
ROM[460] <= 32'b00000000000000000000001110010011;
ROM[461] <= 32'b00000000011100010010000000100011;
ROM[462] <= 32'b00000000010000010000000100010011;
ROM[463] <= 32'b11111111110000010000000100010011;
ROM[464] <= 32'b00000000000000010010001110000011;
ROM[465] <= 32'b00000000011101101010100110100011;
ROM[466] <= 32'b00000000000100000000001110010011;
ROM[467] <= 32'b00000000011100010010000000100011;
ROM[468] <= 32'b00000000010000010000000100010011;
ROM[469] <= 32'b11111111110000010000000100010011;
ROM[470] <= 32'b00000000000000010010001110000011;
ROM[471] <= 32'b01000000011100000000001110110011;
ROM[472] <= 32'b00000000011100010010000000100011;
ROM[473] <= 32'b00000000010000010000000100010011;
ROM[474] <= 32'b11111111110000010000000100010011;
ROM[475] <= 32'b00000000000000010010001110000011;
ROM[476] <= 32'b00000000011101101010101000100011;
ROM[477] <= 32'b00000000111101101010001110000011;
ROM[478] <= 32'b00000000011100010010000000100011;
ROM[479] <= 32'b00000000010000010000000100010011;
ROM[480] <= 32'b00000001000001101010001110000011;
ROM[481] <= 32'b00000000011100010010000000100011;
ROM[482] <= 32'b00000000010000010000000100010011;
ROM[483] <= 32'b11111111110000010000000100010011;
ROM[484] <= 32'b00000000000000010010001110000011;
ROM[485] <= 32'b11111111110000010000000100010011;
ROM[486] <= 32'b00000000000000010010010000000011;
ROM[487] <= 32'b01000000100000111000001110110011;
ROM[488] <= 32'b00000000011100010010000000100011;
ROM[489] <= 32'b00000000010000010000000100010011;
ROM[490] <= 32'b00000001001001101010001110000011;
ROM[491] <= 32'b00000000011100010010000000100011;
ROM[492] <= 32'b00000000010000010000000100010011;
ROM[493] <= 32'b00000001001101101010001110000011;
ROM[494] <= 32'b00000000011100010010000000100011;
ROM[495] <= 32'b00000000010000010000000100010011;
ROM[496] <= 32'b11111111110000010000000100010011;
ROM[497] <= 32'b00000000000000010010001110000011;
ROM[498] <= 32'b11111111110000010000000100010011;
ROM[499] <= 32'b00000000000000010010010000000011;
ROM[500] <= 32'b00000000100000111000001110110011;
ROM[501] <= 32'b00000000011100010010000000100011;
ROM[502] <= 32'b00000000010000010000000100010011;
ROM[503] <= 32'b11111111110000010000000100010011;
ROM[504] <= 32'b00000000000000010010001110000011;
ROM[505] <= 32'b00000000011100110010001000100011;
ROM[506] <= 32'b11111111110000010000000100010011;
ROM[507] <= 32'b00000000000000010010001110000011;
ROM[508] <= 32'b00000000011100110010000000100011;
ROM[509] <= 32'b00000000000000000000001110010011;
ROM[510] <= 32'b00000000011100010010000000100011;
ROM[511] <= 32'b00000000010000010000000100010011;
ROM[512] <= 32'b00000001001001101010001110000011;
ROM[513] <= 32'b00000000011100010010000000100011;
ROM[514] <= 32'b00000000010000010000000100010011;
ROM[515] <= 32'b00000001010001101010001110000011;
ROM[516] <= 32'b00000000011100010010000000100011;
ROM[517] <= 32'b00000000010000010000000100010011;
ROM[518] <= 32'b11111111110000010000000100010011;
ROM[519] <= 32'b00000000000000010010001110000011;
ROM[520] <= 32'b11111111110000010000000100010011;
ROM[521] <= 32'b00000000000000010010010000000011;
ROM[522] <= 32'b00000000100000111000001110110011;
ROM[523] <= 32'b00000000011100010010000000100011;
ROM[524] <= 32'b00000000010000010000000100010011;
ROM[525] <= 32'b11111111110000010000000100010011;
ROM[526] <= 32'b00000000000000010010001110000011;
ROM[527] <= 32'b00000000011100110010001000100011;
ROM[528] <= 32'b11111111110000010000000100010011;
ROM[529] <= 32'b00000000000000010010001110000011;
ROM[530] <= 32'b00000000011100110010000000100011;
ROM[531] <= 32'b00000000000100000000001110010011;
ROM[532] <= 32'b00000000011100010010000000100011;
ROM[533] <= 32'b00000000010000010000000100010011;
ROM[534] <= 32'b11111111110000010000000100010011;
ROM[535] <= 32'b00000000000000010010001110000011;
ROM[536] <= 32'b00000000011101101010101010100011;
ROM[537] <= 32'b00000000000000000000001110010011;
ROM[538] <= 32'b00000000011100010010000000100011;
ROM[539] <= 32'b00000000010000010000000100010011;
ROM[540] <= 32'b11111111110000010000000100010011;
ROM[541] <= 32'b00000000000000010010001110000011;
ROM[542] <= 32'b00000000011100100010000000100011;
ROM[543] <= 32'b00000000010000100000000100010011;
ROM[544] <= 32'b00000001010000000000001110010011;
ROM[545] <= 32'b01000000011100011000001110110011;
ROM[546] <= 32'b00000000000000111010000010000011;
ROM[547] <= 32'b00000000010000111010000110000011;
ROM[548] <= 32'b00000000100000111010001000000011;
ROM[549] <= 32'b00000000110000111010001010000011;
ROM[550] <= 32'b00000001000000111010001100000011;
ROM[551] <= 32'b00000000000000001000000011100111;
ROM[552] <= 32'b00000001000101101010001110000011;
ROM[553] <= 32'b00000000011100010010000000100011;
ROM[554] <= 32'b00000000010000010000000100010011;
ROM[555] <= 32'b00000000000000100010001110000011;
ROM[556] <= 32'b00000000011100010010000000100011;
ROM[557] <= 32'b00000000010000010000000100010011;
ROM[558] <= 32'b11111111110000010000000100010011;
ROM[559] <= 32'b00000000000000010010001110000011;
ROM[560] <= 32'b11111111110000010000000100010011;
ROM[561] <= 32'b00000000000000010010010000000011;
ROM[562] <= 32'b00000000100000111000001110110011;
ROM[563] <= 32'b00000000011100010010000000100011;
ROM[564] <= 32'b00000000010000010000000100010011;
ROM[565] <= 32'b11111111110000010000000100010011;
ROM[566] <= 32'b00000000000000010010001110000011;
ROM[567] <= 32'b00000000011100110010001000100011;
ROM[568] <= 32'b00000000000000110010001110000011;
ROM[569] <= 32'b00000000011100010010000000100011;
ROM[570] <= 32'b00000000010000010000000100010011;
ROM[571] <= 32'b11111111110000010000000100010011;
ROM[572] <= 32'b00000000000000010010001110000011;
ROM[573] <= 32'b00000000011100100010000000100011;
ROM[574] <= 32'b00000000010000100000000100010011;
ROM[575] <= 32'b00000001010000000000001110010011;
ROM[576] <= 32'b01000000011100011000001110110011;
ROM[577] <= 32'b00000000000000111010000010000011;
ROM[578] <= 32'b00000000010000111010000110000011;
ROM[579] <= 32'b00000000100000111010001000000011;
ROM[580] <= 32'b00000000110000111010001010000011;
ROM[581] <= 32'b00000001000000111010001100000011;
ROM[582] <= 32'b00000000000000001000000011100111;
ROM[583] <= 32'b00000000010000100010001110000011;
ROM[584] <= 32'b00000000011100010010000000100011;
ROM[585] <= 32'b00000000010000010000000100010011;
ROM[586] <= 32'b00000001000101101010001110000011;
ROM[587] <= 32'b00000000011100010010000000100011;
ROM[588] <= 32'b00000000010000010000000100010011;
ROM[589] <= 32'b00000000000000100010001110000011;
ROM[590] <= 32'b00000000011100010010000000100011;
ROM[591] <= 32'b00000000010000010000000100010011;
ROM[592] <= 32'b11111111110000010000000100010011;
ROM[593] <= 32'b00000000000000010010001110000011;
ROM[594] <= 32'b11111111110000010000000100010011;
ROM[595] <= 32'b00000000000000010010010000000011;
ROM[596] <= 32'b00000000100000111000001110110011;
ROM[597] <= 32'b00000000011100010010000000100011;
ROM[598] <= 32'b00000000010000010000000100010011;
ROM[599] <= 32'b11111111110000010000000100010011;
ROM[600] <= 32'b00000000000000010010001110000011;
ROM[601] <= 32'b00000000011100110010001000100011;
ROM[602] <= 32'b11111111110000010000000100010011;
ROM[603] <= 32'b00000000000000010010001110000011;
ROM[604] <= 32'b00000000011100110010000000100011;
ROM[605] <= 32'b00000000000000000000001110010011;
ROM[606] <= 32'b00000000011100010010000000100011;
ROM[607] <= 32'b00000000010000010000000100010011;
ROM[608] <= 32'b11111111110000010000000100010011;
ROM[609] <= 32'b00000000000000010010001110000011;
ROM[610] <= 32'b00000000011100100010000000100011;
ROM[611] <= 32'b00000000010000100000000100010011;
ROM[612] <= 32'b00000001010000000000001110010011;
ROM[613] <= 32'b01000000011100011000001110110011;
ROM[614] <= 32'b00000000000000111010000010000011;
ROM[615] <= 32'b00000000010000111010000110000011;
ROM[616] <= 32'b00000000100000111010001000000011;
ROM[617] <= 32'b00000000110000111010001010000011;
ROM[618] <= 32'b00000001000000111010001100000011;
ROM[619] <= 32'b00000000000000001000000011100111;
ROM[620] <= 32'b00000000000000010010000000100011;
ROM[621] <= 32'b00000000010000010000000100010011;
ROM[622] <= 32'b00000000000000010010000000100011;
ROM[623] <= 32'b00000000010000010000000100010011;
ROM[624] <= 32'b00000000000000010010000000100011;
ROM[625] <= 32'b00000000010000010000000100010011;
ROM[626] <= 32'b00000000000000010010000000100011;
ROM[627] <= 32'b00000000010000010000000100010011;
ROM[628] <= 32'b00000000000000000000001110010011;
ROM[629] <= 32'b00000000011100010010000000100011;
ROM[630] <= 32'b00000000010000010000000100010011;
ROM[631] <= 32'b11111111110000010000000100010011;
ROM[632] <= 32'b00000000000000010010001110000011;
ROM[633] <= 32'b00000000011100011010001000100011;
ROM[634] <= 32'b00000000111101101010001110000011;
ROM[635] <= 32'b00000000011100010010000000100011;
ROM[636] <= 32'b00000000010000010000000100010011;
ROM[637] <= 32'b00000001000001101010001110000011;
ROM[638] <= 32'b00000000011100010010000000100011;
ROM[639] <= 32'b00000000010000010000000100010011;
ROM[640] <= 32'b11111111110000010000000100010011;
ROM[641] <= 32'b00000000000000010010001110000011;
ROM[642] <= 32'b11111111110000010000000100010011;
ROM[643] <= 32'b00000000000000010010010000000011;
ROM[644] <= 32'b01000000100000111000001110110011;
ROM[645] <= 32'b00000000011100010010000000100011;
ROM[646] <= 32'b00000000010000010000000100010011;
ROM[647] <= 32'b11111111110000010000000100010011;
ROM[648] <= 32'b00000000000000010010001110000011;
ROM[649] <= 32'b00000000011100011010010000100011;
ROM[650] <= 32'b00000001001001101010001110000011;
ROM[651] <= 32'b00000000011100010010000000100011;
ROM[652] <= 32'b00000000010000010000000100010011;
ROM[653] <= 32'b11111111110000010000000100010011;
ROM[654] <= 32'b00000000000000010010001110000011;
ROM[655] <= 32'b00000000011100011010000000100011;
ROM[656] <= 32'b00000000000000011010001110000011;
ROM[657] <= 32'b00000000011100010010000000100011;
ROM[658] <= 32'b00000000010000010000000100010011;
ROM[659] <= 32'b00000001010001101010001110000011;
ROM[660] <= 32'b00000000011100010010000000100011;
ROM[661] <= 32'b00000000010000010000000100010011;
ROM[662] <= 32'b11111111110000010000000100010011;
ROM[663] <= 32'b00000000000000010010001110000011;
ROM[664] <= 32'b11111111110000010000000100010011;
ROM[665] <= 32'b00000000000000010010010000000011;
ROM[666] <= 32'b00000000100000111000001110110011;
ROM[667] <= 32'b00000000011100010010000000100011;
ROM[668] <= 32'b00000000010000010000000100010011;
ROM[669] <= 32'b11111111110000010000000100010011;
ROM[670] <= 32'b00000000000000010010001110000011;
ROM[671] <= 32'b00000000011100110010001000100011;
ROM[672] <= 32'b00000000000000110010001110000011;
ROM[673] <= 32'b00000000011100010010000000100011;
ROM[674] <= 32'b00000000010000010000000100010011;
ROM[675] <= 32'b00000000000000000000001110010011;
ROM[676] <= 32'b00000000011100010010000000100011;
ROM[677] <= 32'b00000000010000010000000100010011;
ROM[678] <= 32'b11111111110000010000000100010011;
ROM[679] <= 32'b00000000000000010010001110000011;
ROM[680] <= 32'b11111111110000010000000100010011;
ROM[681] <= 32'b00000000000000010010010000000011;
ROM[682] <= 32'b00000000011101000010010010110011;
ROM[683] <= 32'b00000000100000111010010100110011;
ROM[684] <= 32'b00000000101001001000001110110011;
ROM[685] <= 32'b00000000000100111000001110010011;
ROM[686] <= 32'b00000000000100111111001110010011;
ROM[687] <= 32'b00000000011100010010000000100011;
ROM[688] <= 32'b00000000010000010000000100010011;
ROM[689] <= 32'b11111111110000010000000100010011;
ROM[690] <= 32'b00000000000000010010001110000011;
ROM[691] <= 32'b00000000000000111000101001100011;
ROM[692] <= 32'b00000000000000000000001110110111;
ROM[693] <= 32'b10101110010000111000001110010011;
ROM[694] <= 32'b00000000111000111000001110110011;
ROM[695] <= 32'b00000000000000111000000011100111;
ROM[696] <= 32'b00000100000000000000000011101111;
ROM[697] <= 32'b00000000000000011010001110000011;
ROM[698] <= 32'b00000000011100010010000000100011;
ROM[699] <= 32'b00000000010000010000000100010011;
ROM[700] <= 32'b11111111110000010000000100010011;
ROM[701] <= 32'b00000000000000010010001110000011;
ROM[702] <= 32'b00000000011100100010000000100011;
ROM[703] <= 32'b00000000010000100000000100010011;
ROM[704] <= 32'b00000001010000000000001110010011;
ROM[705] <= 32'b01000000011100011000001110110011;
ROM[706] <= 32'b00000000000000111010000010000011;
ROM[707] <= 32'b00000000010000111010000110000011;
ROM[708] <= 32'b00000000100000111010001000000011;
ROM[709] <= 32'b00000000110000111010001010000011;
ROM[710] <= 32'b00000001000000111010001100000011;
ROM[711] <= 32'b00000000000000001000000011100111;
ROM[712] <= 32'b00000000000000011010001110000011;
ROM[713] <= 32'b00000000011100010010000000100011;
ROM[714] <= 32'b00000000010000010000000100010011;
ROM[715] <= 32'b00000000000000000000001110010011;
ROM[716] <= 32'b00000000011100010010000000100011;
ROM[717] <= 32'b00000000010000010000000100010011;
ROM[718] <= 32'b11111111110000010000000100010011;
ROM[719] <= 32'b00000000000000010010001110000011;
ROM[720] <= 32'b11111111110000010000000100010011;
ROM[721] <= 32'b00000000000000010010010000000011;
ROM[722] <= 32'b00000000011101000010010010110011;
ROM[723] <= 32'b00000000100000111010010100110011;
ROM[724] <= 32'b00000000101001001000001110110011;
ROM[725] <= 32'b00000000000100111000001110010011;
ROM[726] <= 32'b00000000000100111111001110010011;
ROM[727] <= 32'b00000000011100010010000000100011;
ROM[728] <= 32'b00000000010000010000000100010011;
ROM[729] <= 32'b11111111110000010000000100010011;
ROM[730] <= 32'b00000000000000010010001110000011;
ROM[731] <= 32'b01000000011100000000001110110011;
ROM[732] <= 32'b00000000000100111000001110010011;
ROM[733] <= 32'b00000000011100010010000000100011;
ROM[734] <= 32'b00000000010000010000000100010011;
ROM[735] <= 32'b11111111110000010000000100010011;
ROM[736] <= 32'b00000000000000010010001110000011;
ROM[737] <= 32'b01000000011100000000001110110011;
ROM[738] <= 32'b00000000000100111000001110010011;
ROM[739] <= 32'b00000000011100010010000000100011;
ROM[740] <= 32'b00000000010000010000000100010011;
ROM[741] <= 32'b11111111110000010000000100010011;
ROM[742] <= 32'b00000000000000010010001110000011;
ROM[743] <= 32'b00000000000000111000101001100011;
ROM[744] <= 32'b00000000000000000000001110110111;
ROM[745] <= 32'b11010111100000111000001110010011;
ROM[746] <= 32'b00000000111000111000001110110011;
ROM[747] <= 32'b00000000000000111000000011100111;
ROM[748] <= 32'b00000000000000011010001110000011;
ROM[749] <= 32'b00000000011100010010000000100011;
ROM[750] <= 32'b00000000010000010000000100010011;
ROM[751] <= 32'b00000001001101101010001110000011;
ROM[752] <= 32'b00000000011100010010000000100011;
ROM[753] <= 32'b00000000010000010000000100010011;
ROM[754] <= 32'b11111111110000010000000100010011;
ROM[755] <= 32'b00000000000000010010001110000011;
ROM[756] <= 32'b11111111110000010000000100010011;
ROM[757] <= 32'b00000000000000010010010000000011;
ROM[758] <= 32'b00000000100000111000001110110011;
ROM[759] <= 32'b00000000011100010010000000100011;
ROM[760] <= 32'b00000000010000010000000100010011;
ROM[761] <= 32'b11111111110000010000000100010011;
ROM[762] <= 32'b00000000000000010010001110000011;
ROM[763] <= 32'b00000000011100110010001000100011;
ROM[764] <= 32'b00000000000000110010001110000011;
ROM[765] <= 32'b00000000011100010010000000100011;
ROM[766] <= 32'b00000000010000010000000100010011;
ROM[767] <= 32'b00000000000100000000001110010011;
ROM[768] <= 32'b00000000011100010010000000100011;
ROM[769] <= 32'b00000000010000010000000100010011;
ROM[770] <= 32'b11111111110000010000000100010011;
ROM[771] <= 32'b00000000000000010010001110000011;
ROM[772] <= 32'b11111111110000010000000100010011;
ROM[773] <= 32'b00000000000000010010010000000011;
ROM[774] <= 32'b01000000100000111000001110110011;
ROM[775] <= 32'b00000000011100010010000000100011;
ROM[776] <= 32'b00000000010000010000000100010011;
ROM[777] <= 32'b11111111110000010000000100010011;
ROM[778] <= 32'b00000000000000010010001110000011;
ROM[779] <= 32'b00000000011100011010011000100011;
ROM[780] <= 32'b00000000110000011010001110000011;
ROM[781] <= 32'b00000000011100010010000000100011;
ROM[782] <= 32'b00000000010000010000000100010011;
ROM[783] <= 32'b00000000000000100010001110000011;
ROM[784] <= 32'b00000000011100010010000000100011;
ROM[785] <= 32'b00000000010000010000000100010011;
ROM[786] <= 32'b11111111110000010000000100010011;
ROM[787] <= 32'b00000000000000010010001110000011;
ROM[788] <= 32'b11111111110000010000000100010011;
ROM[789] <= 32'b00000000000000010010010000000011;
ROM[790] <= 32'b00000000011101000010001110110011;
ROM[791] <= 32'b00000000011100010010000000100011;
ROM[792] <= 32'b00000000010000010000000100010011;
ROM[793] <= 32'b11111111110000010000000100010011;
ROM[794] <= 32'b00000000000000010010001110000011;
ROM[795] <= 32'b01000000011100000000001110110011;
ROM[796] <= 32'b00000000000100111000001110010011;
ROM[797] <= 32'b00000000011100010010000000100011;
ROM[798] <= 32'b00000000010000010000000100010011;
ROM[799] <= 32'b00000000110000011010001110000011;
ROM[800] <= 32'b00000000011100010010000000100011;
ROM[801] <= 32'b00000000010000010000000100010011;
ROM[802] <= 32'b00000000100000011010001110000011;
ROM[803] <= 32'b00000000011100010010000000100011;
ROM[804] <= 32'b00000000010000010000000100010011;
ROM[805] <= 32'b11111111110000010000000100010011;
ROM[806] <= 32'b00000000000000010010001110000011;
ROM[807] <= 32'b11111111110000010000000100010011;
ROM[808] <= 32'b00000000000000010010010000000011;
ROM[809] <= 32'b00000000011101000010001110110011;
ROM[810] <= 32'b00000000011100010010000000100011;
ROM[811] <= 32'b00000000010000010000000100010011;
ROM[812] <= 32'b11111111110000010000000100010011;
ROM[813] <= 32'b00000000000000010010001110000011;
ROM[814] <= 32'b11111111110000010000000100010011;
ROM[815] <= 32'b00000000000000010010010000000011;
ROM[816] <= 32'b00000000100000111111001110110011;
ROM[817] <= 32'b00000000011100010010000000100011;
ROM[818] <= 32'b00000000010000010000000100010011;
ROM[819] <= 32'b11111111110000010000000100010011;
ROM[820] <= 32'b00000000000000010010001110000011;
ROM[821] <= 32'b00000000000000111000101001100011;
ROM[822] <= 32'b00000000000000000000001110110111;
ROM[823] <= 32'b11001110110000111000001110010011;
ROM[824] <= 32'b00000000111000111000001110110011;
ROM[825] <= 32'b00000000000000111000000011100111;
ROM[826] <= 32'b00000011010000000000000011101111;
ROM[827] <= 32'b00000000000000011010001110000011;
ROM[828] <= 32'b00000000011100010010000000100011;
ROM[829] <= 32'b00000000010000010000000100010011;
ROM[830] <= 32'b11111111110000010000000100010011;
ROM[831] <= 32'b00000000000000010010001110000011;
ROM[832] <= 32'b00000000011100011010001000100011;
ROM[833] <= 32'b00000000110000011010001110000011;
ROM[834] <= 32'b00000000011100010010000000100011;
ROM[835] <= 32'b00000000010000010000000100010011;
ROM[836] <= 32'b11111111110000010000000100010011;
ROM[837] <= 32'b00000000000000010010001110000011;
ROM[838] <= 32'b00000000011100011010010000100011;
ROM[839] <= 32'b00000000000000011010001110000011;
ROM[840] <= 32'b00000000011100010010000000100011;
ROM[841] <= 32'b00000000010000010000000100010011;
ROM[842] <= 32'b00000001010001101010001110000011;
ROM[843] <= 32'b00000000011100010010000000100011;
ROM[844] <= 32'b00000000010000010000000100010011;
ROM[845] <= 32'b11111111110000010000000100010011;
ROM[846] <= 32'b00000000000000010010001110000011;
ROM[847] <= 32'b11111111110000010000000100010011;
ROM[848] <= 32'b00000000000000010010010000000011;
ROM[849] <= 32'b00000000100000111000001110110011;
ROM[850] <= 32'b00000000011100010010000000100011;
ROM[851] <= 32'b00000000010000010000000100010011;
ROM[852] <= 32'b11111111110000010000000100010011;
ROM[853] <= 32'b00000000000000010010001110000011;
ROM[854] <= 32'b00000000011100110010001000100011;
ROM[855] <= 32'b00000000000000110010001110000011;
ROM[856] <= 32'b00000000011100010010000000100011;
ROM[857] <= 32'b00000000010000010000000100010011;
ROM[858] <= 32'b11111111110000010000000100010011;
ROM[859] <= 32'b00000000000000010010001110000011;
ROM[860] <= 32'b00000000011100011010000000100011;
ROM[861] <= 32'b11011010110111111111000011101111;
ROM[862] <= 32'b00000000010000011010001110000011;
ROM[863] <= 32'b00000000011100010010000000100011;
ROM[864] <= 32'b00000000010000010000000100010011;
ROM[865] <= 32'b11111111110000010000000100010011;
ROM[866] <= 32'b00000000000000010010001110000011;
ROM[867] <= 32'b00000000011100100010000000100011;
ROM[868] <= 32'b00000000010000100000000100010011;
ROM[869] <= 32'b00000001010000000000001110010011;
ROM[870] <= 32'b01000000011100011000001110110011;
ROM[871] <= 32'b00000000000000111010000010000011;
ROM[872] <= 32'b00000000010000111010000110000011;
ROM[873] <= 32'b00000000100000111010001000000011;
ROM[874] <= 32'b00000000110000111010001010000011;
ROM[875] <= 32'b00000001000000111010001100000011;
ROM[876] <= 32'b00000000000000001000000011100111;
ROM[877] <= 32'b00000000000000010010000000100011;
ROM[878] <= 32'b00000000010000010000000100010011;
ROM[879] <= 32'b00000000000000010010000000100011;
ROM[880] <= 32'b00000000010000010000000100010011;
ROM[881] <= 32'b00000000000000010010000000100011;
ROM[882] <= 32'b00000000010000010000000100010011;
ROM[883] <= 32'b00000000000000100010001110000011;
ROM[884] <= 32'b00000000011100010010000000100011;
ROM[885] <= 32'b00000000010000010000000100010011;
ROM[886] <= 32'b00000000000000000000001110110111;
ROM[887] <= 32'b11100010010000111000001110010011;
ROM[888] <= 32'b00000000111000111000001110110011;
ROM[889] <= 32'b00000000011100010010000000100011;
ROM[890] <= 32'b00000000010000010000000100010011;
ROM[891] <= 32'b00000000001100010010000000100011;
ROM[892] <= 32'b00000000010000010000000100010011;
ROM[893] <= 32'b00000000010000010010000000100011;
ROM[894] <= 32'b00000000010000010000000100010011;
ROM[895] <= 32'b00000000010100010010000000100011;
ROM[896] <= 32'b00000000010000010000000100010011;
ROM[897] <= 32'b00000000011000010010000000100011;
ROM[898] <= 32'b00000000010000010000000100010011;
ROM[899] <= 32'b00000001010000000000001110010011;
ROM[900] <= 32'b00000000010000111000001110010011;
ROM[901] <= 32'b01000000011100010000001110110011;
ROM[902] <= 32'b00000000011100000000001000110011;
ROM[903] <= 32'b00000000001000000000000110110011;
ROM[904] <= 32'b10111001000111111111000011101111;
ROM[905] <= 32'b11111111110000010000000100010011;
ROM[906] <= 32'b00000000000000010010001110000011;
ROM[907] <= 32'b00000000011100011010000000100011;
ROM[908] <= 32'b00000000000000011010001110000011;
ROM[909] <= 32'b00000000011100010010000000100011;
ROM[910] <= 32'b00000000010000010000000100010011;
ROM[911] <= 32'b00000000000100000000001110010011;
ROM[912] <= 32'b00000000011100010010000000100011;
ROM[913] <= 32'b00000000010000010000000100010011;
ROM[914] <= 32'b11111111110000010000000100010011;
ROM[915] <= 32'b00000000000000010010001110000011;
ROM[916] <= 32'b11111111110000010000000100010011;
ROM[917] <= 32'b00000000000000010010010000000011;
ROM[918] <= 32'b01000000100000111000001110110011;
ROM[919] <= 32'b00000000011100010010000000100011;
ROM[920] <= 32'b00000000010000010000000100010011;
ROM[921] <= 32'b11111111110000010000000100010011;
ROM[922] <= 32'b00000000000000010010001110000011;
ROM[923] <= 32'b00000000011100011010010000100011;
ROM[924] <= 32'b00000000000000011010001110000011;
ROM[925] <= 32'b00000000011100010010000000100011;
ROM[926] <= 32'b00000000010000010000000100010011;
ROM[927] <= 32'b00000000000000000000001110010011;
ROM[928] <= 32'b00000000011100010010000000100011;
ROM[929] <= 32'b00000000010000010000000100010011;
ROM[930] <= 32'b11111111110000010000000100010011;
ROM[931] <= 32'b00000000000000010010001110000011;
ROM[932] <= 32'b11111111110000010000000100010011;
ROM[933] <= 32'b00000000000000010010010000000011;
ROM[934] <= 32'b00000000011101000010010010110011;
ROM[935] <= 32'b00000000100000111010010100110011;
ROM[936] <= 32'b00000000101001001000001110110011;
ROM[937] <= 32'b00000000000100111000001110010011;
ROM[938] <= 32'b00000000000100111111001110010011;
ROM[939] <= 32'b00000000011100010010000000100011;
ROM[940] <= 32'b00000000010000010000000100010011;
ROM[941] <= 32'b11111111110000010000000100010011;
ROM[942] <= 32'b00000000000000010010001110000011;
ROM[943] <= 32'b01000000011100000000001110110011;
ROM[944] <= 32'b00000000000100111000001110010011;
ROM[945] <= 32'b00000000011100010010000000100011;
ROM[946] <= 32'b00000000010000010000000100010011;
ROM[947] <= 32'b11111111110000010000000100010011;
ROM[948] <= 32'b00000000000000010010001110000011;
ROM[949] <= 32'b00000000000000111000101001100011;
ROM[950] <= 32'b00000000000000000000001110110111;
ROM[951] <= 32'b11101110110000111000001110010011;
ROM[952] <= 32'b00000000111000111000001110110011;
ROM[953] <= 32'b00000000000000111000000011100111;
ROM[954] <= 32'b01000100100000000000000011101111;
ROM[955] <= 32'b00000000000000011010001110000011;
ROM[956] <= 32'b00000000011100010010000000100011;
ROM[957] <= 32'b00000000010000010000000100010011;
ROM[958] <= 32'b00000001001101101010001110000011;
ROM[959] <= 32'b00000000011100010010000000100011;
ROM[960] <= 32'b00000000010000010000000100010011;
ROM[961] <= 32'b11111111110000010000000100010011;
ROM[962] <= 32'b00000000000000010010001110000011;
ROM[963] <= 32'b11111111110000010000000100010011;
ROM[964] <= 32'b00000000000000010010010000000011;
ROM[965] <= 32'b00000000100000111000001110110011;
ROM[966] <= 32'b00000000011100010010000000100011;
ROM[967] <= 32'b00000000010000010000000100010011;
ROM[968] <= 32'b11111111110000010000000100010011;
ROM[969] <= 32'b00000000000000010010001110000011;
ROM[970] <= 32'b00000000011100110010001000100011;
ROM[971] <= 32'b00000000000000110010001110000011;
ROM[972] <= 32'b00000000011100010010000000100011;
ROM[973] <= 32'b00000000010000010000000100010011;
ROM[974] <= 32'b00000000000000100010001110000011;
ROM[975] <= 32'b00000000011100010010000000100011;
ROM[976] <= 32'b00000000010000010000000100010011;
ROM[977] <= 32'b00000000001100000000001110010011;
ROM[978] <= 32'b00000000011100010010000000100011;
ROM[979] <= 32'b00000000010000010000000100010011;
ROM[980] <= 32'b11111111110000010000000100010011;
ROM[981] <= 32'b00000000000000010010001110000011;
ROM[982] <= 32'b11111111110000010000000100010011;
ROM[983] <= 32'b00000000000000010010010000000011;
ROM[984] <= 32'b00000000100000111000001110110011;
ROM[985] <= 32'b00000000011100010010000000100011;
ROM[986] <= 32'b00000000010000010000000100010011;
ROM[987] <= 32'b11111111110000010000000100010011;
ROM[988] <= 32'b00000000000000010010001110000011;
ROM[989] <= 32'b11111111110000010000000100010011;
ROM[990] <= 32'b00000000000000010010010000000011;
ROM[991] <= 32'b00000000100000111010001110110011;
ROM[992] <= 32'b00000000011100010010000000100011;
ROM[993] <= 32'b00000000010000010000000100010011;
ROM[994] <= 32'b11111111110000010000000100010011;
ROM[995] <= 32'b00000000000000010010001110000011;
ROM[996] <= 32'b00000000000000111000101001100011;
ROM[997] <= 32'b00000000000000000001001110110111;
ROM[998] <= 32'b00001001100000111000001110010011;
ROM[999] <= 32'b00000000111000111000001110110011;
ROM[1000] <= 32'b00000000000000111000000011100111;
ROM[1001] <= 32'b00000000000000011010001110000011;
ROM[1002] <= 32'b00000000011100010010000000100011;
ROM[1003] <= 32'b00000000010000010000000100010011;
ROM[1004] <= 32'b00000001010001101010001110000011;
ROM[1005] <= 32'b00000000011100010010000000100011;
ROM[1006] <= 32'b00000000010000010000000100010011;
ROM[1007] <= 32'b11111111110000010000000100010011;
ROM[1008] <= 32'b00000000000000010010001110000011;
ROM[1009] <= 32'b11111111110000010000000100010011;
ROM[1010] <= 32'b00000000000000010010010000000011;
ROM[1011] <= 32'b00000000100000111000001110110011;
ROM[1012] <= 32'b00000000011100010010000000100011;
ROM[1013] <= 32'b00000000010000010000000100010011;
ROM[1014] <= 32'b11111111110000010000000100010011;
ROM[1015] <= 32'b00000000000000010010001110000011;
ROM[1016] <= 32'b00000000011100110010001000100011;
ROM[1017] <= 32'b00000000000000110010001110000011;
ROM[1018] <= 32'b00000000011100010010000000100011;
ROM[1019] <= 32'b00000000010000010000000100010011;
ROM[1020] <= 32'b11111111110000010000000100010011;
ROM[1021] <= 32'b00000000000000010010001110000011;
ROM[1022] <= 32'b00000000011100011010001000100011;
ROM[1023] <= 32'b00000000000000011010001110000011;
ROM[1024] <= 32'b00000000011100010010000000100011;
ROM[1025] <= 32'b00000000010000010000000100010011;
ROM[1026] <= 32'b00000001001101101010001110000011;
ROM[1027] <= 32'b00000000011100010010000000100011;
ROM[1028] <= 32'b00000000010000010000000100010011;
ROM[1029] <= 32'b11111111110000010000000100010011;
ROM[1030] <= 32'b00000000000000010010001110000011;
ROM[1031] <= 32'b11111111110000010000000100010011;
ROM[1032] <= 32'b00000000000000010010010000000011;
ROM[1033] <= 32'b00000000100000111000001110110011;
ROM[1034] <= 32'b00000000011100010010000000100011;
ROM[1035] <= 32'b00000000010000010000000100010011;
ROM[1036] <= 32'b11111111110000010000000100010011;
ROM[1037] <= 32'b00000000000000010010001110000011;
ROM[1038] <= 32'b00000000011100110010001000100011;
ROM[1039] <= 32'b00000000000000110010001110000011;
ROM[1040] <= 32'b00000000011100010010000000100011;
ROM[1041] <= 32'b00000000010000010000000100010011;
ROM[1042] <= 32'b00000000100000011010001110000011;
ROM[1043] <= 32'b00000000011100010010000000100011;
ROM[1044] <= 32'b00000000010000010000000100010011;
ROM[1045] <= 32'b00000001010101101010001110000011;
ROM[1046] <= 32'b00000000011100010010000000100011;
ROM[1047] <= 32'b00000000010000010000000100010011;
ROM[1048] <= 32'b11111111110000010000000100010011;
ROM[1049] <= 32'b00000000000000010010001110000011;
ROM[1050] <= 32'b11111111110000010000000100010011;
ROM[1051] <= 32'b00000000000000010010010000000011;
ROM[1052] <= 32'b00000000100000111000001110110011;
ROM[1053] <= 32'b00000000011100010010000000100011;
ROM[1054] <= 32'b00000000010000010000000100010011;
ROM[1055] <= 32'b11111111110000010000000100010011;
ROM[1056] <= 32'b00000000000000010010001110000011;
ROM[1057] <= 32'b00000000011100110010001000100011;
ROM[1058] <= 32'b11111111110000010000000100010011;
ROM[1059] <= 32'b00000000000000010010001110000011;
ROM[1060] <= 32'b00000000011100110010000000100011;
ROM[1061] <= 32'b00101000010000000000000011101111;
ROM[1062] <= 32'b00000000000000011010001110000011;
ROM[1063] <= 32'b00000000011100010010000000100011;
ROM[1064] <= 32'b00000000010000010000000100010011;
ROM[1065] <= 32'b00000000000000100010001110000011;
ROM[1066] <= 32'b00000000011100010010000000100011;
ROM[1067] <= 32'b00000000010000010000000100010011;
ROM[1068] <= 32'b11111111110000010000000100010011;
ROM[1069] <= 32'b00000000000000010010001110000011;
ROM[1070] <= 32'b11111111110000010000000100010011;
ROM[1071] <= 32'b00000000000000010010010000000011;
ROM[1072] <= 32'b01000000100000111000001110110011;
ROM[1073] <= 32'b00000000011100010010000000100011;
ROM[1074] <= 32'b00000000010000010000000100010011;
ROM[1075] <= 32'b00000000000100000000001110010011;
ROM[1076] <= 32'b00000000011100010010000000100011;
ROM[1077] <= 32'b00000000010000010000000100010011;
ROM[1078] <= 32'b11111111110000010000000100010011;
ROM[1079] <= 32'b00000000000000010010001110000011;
ROM[1080] <= 32'b11111111110000010000000100010011;
ROM[1081] <= 32'b00000000000000010010010000000011;
ROM[1082] <= 32'b01000000100000111000001110110011;
ROM[1083] <= 32'b00000000011100010010000000100011;
ROM[1084] <= 32'b00000000010000010000000100010011;
ROM[1085] <= 32'b11111111110000010000000100010011;
ROM[1086] <= 32'b00000000000000010010001110000011;
ROM[1087] <= 32'b00000000011100011010001000100011;
ROM[1088] <= 32'b00000000000000011010001110000011;
ROM[1089] <= 32'b00000000011100010010000000100011;
ROM[1090] <= 32'b00000000010000010000000100010011;
ROM[1091] <= 32'b00000001010001101010001110000011;
ROM[1092] <= 32'b00000000011100010010000000100011;
ROM[1093] <= 32'b00000000010000010000000100010011;
ROM[1094] <= 32'b11111111110000010000000100010011;
ROM[1095] <= 32'b00000000000000010010001110000011;
ROM[1096] <= 32'b11111111110000010000000100010011;
ROM[1097] <= 32'b00000000000000010010010000000011;
ROM[1098] <= 32'b00000000100000111000001110110011;
ROM[1099] <= 32'b00000000011100010010000000100011;
ROM[1100] <= 32'b00000000010000010000000100010011;
ROM[1101] <= 32'b11111111110000010000000100010011;
ROM[1102] <= 32'b00000000000000010010001110000011;
ROM[1103] <= 32'b00000000011100110010001000100011;
ROM[1104] <= 32'b00000000000000110010001110000011;
ROM[1105] <= 32'b00000000011100010010000000100011;
ROM[1106] <= 32'b00000000010000010000000100010011;
ROM[1107] <= 32'b00000000010000011010001110000011;
ROM[1108] <= 32'b00000000011100010010000000100011;
ROM[1109] <= 32'b00000000010000010000000100010011;
ROM[1110] <= 32'b00000001010001101010001110000011;
ROM[1111] <= 32'b00000000011100010010000000100011;
ROM[1112] <= 32'b00000000010000010000000100010011;
ROM[1113] <= 32'b11111111110000010000000100010011;
ROM[1114] <= 32'b00000000000000010010001110000011;
ROM[1115] <= 32'b11111111110000010000000100010011;
ROM[1116] <= 32'b00000000000000010010010000000011;
ROM[1117] <= 32'b00000000100000111000001110110011;
ROM[1118] <= 32'b00000000011100010010000000100011;
ROM[1119] <= 32'b00000000010000010000000100010011;
ROM[1120] <= 32'b11111111110000010000000100010011;
ROM[1121] <= 32'b00000000000000010010001110000011;
ROM[1122] <= 32'b00000000011100110010001000100011;
ROM[1123] <= 32'b11111111110000010000000100010011;
ROM[1124] <= 32'b00000000000000010010001110000011;
ROM[1125] <= 32'b00000000011100110010000000100011;
ROM[1126] <= 32'b00000000000000011010001110000011;
ROM[1127] <= 32'b00000000011100010010000000100011;
ROM[1128] <= 32'b00000000010000010000000100010011;
ROM[1129] <= 32'b00000001001101101010001110000011;
ROM[1130] <= 32'b00000000011100010010000000100011;
ROM[1131] <= 32'b00000000010000010000000100010011;
ROM[1132] <= 32'b11111111110000010000000100010011;
ROM[1133] <= 32'b00000000000000010010001110000011;
ROM[1134] <= 32'b11111111110000010000000100010011;
ROM[1135] <= 32'b00000000000000010010010000000011;
ROM[1136] <= 32'b00000000100000111000001110110011;
ROM[1137] <= 32'b00000000011100010010000000100011;
ROM[1138] <= 32'b00000000010000010000000100010011;
ROM[1139] <= 32'b11111111110000010000000100010011;
ROM[1140] <= 32'b00000000000000010010001110000011;
ROM[1141] <= 32'b00000000011100110010001000100011;
ROM[1142] <= 32'b00000000000000110010001110000011;
ROM[1143] <= 32'b00000000011100010010000000100011;
ROM[1144] <= 32'b00000000010000010000000100010011;
ROM[1145] <= 32'b00000000000000100010001110000011;
ROM[1146] <= 32'b00000000011100010010000000100011;
ROM[1147] <= 32'b00000000010000010000000100010011;
ROM[1148] <= 32'b11111111110000010000000100010011;
ROM[1149] <= 32'b00000000000000010010001110000011;
ROM[1150] <= 32'b11111111110000010000000100010011;
ROM[1151] <= 32'b00000000000000010010010000000011;
ROM[1152] <= 32'b01000000100000111000001110110011;
ROM[1153] <= 32'b00000000011100010010000000100011;
ROM[1154] <= 32'b00000000010000010000000100010011;
ROM[1155] <= 32'b00000000000100000000001110010011;
ROM[1156] <= 32'b00000000011100010010000000100011;
ROM[1157] <= 32'b00000000010000010000000100010011;
ROM[1158] <= 32'b11111111110000010000000100010011;
ROM[1159] <= 32'b00000000000000010010001110000011;
ROM[1160] <= 32'b11111111110000010000000100010011;
ROM[1161] <= 32'b00000000000000010010010000000011;
ROM[1162] <= 32'b01000000100000111000001110110011;
ROM[1163] <= 32'b00000000011100010010000000100011;
ROM[1164] <= 32'b00000000010000010000000100010011;
ROM[1165] <= 32'b00000000010000011010001110000011;
ROM[1166] <= 32'b00000000011100010010000000100011;
ROM[1167] <= 32'b00000000010000010000000100010011;
ROM[1168] <= 32'b00000001001101101010001110000011;
ROM[1169] <= 32'b00000000011100010010000000100011;
ROM[1170] <= 32'b00000000010000010000000100010011;
ROM[1171] <= 32'b11111111110000010000000100010011;
ROM[1172] <= 32'b00000000000000010010001110000011;
ROM[1173] <= 32'b11111111110000010000000100010011;
ROM[1174] <= 32'b00000000000000010010010000000011;
ROM[1175] <= 32'b00000000100000111000001110110011;
ROM[1176] <= 32'b00000000011100010010000000100011;
ROM[1177] <= 32'b00000000010000010000000100010011;
ROM[1178] <= 32'b11111111110000010000000100010011;
ROM[1179] <= 32'b00000000000000010010001110000011;
ROM[1180] <= 32'b00000000011100110010001000100011;
ROM[1181] <= 32'b11111111110000010000000100010011;
ROM[1182] <= 32'b00000000000000010010001110000011;
ROM[1183] <= 32'b00000000011100110010000000100011;
ROM[1184] <= 32'b00000000000000100010001110000011;
ROM[1185] <= 32'b00000000011100010010000000100011;
ROM[1186] <= 32'b00000000010000010000000100010011;
ROM[1187] <= 32'b00000000000100000000001110010011;
ROM[1188] <= 32'b00000000011100010010000000100011;
ROM[1189] <= 32'b00000000010000010000000100010011;
ROM[1190] <= 32'b11111111110000010000000100010011;
ROM[1191] <= 32'b00000000000000010010001110000011;
ROM[1192] <= 32'b11111111110000010000000100010011;
ROM[1193] <= 32'b00000000000000010010010000000011;
ROM[1194] <= 32'b00000000100000111000001110110011;
ROM[1195] <= 32'b00000000011100010010000000100011;
ROM[1196] <= 32'b00000000010000010000000100010011;
ROM[1197] <= 32'b00000000100000011010001110000011;
ROM[1198] <= 32'b00000000011100010010000000100011;
ROM[1199] <= 32'b00000000010000010000000100010011;
ROM[1200] <= 32'b00000001010101101010001110000011;
ROM[1201] <= 32'b00000000011100010010000000100011;
ROM[1202] <= 32'b00000000010000010000000100010011;
ROM[1203] <= 32'b11111111110000010000000100010011;
ROM[1204] <= 32'b00000000000000010010001110000011;
ROM[1205] <= 32'b11111111110000010000000100010011;
ROM[1206] <= 32'b00000000000000010010010000000011;
ROM[1207] <= 32'b00000000100000111000001110110011;
ROM[1208] <= 32'b00000000011100010010000000100011;
ROM[1209] <= 32'b00000000010000010000000100010011;
ROM[1210] <= 32'b11111111110000010000000100010011;
ROM[1211] <= 32'b00000000000000010010001110000011;
ROM[1212] <= 32'b00000000011100110010001000100011;
ROM[1213] <= 32'b11111111110000010000000100010011;
ROM[1214] <= 32'b00000000000000010010001110000011;
ROM[1215] <= 32'b00000000011100110010000000100011;
ROM[1216] <= 32'b00000000010000011010001110000011;
ROM[1217] <= 32'b00000000011100010010000000100011;
ROM[1218] <= 32'b00000000010000010000000100010011;
ROM[1219] <= 32'b11111111110000010000000100010011;
ROM[1220] <= 32'b00000000000000010010001110000011;
ROM[1221] <= 32'b00000000011101101010100100100011;
ROM[1222] <= 32'b00000000010000011010001110000011;
ROM[1223] <= 32'b00000000011100010010000000100011;
ROM[1224] <= 32'b00000000010000010000000100010011;
ROM[1225] <= 32'b11111111110000010000000100010011;
ROM[1226] <= 32'b00000000000000010010001110000011;
ROM[1227] <= 32'b00000000011100011010000000100011;
ROM[1228] <= 32'b00000000100000011010001110000011;
ROM[1229] <= 32'b00000000011100010010000000100011;
ROM[1230] <= 32'b00000000010000010000000100010011;
ROM[1231] <= 32'b11111111110000010000000100010011;
ROM[1232] <= 32'b00000000000000010010001110000011;
ROM[1233] <= 32'b00000000011100100010000000100011;
ROM[1234] <= 32'b00000000010000100000000100010011;
ROM[1235] <= 32'b00000001010000000000001110010011;
ROM[1236] <= 32'b01000000011100011000001110110011;
ROM[1237] <= 32'b00000000000000111010000010000011;
ROM[1238] <= 32'b00000000010000111010000110000011;
ROM[1239] <= 32'b00000000100000111010001000000011;
ROM[1240] <= 32'b00000000110000111010001010000011;
ROM[1241] <= 32'b00000001000000111010001100000011;
ROM[1242] <= 32'b00000000000000001000000011100111;
ROM[1243] <= 32'b00000000000000010010000000100011;
ROM[1244] <= 32'b00000000010000010000000100010011;
ROM[1245] <= 32'b00000000000000010010000000100011;
ROM[1246] <= 32'b00000000010000010000000100010011;
ROM[1247] <= 32'b00000000000000010010000000100011;
ROM[1248] <= 32'b00000000010000010000000100010011;
ROM[1249] <= 32'b00000000000000100010001110000011;
ROM[1250] <= 32'b00000000011100010010000000100011;
ROM[1251] <= 32'b00000000010000010000000100010011;
ROM[1252] <= 32'b00000001010101101010001110000011;
ROM[1253] <= 32'b00000000011100010010000000100011;
ROM[1254] <= 32'b00000000010000010000000100010011;
ROM[1255] <= 32'b11111111110000010000000100010011;
ROM[1256] <= 32'b00000000000000010010001110000011;
ROM[1257] <= 32'b11111111110000010000000100010011;
ROM[1258] <= 32'b00000000000000010010010000000011;
ROM[1259] <= 32'b00000000100000111000001110110011;
ROM[1260] <= 32'b00000000011100010010000000100011;
ROM[1261] <= 32'b00000000010000010000000100010011;
ROM[1262] <= 32'b11111111110000010000000100010011;
ROM[1263] <= 32'b00000000000000010010001110000011;
ROM[1264] <= 32'b00000000011100110010001000100011;
ROM[1265] <= 32'b00000000000000110010001110000011;
ROM[1266] <= 32'b00000000011100010010000000100011;
ROM[1267] <= 32'b00000000010000010000000100010011;
ROM[1268] <= 32'b11111111110000010000000100010011;
ROM[1269] <= 32'b00000000000000010010001110000011;
ROM[1270] <= 32'b00000000011100011010010000100011;
ROM[1271] <= 32'b00000000000000100010001110000011;
ROM[1272] <= 32'b00000000011100010010000000100011;
ROM[1273] <= 32'b00000000010000010000000100010011;
ROM[1274] <= 32'b00000000000100000000001110010011;
ROM[1275] <= 32'b00000000011100010010000000100011;
ROM[1276] <= 32'b00000000010000010000000100010011;
ROM[1277] <= 32'b11111111110000010000000100010011;
ROM[1278] <= 32'b00000000000000010010001110000011;
ROM[1279] <= 32'b11111111110000010000000100010011;
ROM[1280] <= 32'b00000000000000010010010000000011;
ROM[1281] <= 32'b00000000100000111000001110110011;
ROM[1282] <= 32'b00000000011100010010000000100011;
ROM[1283] <= 32'b00000000010000010000000100010011;
ROM[1284] <= 32'b11111111110000010000000100010011;
ROM[1285] <= 32'b00000000000000010010001110000011;
ROM[1286] <= 32'b00000000011100100010000000100011;
ROM[1287] <= 32'b00000000000000100010001110000011;
ROM[1288] <= 32'b00000000011100010010000000100011;
ROM[1289] <= 32'b00000000010000010000000100010011;
ROM[1290] <= 32'b00000000000000000001001110110111;
ROM[1291] <= 32'b01000111010000111000001110010011;
ROM[1292] <= 32'b00000000111000111000001110110011;
ROM[1293] <= 32'b00000000011100010010000000100011;
ROM[1294] <= 32'b00000000010000010000000100010011;
ROM[1295] <= 32'b00000000001100010010000000100011;
ROM[1296] <= 32'b00000000010000010000000100010011;
ROM[1297] <= 32'b00000000010000010010000000100011;
ROM[1298] <= 32'b00000000010000010000000100010011;
ROM[1299] <= 32'b00000000010100010010000000100011;
ROM[1300] <= 32'b00000000010000010000000100010011;
ROM[1301] <= 32'b00000000011000010010000000100011;
ROM[1302] <= 32'b00000000010000010000000100010011;
ROM[1303] <= 32'b00000001010000000000001110010011;
ROM[1304] <= 32'b00000000010000111000001110010011;
ROM[1305] <= 32'b01000000011100010000001110110011;
ROM[1306] <= 32'b00000000011100000000001000110011;
ROM[1307] <= 32'b00000000001000000000000110110011;
ROM[1308] <= 32'b01110110000000000000000011101111;
ROM[1309] <= 32'b11111111110000010000000100010011;
ROM[1310] <= 32'b00000000000000010010001110000011;
ROM[1311] <= 32'b00000000011100011010000000100011;
ROM[1312] <= 32'b00000000000000011010001110000011;
ROM[1313] <= 32'b00000000011100010010000000100011;
ROM[1314] <= 32'b00000000010000010000000100010011;
ROM[1315] <= 32'b00000000000000000000001110010011;
ROM[1316] <= 32'b00000000011100010010000000100011;
ROM[1317] <= 32'b00000000010000010000000100010011;
ROM[1318] <= 32'b11111111110000010000000100010011;
ROM[1319] <= 32'b00000000000000010010001110000011;
ROM[1320] <= 32'b11111111110000010000000100010011;
ROM[1321] <= 32'b00000000000000010010010000000011;
ROM[1322] <= 32'b00000000011101000010010010110011;
ROM[1323] <= 32'b00000000100000111010010100110011;
ROM[1324] <= 32'b00000000101001001000001110110011;
ROM[1325] <= 32'b00000000000100111000001110010011;
ROM[1326] <= 32'b00000000000100111111001110010011;
ROM[1327] <= 32'b00000000011100010010000000100011;
ROM[1328] <= 32'b00000000010000010000000100010011;
ROM[1329] <= 32'b11111111110000010000000100010011;
ROM[1330] <= 32'b00000000000000010010001110000011;
ROM[1331] <= 32'b00000000000000111000101001100011;
ROM[1332] <= 32'b00000000000000000001001110110111;
ROM[1333] <= 32'b01111101000000111000001110010011;
ROM[1334] <= 32'b00000000111000111000001110110011;
ROM[1335] <= 32'b00000000000000111000000011100111;
ROM[1336] <= 32'b00000000000000011010001110000011;
ROM[1337] <= 32'b00000000011100010010000000100011;
ROM[1338] <= 32'b00000000010000010000000100010011;
ROM[1339] <= 32'b00000000000000011010001110000011;
ROM[1340] <= 32'b00000000011100010010000000100011;
ROM[1341] <= 32'b00000000010000010000000100010011;
ROM[1342] <= 32'b00000001001101101010001110000011;
ROM[1343] <= 32'b00000000011100010010000000100011;
ROM[1344] <= 32'b00000000010000010000000100010011;
ROM[1345] <= 32'b11111111110000010000000100010011;
ROM[1346] <= 32'b00000000000000010010001110000011;
ROM[1347] <= 32'b11111111110000010000000100010011;
ROM[1348] <= 32'b00000000000000010010010000000011;
ROM[1349] <= 32'b00000000100000111000001110110011;
ROM[1350] <= 32'b00000000011100010010000000100011;
ROM[1351] <= 32'b00000000010000010000000100010011;
ROM[1352] <= 32'b11111111110000010000000100010011;
ROM[1353] <= 32'b00000000000000010010001110000011;
ROM[1354] <= 32'b00000000011100110010001000100011;
ROM[1355] <= 32'b00000000000000110010001110000011;
ROM[1356] <= 32'b00000000011100010010000000100011;
ROM[1357] <= 32'b00000000010000010000000100010011;
ROM[1358] <= 32'b11111111110000010000000100010011;
ROM[1359] <= 32'b00000000000000010010001110000011;
ROM[1360] <= 32'b11111111110000010000000100010011;
ROM[1361] <= 32'b00000000000000010010010000000011;
ROM[1362] <= 32'b01000000100000111000001110110011;
ROM[1363] <= 32'b00000000011100010010000000100011;
ROM[1364] <= 32'b00000000010000010000000100010011;
ROM[1365] <= 32'b00000000000000100010001110000011;
ROM[1366] <= 32'b00000000011100010010000000100011;
ROM[1367] <= 32'b00000000010000010000000100010011;
ROM[1368] <= 32'b11111111110000010000000100010011;
ROM[1369] <= 32'b00000000000000010010001110000011;
ROM[1370] <= 32'b11111111110000010000000100010011;
ROM[1371] <= 32'b00000000000000010010010000000011;
ROM[1372] <= 32'b00000000011101000010010010110011;
ROM[1373] <= 32'b00000000100000111010010100110011;
ROM[1374] <= 32'b00000000101001001000001110110011;
ROM[1375] <= 32'b00000000000100111000001110010011;
ROM[1376] <= 32'b00000000000100111111001110010011;
ROM[1377] <= 32'b00000000011100010010000000100011;
ROM[1378] <= 32'b00000000010000010000000100010011;
ROM[1379] <= 32'b11111111110000010000000100010011;
ROM[1380] <= 32'b00000000000000010010001110000011;
ROM[1381] <= 32'b00000000000000111000101001100011;
ROM[1382] <= 32'b00000000000000000001001110110111;
ROM[1383] <= 32'b01101111010000111000001110010011;
ROM[1384] <= 32'b00000000111000111000001110110011;
ROM[1385] <= 32'b00000000000000111000000011100111;
ROM[1386] <= 32'b00000000100000011010001110000011;
ROM[1387] <= 32'b00000000011100010010000000100011;
ROM[1388] <= 32'b00000000010000010000000100010011;
ROM[1389] <= 32'b00000000000000100010001110000011;
ROM[1390] <= 32'b00000000011100010010000000100011;
ROM[1391] <= 32'b00000000010000010000000100010011;
ROM[1392] <= 32'b00000001001101101010001110000011;
ROM[1393] <= 32'b00000000011100010010000000100011;
ROM[1394] <= 32'b00000000010000010000000100010011;
ROM[1395] <= 32'b11111111110000010000000100010011;
ROM[1396] <= 32'b00000000000000010010001110000011;
ROM[1397] <= 32'b11111111110000010000000100010011;
ROM[1398] <= 32'b00000000000000010010010000000011;
ROM[1399] <= 32'b00000000100000111000001110110011;
ROM[1400] <= 32'b00000000011100010010000000100011;
ROM[1401] <= 32'b00000000010000010000000100010011;
ROM[1402] <= 32'b11111111110000010000000100010011;
ROM[1403] <= 32'b00000000000000010010001110000011;
ROM[1404] <= 32'b00000000011100110010001000100011;
ROM[1405] <= 32'b11111111110000010000000100010011;
ROM[1406] <= 32'b00000000000000010010001110000011;
ROM[1407] <= 32'b00000000011100110010000000100011;
ROM[1408] <= 32'b00000000000000011010001110000011;
ROM[1409] <= 32'b00000000011100010010000000100011;
ROM[1410] <= 32'b00000000010000010000000100010011;
ROM[1411] <= 32'b00000001010001101010001110000011;
ROM[1412] <= 32'b00000000011100010010000000100011;
ROM[1413] <= 32'b00000000010000010000000100010011;
ROM[1414] <= 32'b11111111110000010000000100010011;
ROM[1415] <= 32'b00000000000000010010001110000011;
ROM[1416] <= 32'b11111111110000010000000100010011;
ROM[1417] <= 32'b00000000000000010010010000000011;
ROM[1418] <= 32'b00000000100000111000001110110011;
ROM[1419] <= 32'b00000000011100010010000000100011;
ROM[1420] <= 32'b00000000010000010000000100010011;
ROM[1421] <= 32'b11111111110000010000000100010011;
ROM[1422] <= 32'b00000000000000010010001110000011;
ROM[1423] <= 32'b00000000011100110010001000100011;
ROM[1424] <= 32'b00000000000000110010001110000011;
ROM[1425] <= 32'b00000000011100010010000000100011;
ROM[1426] <= 32'b00000000010000010000000100010011;
ROM[1427] <= 32'b00000000000000100010001110000011;
ROM[1428] <= 32'b00000000011100010010000000100011;
ROM[1429] <= 32'b00000000010000010000000100010011;
ROM[1430] <= 32'b00000001010001101010001110000011;
ROM[1431] <= 32'b00000000011100010010000000100011;
ROM[1432] <= 32'b00000000010000010000000100010011;
ROM[1433] <= 32'b11111111110000010000000100010011;
ROM[1434] <= 32'b00000000000000010010001110000011;
ROM[1435] <= 32'b11111111110000010000000100010011;
ROM[1436] <= 32'b00000000000000010010010000000011;
ROM[1437] <= 32'b00000000100000111000001110110011;
ROM[1438] <= 32'b00000000011100010010000000100011;
ROM[1439] <= 32'b00000000010000010000000100010011;
ROM[1440] <= 32'b11111111110000010000000100010011;
ROM[1441] <= 32'b00000000000000010010001110000011;
ROM[1442] <= 32'b00000000011100110010001000100011;
ROM[1443] <= 32'b11111111110000010000000100010011;
ROM[1444] <= 32'b00000000000000010010001110000011;
ROM[1445] <= 32'b00000000011100110010000000100011;
ROM[1446] <= 32'b00000000000000100010001110000011;
ROM[1447] <= 32'b00000000011100010010000000100011;
ROM[1448] <= 32'b00000000010000010000000100010011;
ROM[1449] <= 32'b00000000000000011010001110000011;
ROM[1450] <= 32'b00000000011100010010000000100011;
ROM[1451] <= 32'b00000000010000010000000100010011;
ROM[1452] <= 32'b00000001010001101010001110000011;
ROM[1453] <= 32'b00000000011100010010000000100011;
ROM[1454] <= 32'b00000000010000010000000100010011;
ROM[1455] <= 32'b11111111110000010000000100010011;
ROM[1456] <= 32'b00000000000000010010001110000011;
ROM[1457] <= 32'b11111111110000010000000100010011;
ROM[1458] <= 32'b00000000000000010010010000000011;
ROM[1459] <= 32'b00000000100000111000001110110011;
ROM[1460] <= 32'b00000000011100010010000000100011;
ROM[1461] <= 32'b00000000010000010000000100010011;
ROM[1462] <= 32'b11111111110000010000000100010011;
ROM[1463] <= 32'b00000000000000010010001110000011;
ROM[1464] <= 32'b00000000011100110010001000100011;
ROM[1465] <= 32'b11111111110000010000000100010011;
ROM[1466] <= 32'b00000000000000010010001110000011;
ROM[1467] <= 32'b00000000011100110010000000100011;
ROM[1468] <= 32'b00001101110000000000000011101111;
ROM[1469] <= 32'b00000000000000011010001110000011;
ROM[1470] <= 32'b00000000011100010010000000100011;
ROM[1471] <= 32'b00000000010000010000000100010011;
ROM[1472] <= 32'b00000001001101101010001110000011;
ROM[1473] <= 32'b00000000011100010010000000100011;
ROM[1474] <= 32'b00000000010000010000000100010011;
ROM[1475] <= 32'b11111111110000010000000100010011;
ROM[1476] <= 32'b00000000000000010010001110000011;
ROM[1477] <= 32'b11111111110000010000000100010011;
ROM[1478] <= 32'b00000000000000010010010000000011;
ROM[1479] <= 32'b00000000100000111000001110110011;
ROM[1480] <= 32'b00000000011100010010000000100011;
ROM[1481] <= 32'b00000000010000010000000100010011;
ROM[1482] <= 32'b11111111110000010000000100010011;
ROM[1483] <= 32'b00000000000000010010001110000011;
ROM[1484] <= 32'b00000000011100110010001000100011;
ROM[1485] <= 32'b00000000000000110010001110000011;
ROM[1486] <= 32'b00000000011100010010000000100011;
ROM[1487] <= 32'b00000000010000010000000100010011;
ROM[1488] <= 32'b00000000100000011010001110000011;
ROM[1489] <= 32'b00000000011100010010000000100011;
ROM[1490] <= 32'b00000000010000010000000100010011;
ROM[1491] <= 32'b11111111110000010000000100010011;
ROM[1492] <= 32'b00000000000000010010001110000011;
ROM[1493] <= 32'b11111111110000010000000100010011;
ROM[1494] <= 32'b00000000000000010010010000000011;
ROM[1495] <= 32'b00000000100000111000001110110011;
ROM[1496] <= 32'b00000000011100010010000000100011;
ROM[1497] <= 32'b00000000010000010000000100010011;
ROM[1498] <= 32'b00000000000000011010001110000011;
ROM[1499] <= 32'b00000000011100010010000000100011;
ROM[1500] <= 32'b00000000010000010000000100010011;
ROM[1501] <= 32'b00000001001101101010001110000011;
ROM[1502] <= 32'b00000000011100010010000000100011;
ROM[1503] <= 32'b00000000010000010000000100010011;
ROM[1504] <= 32'b11111111110000010000000100010011;
ROM[1505] <= 32'b00000000000000010010001110000011;
ROM[1506] <= 32'b11111111110000010000000100010011;
ROM[1507] <= 32'b00000000000000010010010000000011;
ROM[1508] <= 32'b00000000100000111000001110110011;
ROM[1509] <= 32'b00000000011100010010000000100011;
ROM[1510] <= 32'b00000000010000010000000100010011;
ROM[1511] <= 32'b11111111110000010000000100010011;
ROM[1512] <= 32'b00000000000000010010001110000011;
ROM[1513] <= 32'b00000000011100110010001000100011;
ROM[1514] <= 32'b11111111110000010000000100010011;
ROM[1515] <= 32'b00000000000000010010001110000011;
ROM[1516] <= 32'b00000000011100110010000000100011;
ROM[1517] <= 32'b00000000000000011010001110000011;
ROM[1518] <= 32'b00000000011100010010000000100011;
ROM[1519] <= 32'b00000000010000010000000100010011;
ROM[1520] <= 32'b11111111110000010000000100010011;
ROM[1521] <= 32'b00000000000000010010001110000011;
ROM[1522] <= 32'b00000000011100100010000000100011;
ROM[1523] <= 32'b00001100110000000000000011101111;
ROM[1524] <= 32'b00000000100000011010001110000011;
ROM[1525] <= 32'b00000000011100010010000000100011;
ROM[1526] <= 32'b00000000010000010000000100010011;
ROM[1527] <= 32'b00000000000000100010001110000011;
ROM[1528] <= 32'b00000000011100010010000000100011;
ROM[1529] <= 32'b00000000010000010000000100010011;
ROM[1530] <= 32'b00000001001101101010001110000011;
ROM[1531] <= 32'b00000000011100010010000000100011;
ROM[1532] <= 32'b00000000010000010000000100010011;
ROM[1533] <= 32'b11111111110000010000000100010011;
ROM[1534] <= 32'b00000000000000010010001110000011;
ROM[1535] <= 32'b11111111110000010000000100010011;
ROM[1536] <= 32'b00000000000000010010010000000011;
ROM[1537] <= 32'b00000000100000111000001110110011;
ROM[1538] <= 32'b00000000011100010010000000100011;
ROM[1539] <= 32'b00000000010000010000000100010011;
ROM[1540] <= 32'b11111111110000010000000100010011;
ROM[1541] <= 32'b00000000000000010010001110000011;
ROM[1542] <= 32'b00000000011100110010001000100011;
ROM[1543] <= 32'b11111111110000010000000100010011;
ROM[1544] <= 32'b00000000000000010010001110000011;
ROM[1545] <= 32'b00000000011100110010000000100011;
ROM[1546] <= 32'b00000001001001101010001110000011;
ROM[1547] <= 32'b00000000011100010010000000100011;
ROM[1548] <= 32'b00000000010000010000000100010011;
ROM[1549] <= 32'b00000000000000100010001110000011;
ROM[1550] <= 32'b00000000011100010010000000100011;
ROM[1551] <= 32'b00000000010000010000000100010011;
ROM[1552] <= 32'b00000001010001101010001110000011;
ROM[1553] <= 32'b00000000011100010010000000100011;
ROM[1554] <= 32'b00000000010000010000000100010011;
ROM[1555] <= 32'b11111111110000010000000100010011;
ROM[1556] <= 32'b00000000000000010010001110000011;
ROM[1557] <= 32'b11111111110000010000000100010011;
ROM[1558] <= 32'b00000000000000010010010000000011;
ROM[1559] <= 32'b00000000100000111000001110110011;
ROM[1560] <= 32'b00000000011100010010000000100011;
ROM[1561] <= 32'b00000000010000010000000100010011;
ROM[1562] <= 32'b11111111110000010000000100010011;
ROM[1563] <= 32'b00000000000000010010001110000011;
ROM[1564] <= 32'b00000000011100110010001000100011;
ROM[1565] <= 32'b11111111110000010000000100010011;
ROM[1566] <= 32'b00000000000000010010001110000011;
ROM[1567] <= 32'b00000000011100110010000000100011;
ROM[1568] <= 32'b00000000000000100010001110000011;
ROM[1569] <= 32'b00000000011100010010000000100011;
ROM[1570] <= 32'b00000000010000010000000100010011;
ROM[1571] <= 32'b11111111110000010000000100010011;
ROM[1572] <= 32'b00000000000000010010001110000011;
ROM[1573] <= 32'b00000000011101101010100100100011;
ROM[1574] <= 32'b00000000000000100010001110000011;
ROM[1575] <= 32'b00000000011100010010000000100011;
ROM[1576] <= 32'b00000000010000010000000100010011;
ROM[1577] <= 32'b00000000000000100010001110000011;
ROM[1578] <= 32'b00000000011100010010000000100011;
ROM[1579] <= 32'b00000000010000010000000100010011;
ROM[1580] <= 32'b00000001001101101010001110000011;
ROM[1581] <= 32'b00000000011100010010000000100011;
ROM[1582] <= 32'b00000000010000010000000100010011;
ROM[1583] <= 32'b11111111110000010000000100010011;
ROM[1584] <= 32'b00000000000000010010001110000011;
ROM[1585] <= 32'b11111111110000010000000100010011;
ROM[1586] <= 32'b00000000000000010010010000000011;
ROM[1587] <= 32'b00000000100000111000001110110011;
ROM[1588] <= 32'b00000000011100010010000000100011;
ROM[1589] <= 32'b00000000010000010000000100010011;
ROM[1590] <= 32'b11111111110000010000000100010011;
ROM[1591] <= 32'b00000000000000010010001110000011;
ROM[1592] <= 32'b00000000011100110010001000100011;
ROM[1593] <= 32'b00000000000000110010001110000011;
ROM[1594] <= 32'b00000000011100010010000000100011;
ROM[1595] <= 32'b00000000010000010000000100010011;
ROM[1596] <= 32'b11111111110000010000000100010011;
ROM[1597] <= 32'b00000000000000010010001110000011;
ROM[1598] <= 32'b11111111110000010000000100010011;
ROM[1599] <= 32'b00000000000000010010010000000011;
ROM[1600] <= 32'b01000000100000111000001110110011;
ROM[1601] <= 32'b00000000011100010010000000100011;
ROM[1602] <= 32'b00000000010000010000000100010011;
ROM[1603] <= 32'b00000000000000100010001110000011;
ROM[1604] <= 32'b00000000011100010010000000100011;
ROM[1605] <= 32'b00000000010000010000000100010011;
ROM[1606] <= 32'b00000001010001101010001110000011;
ROM[1607] <= 32'b00000000011100010010000000100011;
ROM[1608] <= 32'b00000000010000010000000100010011;
ROM[1609] <= 32'b11111111110000010000000100010011;
ROM[1610] <= 32'b00000000000000010010001110000011;
ROM[1611] <= 32'b11111111110000010000000100010011;
ROM[1612] <= 32'b00000000000000010010010000000011;
ROM[1613] <= 32'b00000000100000111000001110110011;
ROM[1614] <= 32'b00000000011100010010000000100011;
ROM[1615] <= 32'b00000000010000010000000100010011;
ROM[1616] <= 32'b11111111110000010000000100010011;
ROM[1617] <= 32'b00000000000000010010001110000011;
ROM[1618] <= 32'b00000000011100110010001000100011;
ROM[1619] <= 32'b00000000000000110010001110000011;
ROM[1620] <= 32'b00000000011100010010000000100011;
ROM[1621] <= 32'b00000000010000010000000100010011;
ROM[1622] <= 32'b11111111110000010000000100010011;
ROM[1623] <= 32'b00000000000000010010001110000011;
ROM[1624] <= 32'b11111111110000010000000100010011;
ROM[1625] <= 32'b00000000000000010010010000000011;
ROM[1626] <= 32'b00000000011101000010010010110011;
ROM[1627] <= 32'b00000000100000111010010100110011;
ROM[1628] <= 32'b00000000101001001000001110110011;
ROM[1629] <= 32'b00000000000100111000001110010011;
ROM[1630] <= 32'b00000000000100111111001110010011;
ROM[1631] <= 32'b00000000011100010010000000100011;
ROM[1632] <= 32'b00000000010000010000000100010011;
ROM[1633] <= 32'b11111111110000010000000100010011;
ROM[1634] <= 32'b00000000000000010010001110000011;
ROM[1635] <= 32'b00000000000000111000101001100011;
ROM[1636] <= 32'b00000000000000000001001110110111;
ROM[1637] <= 32'b10011010010000111000001110010011;
ROM[1638] <= 32'b00000000111000111000001110110011;
ROM[1639] <= 32'b00000000000000111000000011100111;
ROM[1640] <= 32'b00011111010000000000000011101111;
ROM[1641] <= 32'b00000000000000100010001110000011;
ROM[1642] <= 32'b00000000011100010010000000100011;
ROM[1643] <= 32'b00000000010000010000000100010011;
ROM[1644] <= 32'b00000001010001101010001110000011;
ROM[1645] <= 32'b00000000011100010010000000100011;
ROM[1646] <= 32'b00000000010000010000000100010011;
ROM[1647] <= 32'b11111111110000010000000100010011;
ROM[1648] <= 32'b00000000000000010010001110000011;
ROM[1649] <= 32'b11111111110000010000000100010011;
ROM[1650] <= 32'b00000000000000010010010000000011;
ROM[1651] <= 32'b00000000100000111000001110110011;
ROM[1652] <= 32'b00000000011100010010000000100011;
ROM[1653] <= 32'b00000000010000010000000100010011;
ROM[1654] <= 32'b11111111110000010000000100010011;
ROM[1655] <= 32'b00000000000000010010001110000011;
ROM[1656] <= 32'b00000000011100110010001000100011;
ROM[1657] <= 32'b00000000000000110010001110000011;
ROM[1658] <= 32'b00000000011100010010000000100011;
ROM[1659] <= 32'b00000000010000010000000100010011;
ROM[1660] <= 32'b11111111110000010000000100010011;
ROM[1661] <= 32'b00000000000000010010001110000011;
ROM[1662] <= 32'b00000000011100011010001000100011;
ROM[1663] <= 32'b00000000000000100010001110000011;
ROM[1664] <= 32'b00000000011100010010000000100011;
ROM[1665] <= 32'b00000000010000010000000100010011;
ROM[1666] <= 32'b00000001001101101010001110000011;
ROM[1667] <= 32'b00000000011100010010000000100011;
ROM[1668] <= 32'b00000000010000010000000100010011;
ROM[1669] <= 32'b11111111110000010000000100010011;
ROM[1670] <= 32'b00000000000000010010001110000011;
ROM[1671] <= 32'b11111111110000010000000100010011;
ROM[1672] <= 32'b00000000000000010010010000000011;
ROM[1673] <= 32'b00000000100000111000001110110011;
ROM[1674] <= 32'b00000000011100010010000000100011;
ROM[1675] <= 32'b00000000010000010000000100010011;
ROM[1676] <= 32'b11111111110000010000000100010011;
ROM[1677] <= 32'b00000000000000010010001110000011;
ROM[1678] <= 32'b00000000011100110010001000100011;
ROM[1679] <= 32'b00000000000000110010001110000011;
ROM[1680] <= 32'b00000000011100010010000000100011;
ROM[1681] <= 32'b00000000010000010000000100010011;
ROM[1682] <= 32'b00000000010000011010001110000011;
ROM[1683] <= 32'b00000000011100010010000000100011;
ROM[1684] <= 32'b00000000010000010000000100010011;
ROM[1685] <= 32'b00000001001101101010001110000011;
ROM[1686] <= 32'b00000000011100010010000000100011;
ROM[1687] <= 32'b00000000010000010000000100010011;
ROM[1688] <= 32'b11111111110000010000000100010011;
ROM[1689] <= 32'b00000000000000010010001110000011;
ROM[1690] <= 32'b11111111110000010000000100010011;
ROM[1691] <= 32'b00000000000000010010010000000011;
ROM[1692] <= 32'b00000000100000111000001110110011;
ROM[1693] <= 32'b00000000011100010010000000100011;
ROM[1694] <= 32'b00000000010000010000000100010011;
ROM[1695] <= 32'b11111111110000010000000100010011;
ROM[1696] <= 32'b00000000000000010010001110000011;
ROM[1697] <= 32'b00000000011100110010001000100011;
ROM[1698] <= 32'b00000000000000110010001110000011;
ROM[1699] <= 32'b00000000011100010010000000100011;
ROM[1700] <= 32'b00000000010000010000000100010011;
ROM[1701] <= 32'b11111111110000010000000100010011;
ROM[1702] <= 32'b00000000000000010010001110000011;
ROM[1703] <= 32'b11111111110000010000000100010011;
ROM[1704] <= 32'b00000000000000010010010000000011;
ROM[1705] <= 32'b00000000100000111000001110110011;
ROM[1706] <= 32'b00000000011100010010000000100011;
ROM[1707] <= 32'b00000000010000010000000100010011;
ROM[1708] <= 32'b00000000000000100010001110000011;
ROM[1709] <= 32'b00000000011100010010000000100011;
ROM[1710] <= 32'b00000000010000010000000100010011;
ROM[1711] <= 32'b00000001001101101010001110000011;
ROM[1712] <= 32'b00000000011100010010000000100011;
ROM[1713] <= 32'b00000000010000010000000100010011;
ROM[1714] <= 32'b11111111110000010000000100010011;
ROM[1715] <= 32'b00000000000000010010001110000011;
ROM[1716] <= 32'b11111111110000010000000100010011;
ROM[1717] <= 32'b00000000000000010010010000000011;
ROM[1718] <= 32'b00000000100000111000001110110011;
ROM[1719] <= 32'b00000000011100010010000000100011;
ROM[1720] <= 32'b00000000010000010000000100010011;
ROM[1721] <= 32'b11111111110000010000000100010011;
ROM[1722] <= 32'b00000000000000010010001110000011;
ROM[1723] <= 32'b00000000011100110010001000100011;
ROM[1724] <= 32'b11111111110000010000000100010011;
ROM[1725] <= 32'b00000000000000010010001110000011;
ROM[1726] <= 32'b00000000011100110010000000100011;
ROM[1727] <= 32'b00000000010000011010001110000011;
ROM[1728] <= 32'b00000000011100010010000000100011;
ROM[1729] <= 32'b00000000010000010000000100010011;
ROM[1730] <= 32'b00000001010001101010001110000011;
ROM[1731] <= 32'b00000000011100010010000000100011;
ROM[1732] <= 32'b00000000010000010000000100010011;
ROM[1733] <= 32'b11111111110000010000000100010011;
ROM[1734] <= 32'b00000000000000010010001110000011;
ROM[1735] <= 32'b11111111110000010000000100010011;
ROM[1736] <= 32'b00000000000000010010010000000011;
ROM[1737] <= 32'b00000000100000111000001110110011;
ROM[1738] <= 32'b00000000011100010010000000100011;
ROM[1739] <= 32'b00000000010000010000000100010011;
ROM[1740] <= 32'b11111111110000010000000100010011;
ROM[1741] <= 32'b00000000000000010010001110000011;
ROM[1742] <= 32'b00000000011100110010001000100011;
ROM[1743] <= 32'b00000000000000110010001110000011;
ROM[1744] <= 32'b00000000011100010010000000100011;
ROM[1745] <= 32'b00000000010000010000000100010011;
ROM[1746] <= 32'b00000000000000100010001110000011;
ROM[1747] <= 32'b00000000011100010010000000100011;
ROM[1748] <= 32'b00000000010000010000000100010011;
ROM[1749] <= 32'b00000001010001101010001110000011;
ROM[1750] <= 32'b00000000011100010010000000100011;
ROM[1751] <= 32'b00000000010000010000000100010011;
ROM[1752] <= 32'b11111111110000010000000100010011;
ROM[1753] <= 32'b00000000000000010010001110000011;
ROM[1754] <= 32'b11111111110000010000000100010011;
ROM[1755] <= 32'b00000000000000010010010000000011;
ROM[1756] <= 32'b00000000100000111000001110110011;
ROM[1757] <= 32'b00000000011100010010000000100011;
ROM[1758] <= 32'b00000000010000010000000100010011;
ROM[1759] <= 32'b11111111110000010000000100010011;
ROM[1760] <= 32'b00000000000000010010001110000011;
ROM[1761] <= 32'b00000000011100110010001000100011;
ROM[1762] <= 32'b11111111110000010000000100010011;
ROM[1763] <= 32'b00000000000000010010001110000011;
ROM[1764] <= 32'b00000000011100110010000000100011;
ROM[1765] <= 32'b00000000000000000000001110010011;
ROM[1766] <= 32'b00000000011100010010000000100011;
ROM[1767] <= 32'b00000000010000010000000100010011;
ROM[1768] <= 32'b11111111110000010000000100010011;
ROM[1769] <= 32'b00000000000000010010001110000011;
ROM[1770] <= 32'b00000000011100100010000000100011;
ROM[1771] <= 32'b00000000010000100000000100010011;
ROM[1772] <= 32'b00000001010000000000001110010011;
ROM[1773] <= 32'b01000000011100011000001110110011;
ROM[1774] <= 32'b00000000000000111010000010000011;
ROM[1775] <= 32'b00000000010000111010000110000011;
ROM[1776] <= 32'b00000000100000111010001000000011;
ROM[1777] <= 32'b00000000110000111010001010000011;
ROM[1778] <= 32'b00000001000000111010001100000011;
ROM[1779] <= 32'b00000000000000001000000011100111;
ROM[1780] <= 32'b00000000000000010010000000100011;
ROM[1781] <= 32'b00000000010000010000000100010011;
ROM[1782] <= 32'b00000001001001101010001110000011;
ROM[1783] <= 32'b00000000011100010010000000100011;
ROM[1784] <= 32'b00000000010000010000000100010011;
ROM[1785] <= 32'b00000000000000100010001110000011;
ROM[1786] <= 32'b00000000011100010010000000100011;
ROM[1787] <= 32'b00000000010000010000000100010011;
ROM[1788] <= 32'b11111111110000010000000100010011;
ROM[1789] <= 32'b00000000000000010010001110000011;
ROM[1790] <= 32'b11111111110000010000000100010011;
ROM[1791] <= 32'b00000000000000010010010000000011;
ROM[1792] <= 32'b00000000011101000010001110110011;
ROM[1793] <= 32'b00000000011100010010000000100011;
ROM[1794] <= 32'b00000000010000010000000100010011;
ROM[1795] <= 32'b11111111110000010000000100010011;
ROM[1796] <= 32'b00000000000000010010001110000011;
ROM[1797] <= 32'b00000000000000111000101001100011;
ROM[1798] <= 32'b00000000000000000001001110110111;
ROM[1799] <= 32'b11000010110000111000001110010011;
ROM[1800] <= 32'b00000000111000111000001110110011;
ROM[1801] <= 32'b00000000000000111000000011100111;
ROM[1802] <= 32'b00000100000000000000000011101111;
ROM[1803] <= 32'b00000000000000000000001110010011;
ROM[1804] <= 32'b00000000011100010010000000100011;
ROM[1805] <= 32'b00000000010000010000000100010011;
ROM[1806] <= 32'b11111111110000010000000100010011;
ROM[1807] <= 32'b00000000000000010010001110000011;
ROM[1808] <= 32'b00000000011100100010000000100011;
ROM[1809] <= 32'b00000000010000100000000100010011;
ROM[1810] <= 32'b00000001010000000000001110010011;
ROM[1811] <= 32'b01000000011100011000001110110011;
ROM[1812] <= 32'b00000000000000111010000010000011;
ROM[1813] <= 32'b00000000010000111010000110000011;
ROM[1814] <= 32'b00000000100000111010001000000011;
ROM[1815] <= 32'b00000000110000111010001010000011;
ROM[1816] <= 32'b00000001000000111010001100000011;
ROM[1817] <= 32'b00000000000000001000000011100111;
ROM[1818] <= 32'b00000001001001101010001110000011;
ROM[1819] <= 32'b00000000011100010010000000100011;
ROM[1820] <= 32'b00000000010000010000000100010011;
ROM[1821] <= 32'b11111111110000010000000100010011;
ROM[1822] <= 32'b00000000000000010010001110000011;
ROM[1823] <= 32'b00000000011100011010000000100011;
ROM[1824] <= 32'b00000000000000011010001110000011;
ROM[1825] <= 32'b00000000011100010010000000100011;
ROM[1826] <= 32'b00000000010000010000000100010011;
ROM[1827] <= 32'b00000001010001101010001110000011;
ROM[1828] <= 32'b00000000011100010010000000100011;
ROM[1829] <= 32'b00000000010000010000000100010011;
ROM[1830] <= 32'b11111111110000010000000100010011;
ROM[1831] <= 32'b00000000000000010010001110000011;
ROM[1832] <= 32'b11111111110000010000000100010011;
ROM[1833] <= 32'b00000000000000010010010000000011;
ROM[1834] <= 32'b00000000100000111000001110110011;
ROM[1835] <= 32'b00000000011100010010000000100011;
ROM[1836] <= 32'b00000000010000010000000100010011;
ROM[1837] <= 32'b11111111110000010000000100010011;
ROM[1838] <= 32'b00000000000000010010001110000011;
ROM[1839] <= 32'b00000000011100110010001000100011;
ROM[1840] <= 32'b00000000000000110010001110000011;
ROM[1841] <= 32'b00000000011100010010000000100011;
ROM[1842] <= 32'b00000000010000010000000100010011;
ROM[1843] <= 32'b00000000000000000000001110010011;
ROM[1844] <= 32'b00000000011100010010000000100011;
ROM[1845] <= 32'b00000000010000010000000100010011;
ROM[1846] <= 32'b11111111110000010000000100010011;
ROM[1847] <= 32'b00000000000000010010001110000011;
ROM[1848] <= 32'b11111111110000010000000100010011;
ROM[1849] <= 32'b00000000000000010010010000000011;
ROM[1850] <= 32'b00000000011101000010010010110011;
ROM[1851] <= 32'b00000000100000111010010100110011;
ROM[1852] <= 32'b00000000101001001000001110110011;
ROM[1853] <= 32'b00000000000100111000001110010011;
ROM[1854] <= 32'b00000000000100111111001110010011;
ROM[1855] <= 32'b00000000011100010010000000100011;
ROM[1856] <= 32'b00000000010000010000000100010011;
ROM[1857] <= 32'b11111111110000010000000100010011;
ROM[1858] <= 32'b00000000000000010010001110000011;
ROM[1859] <= 32'b01000000011100000000001110110011;
ROM[1860] <= 32'b00000000000100111000001110010011;
ROM[1861] <= 32'b00000000011100010010000000100011;
ROM[1862] <= 32'b00000000010000010000000100010011;
ROM[1863] <= 32'b00000000000000011010001110000011;
ROM[1864] <= 32'b00000000011100010010000000100011;
ROM[1865] <= 32'b00000000010000010000000100010011;
ROM[1866] <= 32'b00000001010001101010001110000011;
ROM[1867] <= 32'b00000000011100010010000000100011;
ROM[1868] <= 32'b00000000010000010000000100010011;
ROM[1869] <= 32'b11111111110000010000000100010011;
ROM[1870] <= 32'b00000000000000010010001110000011;
ROM[1871] <= 32'b11111111110000010000000100010011;
ROM[1872] <= 32'b00000000000000010010010000000011;
ROM[1873] <= 32'b00000000100000111000001110110011;
ROM[1874] <= 32'b00000000011100010010000000100011;
ROM[1875] <= 32'b00000000010000010000000100010011;
ROM[1876] <= 32'b11111111110000010000000100010011;
ROM[1877] <= 32'b00000000000000010010001110000011;
ROM[1878] <= 32'b00000000011100110010001000100011;
ROM[1879] <= 32'b00000000000000110010001110000011;
ROM[1880] <= 32'b00000000011100010010000000100011;
ROM[1881] <= 32'b00000000010000010000000100010011;
ROM[1882] <= 32'b00000000000000100010001110000011;
ROM[1883] <= 32'b00000000011100010010000000100011;
ROM[1884] <= 32'b00000000010000010000000100010011;
ROM[1885] <= 32'b11111111110000010000000100010011;
ROM[1886] <= 32'b00000000000000010010001110000011;
ROM[1887] <= 32'b11111111110000010000000100010011;
ROM[1888] <= 32'b00000000000000010010010000000011;
ROM[1889] <= 32'b00000000100000111010001110110011;
ROM[1890] <= 32'b00000000011100010010000000100011;
ROM[1891] <= 32'b00000000010000010000000100010011;
ROM[1892] <= 32'b11111111110000010000000100010011;
ROM[1893] <= 32'b00000000000000010010001110000011;
ROM[1894] <= 32'b11111111110000010000000100010011;
ROM[1895] <= 32'b00000000000000010010010000000011;
ROM[1896] <= 32'b00000000100000111111001110110011;
ROM[1897] <= 32'b00000000011100010010000000100011;
ROM[1898] <= 32'b00000000010000010000000100010011;
ROM[1899] <= 32'b11111111110000010000000100010011;
ROM[1900] <= 32'b00000000000000010010001110000011;
ROM[1901] <= 32'b01000000011100000000001110110011;
ROM[1902] <= 32'b00000000000100111000001110010011;
ROM[1903] <= 32'b00000000011100010010000000100011;
ROM[1904] <= 32'b00000000010000010000000100010011;
ROM[1905] <= 32'b11111111110000010000000100010011;
ROM[1906] <= 32'b00000000000000010010001110000011;
ROM[1907] <= 32'b00000000000000111000101001100011;
ROM[1908] <= 32'b00000000000000000001001110110111;
ROM[1909] <= 32'b11100011110000111000001110010011;
ROM[1910] <= 32'b00000000111000111000001110110011;
ROM[1911] <= 32'b00000000000000111000000011100111;
ROM[1912] <= 32'b00000000000000011010001110000011;
ROM[1913] <= 32'b00000000011100010010000000100011;
ROM[1914] <= 32'b00000000010000010000000100010011;
ROM[1915] <= 32'b00000001010001101010001110000011;
ROM[1916] <= 32'b00000000011100010010000000100011;
ROM[1917] <= 32'b00000000010000010000000100010011;
ROM[1918] <= 32'b11111111110000010000000100010011;
ROM[1919] <= 32'b00000000000000010010001110000011;
ROM[1920] <= 32'b11111111110000010000000100010011;
ROM[1921] <= 32'b00000000000000010010010000000011;
ROM[1922] <= 32'b00000000100000111000001110110011;
ROM[1923] <= 32'b00000000011100010010000000100011;
ROM[1924] <= 32'b00000000010000010000000100010011;
ROM[1925] <= 32'b11111111110000010000000100010011;
ROM[1926] <= 32'b00000000000000010010001110000011;
ROM[1927] <= 32'b00000000011100110010001000100011;
ROM[1928] <= 32'b00000000000000110010001110000011;
ROM[1929] <= 32'b00000000011100010010000000100011;
ROM[1930] <= 32'b00000000010000010000000100010011;
ROM[1931] <= 32'b11111111110000010000000100010011;
ROM[1932] <= 32'b00000000000000010010001110000011;
ROM[1933] <= 32'b00000000011100011010000000100011;
ROM[1934] <= 32'b11100100100111111111000011101111;
ROM[1935] <= 32'b00000000000000011010001110000011;
ROM[1936] <= 32'b00000000011100010010000000100011;
ROM[1937] <= 32'b00000000010000010000000100010011;
ROM[1938] <= 32'b11111111110000010000000100010011;
ROM[1939] <= 32'b00000000000000010010001110000011;
ROM[1940] <= 32'b00000000011100100010000000100011;
ROM[1941] <= 32'b00000000010000100000000100010011;
ROM[1942] <= 32'b00000001010000000000001110010011;
ROM[1943] <= 32'b01000000011100011000001110110011;
ROM[1944] <= 32'b00000000000000111010000010000011;
ROM[1945] <= 32'b00000000010000111010000110000011;
ROM[1946] <= 32'b00000000100000111010001000000011;
ROM[1947] <= 32'b00000000110000111010001010000011;
ROM[1948] <= 32'b00000001000000111010001100000011;
ROM[1949] <= 32'b00000000000000001000000011100111;
ROM[1950] <= 32'b00000000000000111000000010010011;

        end
    assign address = addr[16:2];
    assign Inst = ROM[address];
        
endmodule


						
						

// module ROM ( //Instruction Memory
//     input [15:0] address,
//     input clock,
//     input IRWrite,
//     output reg [31:0] IR
//     );
    
//     (* ram_style="block" *)
//     reg [31:0] ROM[16383:0];

//     initial
//         begin
//             $readmemb("os.mem", ROM, 0, 16383);
//             IR <= 32'd15;
//         end
    
//     always @(posedge clock)
//         begin
//             if( IRWrite )
//                 IR <= ROM[address];
//         end
        
// endmodule

						
						


						
						
