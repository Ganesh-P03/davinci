module ROM ( //Instruction Memory
    input [16:0] addr,
    input clock,
    output [31:0] Inst
    );
    wire [14:0] address;
    
    (* ram_style="block" *)
    reg [31:0] ROM[32767:0];

    initial
        begin
    ROM[0] <= 32'b00000000000000000010011100110111;
ROM[1] <= 32'b01011000000001110000011100010011;
ROM[2] <= 32'b00000000000000100010011010110111;
ROM[3] <= 32'b01011000000001101000011010010011;
ROM[4] <= 32'b00000000000001101000011000010011;
ROM[5] <= 32'b01000000000001101000000100010011;
ROM[6] <= 32'b00000000000000010000000110010011;
ROM[7] <= 32'b00000000000000010000001000010011;
ROM[8] <= 32'b00000000000000010000001010010011;
ROM[9] <= 32'b00000000000000010000001100010011;
ROM[10] <= 32'b00000000000000000000001110110111;
ROM[11] <= 32'b00000111010000111000001110010011;
ROM[12] <= 32'b00000000111000111000001110110011;
ROM[13] <= 32'b00000000011100010010000000100011;
ROM[14] <= 32'b00000000010000010000000100010011;
ROM[15] <= 32'b00000000001100010010000000100011;
ROM[16] <= 32'b00000000010000010000000100010011;
ROM[17] <= 32'b00000000010000010010000000100011;
ROM[18] <= 32'b00000000010000010000000100010011;
ROM[19] <= 32'b00000000010100010010000000100011;
ROM[20] <= 32'b00000000010000010000000100010011;
ROM[21] <= 32'b00000000011000010010000000100011;
ROM[22] <= 32'b00000000010000010000000100010011;
ROM[23] <= 32'b00000001010000000000001110010011;
ROM[24] <= 32'b00000000000000111000001110010011;
ROM[25] <= 32'b01000000011100010000001110110011;
ROM[26] <= 32'b00000000011100000000001000110011;
ROM[27] <= 32'b00000000001000000000000110110011;
ROM[28] <= 32'b01010110010100101010000011101111;
ROM[29] <= 32'b11111111110000010000000100010011;
ROM[30] <= 32'b00000000000000010010001110000011;
ROM[31] <= 32'b01010001010100101011000011101111;
ROM[32] <= 32'b00000000000000100010001110000011;
ROM[33] <= 32'b00000000011100010010000000100011;
ROM[34] <= 32'b00000000010000010000000100010011;
ROM[35] <= 32'b00000000000000000000001110110111;
ROM[36] <= 32'b00001101100000111000001110010011;
ROM[37] <= 32'b00000000111000111000001110110011;
ROM[38] <= 32'b00000000011100010010000000100011;
ROM[39] <= 32'b00000000010000010000000100010011;
ROM[40] <= 32'b00000000001100010010000000100011;
ROM[41] <= 32'b00000000010000010000000100010011;
ROM[42] <= 32'b00000000010000010010000000100011;
ROM[43] <= 32'b00000000010000010000000100010011;
ROM[44] <= 32'b00000000010100010010000000100011;
ROM[45] <= 32'b00000000010000010000000100010011;
ROM[46] <= 32'b00000000011000010010000000100011;
ROM[47] <= 32'b00000000010000010000000100010011;
ROM[48] <= 32'b00000001010000000000001110010011;
ROM[49] <= 32'b00000000010000111000001110010011;
ROM[50] <= 32'b01000000011100010000001110110011;
ROM[51] <= 32'b00000000011100000000001000110011;
ROM[52] <= 32'b00000000001000000000000110110011;
ROM[53] <= 32'b01100000000000010100000011101111;
ROM[54] <= 32'b00000001010000000000001110010011;
ROM[55] <= 32'b01000000011100011000001110110011;
ROM[56] <= 32'b00000000000000111010000010000011;
ROM[57] <= 32'b11111111110000010000000100010011;
ROM[58] <= 32'b00000000000000010010001110000011;
ROM[59] <= 32'b00000000011100100010000000100011;
ROM[60] <= 32'b00000000010000100000000100010011;
ROM[61] <= 32'b00000001010000000000001110010011;
ROM[62] <= 32'b01000000011100011000001110110011;
ROM[63] <= 32'b00000000010000111010000110000011;
ROM[64] <= 32'b00000000100000111010001000000011;
ROM[65] <= 32'b00000000110000111010001010000011;
ROM[66] <= 32'b00000001000000111010001100000011;
ROM[67] <= 32'b00000000000000001000000011100111;
ROM[68] <= 32'b00000000000000100010001110000011;
ROM[69] <= 32'b00000000011100010010000000100011;
ROM[70] <= 32'b00000000010000010000000100010011;
ROM[71] <= 32'b11111111110000010000000100010011;
ROM[72] <= 32'b00000000000000010010001110000011;
ROM[73] <= 32'b00000000000000111000001010010011;
ROM[74] <= 32'b00000000010100010010000000100011;
ROM[75] <= 32'b00000000010000010000000100010011;
ROM[76] <= 32'b00000000000000000000001110110111;
ROM[77] <= 32'b00010111110000111000001110010011;
ROM[78] <= 32'b00000000111000111000001110110011;
ROM[79] <= 32'b00000000011100010010000000100011;
ROM[80] <= 32'b00000000010000010000000100010011;
ROM[81] <= 32'b00000000001100010010000000100011;
ROM[82] <= 32'b00000000010000010000000100010011;
ROM[83] <= 32'b00000000010000010010000000100011;
ROM[84] <= 32'b00000000010000010000000100010011;
ROM[85] <= 32'b00000000010100010010000000100011;
ROM[86] <= 32'b00000000010000010000000100010011;
ROM[87] <= 32'b00000000011000010010000000100011;
ROM[88] <= 32'b00000000010000010000000100010011;
ROM[89] <= 32'b00000001010000000000001110010011;
ROM[90] <= 32'b00000000010000111000001110010011;
ROM[91] <= 32'b01000000011100010000001110110011;
ROM[92] <= 32'b00000000011100000000001000110011;
ROM[93] <= 32'b00000000001000000000000110110011;
ROM[94] <= 32'b00011110010100010011000011101111;
ROM[95] <= 32'b11111111110000010000000100010011;
ROM[96] <= 32'b00000000000000010010001110000011;
ROM[97] <= 32'b00000000011101100010000000100011;
ROM[98] <= 32'b00000000000000000000001110010011;
ROM[99] <= 32'b00000000011100010010000000100011;
ROM[100] <= 32'b00000000010000010000000100010011;
ROM[101] <= 32'b00000001010000000000001110010011;
ROM[102] <= 32'b01000000011100011000001110110011;
ROM[103] <= 32'b00000000000000111010000010000011;
ROM[104] <= 32'b11111111110000010000000100010011;
ROM[105] <= 32'b00000000000000010010001110000011;
ROM[106] <= 32'b00000000011100100010000000100011;
ROM[107] <= 32'b00000000010000100000000100010011;
ROM[108] <= 32'b00000001010000000000001110010011;
ROM[109] <= 32'b01000000011100011000001110110011;
ROM[110] <= 32'b00000000010000111010000110000011;
ROM[111] <= 32'b00000000100000111010001000000011;
ROM[112] <= 32'b00000000110000111010001010000011;
ROM[113] <= 32'b00000001000000111010001100000011;
ROM[114] <= 32'b00000000000000001000000011100111;
ROM[115] <= 32'b00000000000000010010000000100011;
ROM[116] <= 32'b00000000010000010000000100010011;
ROM[117] <= 32'b00000000000000010010000000100011;
ROM[118] <= 32'b00000000010000010000000100010011;
ROM[119] <= 32'b00000000000000010010000000100011;
ROM[120] <= 32'b00000000010000010000000100010011;
ROM[121] <= 32'b00000000000000010010000000100011;
ROM[122] <= 32'b00000000010000010000000100010011;
ROM[123] <= 32'b00000000000000010010000000100011;
ROM[124] <= 32'b00000000010000010000000100010011;
ROM[125] <= 32'b00000011000000000000001110010011;
ROM[126] <= 32'b00000000011100010010000000100011;
ROM[127] <= 32'b00000000010000010000000100010011;
ROM[128] <= 32'b00000000000000000000001110110111;
ROM[129] <= 32'b00100100110000111000001110010011;
ROM[130] <= 32'b00000000111000111000001110110011;
ROM[131] <= 32'b00000000011100010010000000100011;
ROM[132] <= 32'b00000000010000010000000100010011;
ROM[133] <= 32'b00000000001100010010000000100011;
ROM[134] <= 32'b00000000010000010000000100010011;
ROM[135] <= 32'b00000000010000010010000000100011;
ROM[136] <= 32'b00000000010000010000000100010011;
ROM[137] <= 32'b00000000010100010010000000100011;
ROM[138] <= 32'b00000000010000010000000100010011;
ROM[139] <= 32'b00000000011000010010000000100011;
ROM[140] <= 32'b00000000010000010000000100010011;
ROM[141] <= 32'b00000001010000000000001110010011;
ROM[142] <= 32'b00000000010000111000001110010011;
ROM[143] <= 32'b01000000011100010000001110110011;
ROM[144] <= 32'b00000000011100000000001000110011;
ROM[145] <= 32'b00000000001000000000000110110011;
ROM[146] <= 32'b01001111010000101001000011101111;
ROM[147] <= 32'b00000100010100000000001110010011;
ROM[148] <= 32'b00000000011100010010000000100011;
ROM[149] <= 32'b00000000010000010000000100010011;
ROM[150] <= 32'b00000000000000000000001110110111;
ROM[151] <= 32'b00101010010000111000001110010011;
ROM[152] <= 32'b00000000111000111000001110110011;
ROM[153] <= 32'b00000000011100010010000000100011;
ROM[154] <= 32'b00000000010000010000000100010011;
ROM[155] <= 32'b00000000001100010010000000100011;
ROM[156] <= 32'b00000000010000010000000100010011;
ROM[157] <= 32'b00000000010000010010000000100011;
ROM[158] <= 32'b00000000010000010000000100010011;
ROM[159] <= 32'b00000000010100010010000000100011;
ROM[160] <= 32'b00000000010000010000000100010011;
ROM[161] <= 32'b00000000011000010010000000100011;
ROM[162] <= 32'b00000000010000010000000100010011;
ROM[163] <= 32'b00000001010000000000001110010011;
ROM[164] <= 32'b00000000100000111000001110010011;
ROM[165] <= 32'b01000000011100010000001110110011;
ROM[166] <= 32'b00000000011100000000001000110011;
ROM[167] <= 32'b00000000001000000000000110110011;
ROM[168] <= 32'b00010000110100101001000011101111;
ROM[169] <= 32'b00000110111000000000001110010011;
ROM[170] <= 32'b00000000011100010010000000100011;
ROM[171] <= 32'b00000000010000010000000100010011;
ROM[172] <= 32'b00000000000000000000001110110111;
ROM[173] <= 32'b00101111110000111000001110010011;
ROM[174] <= 32'b00000000111000111000001110110011;
ROM[175] <= 32'b00000000011100010010000000100011;
ROM[176] <= 32'b00000000010000010000000100010011;
ROM[177] <= 32'b00000000001100010010000000100011;
ROM[178] <= 32'b00000000010000010000000100010011;
ROM[179] <= 32'b00000000010000010010000000100011;
ROM[180] <= 32'b00000000010000010000000100010011;
ROM[181] <= 32'b00000000010100010010000000100011;
ROM[182] <= 32'b00000000010000010000000100010011;
ROM[183] <= 32'b00000000011000010010000000100011;
ROM[184] <= 32'b00000000010000010000000100010011;
ROM[185] <= 32'b00000001010000000000001110010011;
ROM[186] <= 32'b00000000100000111000001110010011;
ROM[187] <= 32'b01000000011100010000001110110011;
ROM[188] <= 32'b00000000011100000000001000110011;
ROM[189] <= 32'b00000000001000000000000110110011;
ROM[190] <= 32'b00001011010100101001000011101111;
ROM[191] <= 32'b00000111010000000000001110010011;
ROM[192] <= 32'b00000000011100010010000000100011;
ROM[193] <= 32'b00000000010000010000000100010011;
ROM[194] <= 32'b00000000000000000000001110110111;
ROM[195] <= 32'b00110101010000111000001110010011;
ROM[196] <= 32'b00000000111000111000001110110011;
ROM[197] <= 32'b00000000011100010010000000100011;
ROM[198] <= 32'b00000000010000010000000100010011;
ROM[199] <= 32'b00000000001100010010000000100011;
ROM[200] <= 32'b00000000010000010000000100010011;
ROM[201] <= 32'b00000000010000010010000000100011;
ROM[202] <= 32'b00000000010000010000000100010011;
ROM[203] <= 32'b00000000010100010010000000100011;
ROM[204] <= 32'b00000000010000010000000100010011;
ROM[205] <= 32'b00000000011000010010000000100011;
ROM[206] <= 32'b00000000010000010000000100010011;
ROM[207] <= 32'b00000001010000000000001110010011;
ROM[208] <= 32'b00000000100000111000001110010011;
ROM[209] <= 32'b01000000011100010000001110110011;
ROM[210] <= 32'b00000000011100000000001000110011;
ROM[211] <= 32'b00000000001000000000000110110011;
ROM[212] <= 32'b00000101110100101001000011101111;
ROM[213] <= 32'b00000110010100000000001110010011;
ROM[214] <= 32'b00000000011100010010000000100011;
ROM[215] <= 32'b00000000010000010000000100010011;
ROM[216] <= 32'b00000000000000000000001110110111;
ROM[217] <= 32'b00111010110000111000001110010011;
ROM[218] <= 32'b00000000111000111000001110110011;
ROM[219] <= 32'b00000000011100010010000000100011;
ROM[220] <= 32'b00000000010000010000000100010011;
ROM[221] <= 32'b00000000001100010010000000100011;
ROM[222] <= 32'b00000000010000010000000100010011;
ROM[223] <= 32'b00000000010000010010000000100011;
ROM[224] <= 32'b00000000010000010000000100010011;
ROM[225] <= 32'b00000000010100010010000000100011;
ROM[226] <= 32'b00000000010000010000000100010011;
ROM[227] <= 32'b00000000011000010010000000100011;
ROM[228] <= 32'b00000000010000010000000100010011;
ROM[229] <= 32'b00000001010000000000001110010011;
ROM[230] <= 32'b00000000100000111000001110010011;
ROM[231] <= 32'b01000000011100010000001110110011;
ROM[232] <= 32'b00000000011100000000001000110011;
ROM[233] <= 32'b00000000001000000000000110110011;
ROM[234] <= 32'b00000000010100101001000011101111;
ROM[235] <= 32'b00000111001000000000001110010011;
ROM[236] <= 32'b00000000011100010010000000100011;
ROM[237] <= 32'b00000000010000010000000100010011;
ROM[238] <= 32'b00000000000000000000001110110111;
ROM[239] <= 32'b01000000010000111000001110010011;
ROM[240] <= 32'b00000000111000111000001110110011;
ROM[241] <= 32'b00000000011100010010000000100011;
ROM[242] <= 32'b00000000010000010000000100010011;
ROM[243] <= 32'b00000000001100010010000000100011;
ROM[244] <= 32'b00000000010000010000000100010011;
ROM[245] <= 32'b00000000010000010010000000100011;
ROM[246] <= 32'b00000000010000010000000100010011;
ROM[247] <= 32'b00000000010100010010000000100011;
ROM[248] <= 32'b00000000010000010000000100010011;
ROM[249] <= 32'b00000000011000010010000000100011;
ROM[250] <= 32'b00000000010000010000000100010011;
ROM[251] <= 32'b00000001010000000000001110010011;
ROM[252] <= 32'b00000000100000111000001110010011;
ROM[253] <= 32'b01000000011100010000001110110011;
ROM[254] <= 32'b00000000011100000000001000110011;
ROM[255] <= 32'b00000000001000000000000110110011;
ROM[256] <= 32'b01111010110000101001000011101111;
ROM[257] <= 32'b00000010000000000000001110010011;
ROM[258] <= 32'b00000000011100010010000000100011;
ROM[259] <= 32'b00000000010000010000000100010011;
ROM[260] <= 32'b00000000000000000000001110110111;
ROM[261] <= 32'b01000101110000111000001110010011;
ROM[262] <= 32'b00000000111000111000001110110011;
ROM[263] <= 32'b00000000011100010010000000100011;
ROM[264] <= 32'b00000000010000010000000100010011;
ROM[265] <= 32'b00000000001100010010000000100011;
ROM[266] <= 32'b00000000010000010000000100010011;
ROM[267] <= 32'b00000000010000010010000000100011;
ROM[268] <= 32'b00000000010000010000000100010011;
ROM[269] <= 32'b00000000010100010010000000100011;
ROM[270] <= 32'b00000000010000010000000100010011;
ROM[271] <= 32'b00000000011000010010000000100011;
ROM[272] <= 32'b00000000010000010000000100010011;
ROM[273] <= 32'b00000001010000000000001110010011;
ROM[274] <= 32'b00000000100000111000001110010011;
ROM[275] <= 32'b01000000011100010000001110110011;
ROM[276] <= 32'b00000000011100000000001000110011;
ROM[277] <= 32'b00000000001000000000000110110011;
ROM[278] <= 32'b01110101010000101001000011101111;
ROM[279] <= 32'b00000111010000000000001110010011;
ROM[280] <= 32'b00000000011100010010000000100011;
ROM[281] <= 32'b00000000010000010000000100010011;
ROM[282] <= 32'b00000000000000000000001110110111;
ROM[283] <= 32'b01001011010000111000001110010011;
ROM[284] <= 32'b00000000111000111000001110110011;
ROM[285] <= 32'b00000000011100010010000000100011;
ROM[286] <= 32'b00000000010000010000000100010011;
ROM[287] <= 32'b00000000001100010010000000100011;
ROM[288] <= 32'b00000000010000010000000100010011;
ROM[289] <= 32'b00000000010000010010000000100011;
ROM[290] <= 32'b00000000010000010000000100010011;
ROM[291] <= 32'b00000000010100010010000000100011;
ROM[292] <= 32'b00000000010000010000000100010011;
ROM[293] <= 32'b00000000011000010010000000100011;
ROM[294] <= 32'b00000000010000010000000100010011;
ROM[295] <= 32'b00000001010000000000001110010011;
ROM[296] <= 32'b00000000100000111000001110010011;
ROM[297] <= 32'b01000000011100010000001110110011;
ROM[298] <= 32'b00000000011100000000001000110011;
ROM[299] <= 32'b00000000001000000000000110110011;
ROM[300] <= 32'b01101111110000101001000011101111;
ROM[301] <= 32'b00000110100000000000001110010011;
ROM[302] <= 32'b00000000011100010010000000100011;
ROM[303] <= 32'b00000000010000010000000100010011;
ROM[304] <= 32'b00000000000000000000001110110111;
ROM[305] <= 32'b01010000110000111000001110010011;
ROM[306] <= 32'b00000000111000111000001110110011;
ROM[307] <= 32'b00000000011100010010000000100011;
ROM[308] <= 32'b00000000010000010000000100010011;
ROM[309] <= 32'b00000000001100010010000000100011;
ROM[310] <= 32'b00000000010000010000000100010011;
ROM[311] <= 32'b00000000010000010010000000100011;
ROM[312] <= 32'b00000000010000010000000100010011;
ROM[313] <= 32'b00000000010100010010000000100011;
ROM[314] <= 32'b00000000010000010000000100010011;
ROM[315] <= 32'b00000000011000010010000000100011;
ROM[316] <= 32'b00000000010000010000000100010011;
ROM[317] <= 32'b00000001010000000000001110010011;
ROM[318] <= 32'b00000000100000111000001110010011;
ROM[319] <= 32'b01000000011100010000001110110011;
ROM[320] <= 32'b00000000011100000000001000110011;
ROM[321] <= 32'b00000000001000000000000110110011;
ROM[322] <= 32'b01101010010000101001000011101111;
ROM[323] <= 32'b00000110010100000000001110010011;
ROM[324] <= 32'b00000000011100010010000000100011;
ROM[325] <= 32'b00000000010000010000000100010011;
ROM[326] <= 32'b00000000000000000000001110110111;
ROM[327] <= 32'b01010110010000111000001110010011;
ROM[328] <= 32'b00000000111000111000001110110011;
ROM[329] <= 32'b00000000011100010010000000100011;
ROM[330] <= 32'b00000000010000010000000100010011;
ROM[331] <= 32'b00000000001100010010000000100011;
ROM[332] <= 32'b00000000010000010000000100010011;
ROM[333] <= 32'b00000000010000010010000000100011;
ROM[334] <= 32'b00000000010000010000000100010011;
ROM[335] <= 32'b00000000010100010010000000100011;
ROM[336] <= 32'b00000000010000010000000100010011;
ROM[337] <= 32'b00000000011000010010000000100011;
ROM[338] <= 32'b00000000010000010000000100010011;
ROM[339] <= 32'b00000001010000000000001110010011;
ROM[340] <= 32'b00000000100000111000001110010011;
ROM[341] <= 32'b01000000011100010000001110110011;
ROM[342] <= 32'b00000000011100000000001000110011;
ROM[343] <= 32'b00000000001000000000000110110011;
ROM[344] <= 32'b01100100110000101001000011101111;
ROM[345] <= 32'b00000010000000000000001110010011;
ROM[346] <= 32'b00000000011100010010000000100011;
ROM[347] <= 32'b00000000010000010000000100010011;
ROM[348] <= 32'b00000000000000000000001110110111;
ROM[349] <= 32'b01011011110000111000001110010011;
ROM[350] <= 32'b00000000111000111000001110110011;
ROM[351] <= 32'b00000000011100010010000000100011;
ROM[352] <= 32'b00000000010000010000000100010011;
ROM[353] <= 32'b00000000001100010010000000100011;
ROM[354] <= 32'b00000000010000010000000100010011;
ROM[355] <= 32'b00000000010000010010000000100011;
ROM[356] <= 32'b00000000010000010000000100010011;
ROM[357] <= 32'b00000000010100010010000000100011;
ROM[358] <= 32'b00000000010000010000000100010011;
ROM[359] <= 32'b00000000011000010010000000100011;
ROM[360] <= 32'b00000000010000010000000100010011;
ROM[361] <= 32'b00000001010000000000001110010011;
ROM[362] <= 32'b00000000100000111000001110010011;
ROM[363] <= 32'b01000000011100010000001110110011;
ROM[364] <= 32'b00000000011100000000001000110011;
ROM[365] <= 32'b00000000001000000000000110110011;
ROM[366] <= 32'b01011111010000101001000011101111;
ROM[367] <= 32'b00000110111000000000001110010011;
ROM[368] <= 32'b00000000011100010010000000100011;
ROM[369] <= 32'b00000000010000010000000100010011;
ROM[370] <= 32'b00000000000000000000001110110111;
ROM[371] <= 32'b01100001010000111000001110010011;
ROM[372] <= 32'b00000000111000111000001110110011;
ROM[373] <= 32'b00000000011100010010000000100011;
ROM[374] <= 32'b00000000010000010000000100010011;
ROM[375] <= 32'b00000000001100010010000000100011;
ROM[376] <= 32'b00000000010000010000000100010011;
ROM[377] <= 32'b00000000010000010010000000100011;
ROM[378] <= 32'b00000000010000010000000100010011;
ROM[379] <= 32'b00000000010100010010000000100011;
ROM[380] <= 32'b00000000010000010000000100010011;
ROM[381] <= 32'b00000000011000010010000000100011;
ROM[382] <= 32'b00000000010000010000000100010011;
ROM[383] <= 32'b00000001010000000000001110010011;
ROM[384] <= 32'b00000000100000111000001110010011;
ROM[385] <= 32'b01000000011100010000001110110011;
ROM[386] <= 32'b00000000011100000000001000110011;
ROM[387] <= 32'b00000000001000000000000110110011;
ROM[388] <= 32'b01011001110000101001000011101111;
ROM[389] <= 32'b00000111010100000000001110010011;
ROM[390] <= 32'b00000000011100010010000000100011;
ROM[391] <= 32'b00000000010000010000000100010011;
ROM[392] <= 32'b00000000000000000000001110110111;
ROM[393] <= 32'b01100110110000111000001110010011;
ROM[394] <= 32'b00000000111000111000001110110011;
ROM[395] <= 32'b00000000011100010010000000100011;
ROM[396] <= 32'b00000000010000010000000100010011;
ROM[397] <= 32'b00000000001100010010000000100011;
ROM[398] <= 32'b00000000010000010000000100010011;
ROM[399] <= 32'b00000000010000010010000000100011;
ROM[400] <= 32'b00000000010000010000000100010011;
ROM[401] <= 32'b00000000010100010010000000100011;
ROM[402] <= 32'b00000000010000010000000100010011;
ROM[403] <= 32'b00000000011000010010000000100011;
ROM[404] <= 32'b00000000010000010000000100010011;
ROM[405] <= 32'b00000001010000000000001110010011;
ROM[406] <= 32'b00000000100000111000001110010011;
ROM[407] <= 32'b01000000011100010000001110110011;
ROM[408] <= 32'b00000000011100000000001000110011;
ROM[409] <= 32'b00000000001000000000000110110011;
ROM[410] <= 32'b01010100010000101001000011101111;
ROM[411] <= 32'b00000110110100000000001110010011;
ROM[412] <= 32'b00000000011100010010000000100011;
ROM[413] <= 32'b00000000010000010000000100010011;
ROM[414] <= 32'b00000000000000000000001110110111;
ROM[415] <= 32'b01101100010000111000001110010011;
ROM[416] <= 32'b00000000111000111000001110110011;
ROM[417] <= 32'b00000000011100010010000000100011;
ROM[418] <= 32'b00000000010000010000000100010011;
ROM[419] <= 32'b00000000001100010010000000100011;
ROM[420] <= 32'b00000000010000010000000100010011;
ROM[421] <= 32'b00000000010000010010000000100011;
ROM[422] <= 32'b00000000010000010000000100010011;
ROM[423] <= 32'b00000000010100010010000000100011;
ROM[424] <= 32'b00000000010000010000000100010011;
ROM[425] <= 32'b00000000011000010010000000100011;
ROM[426] <= 32'b00000000010000010000000100010011;
ROM[427] <= 32'b00000001010000000000001110010011;
ROM[428] <= 32'b00000000100000111000001110010011;
ROM[429] <= 32'b01000000011100010000001110110011;
ROM[430] <= 32'b00000000011100000000001000110011;
ROM[431] <= 32'b00000000001000000000000110110011;
ROM[432] <= 32'b01001110110000101001000011101111;
ROM[433] <= 32'b00000110001000000000001110010011;
ROM[434] <= 32'b00000000011100010010000000100011;
ROM[435] <= 32'b00000000010000010000000100010011;
ROM[436] <= 32'b00000000000000000000001110110111;
ROM[437] <= 32'b01110001110000111000001110010011;
ROM[438] <= 32'b00000000111000111000001110110011;
ROM[439] <= 32'b00000000011100010010000000100011;
ROM[440] <= 32'b00000000010000010000000100010011;
ROM[441] <= 32'b00000000001100010010000000100011;
ROM[442] <= 32'b00000000010000010000000100010011;
ROM[443] <= 32'b00000000010000010010000000100011;
ROM[444] <= 32'b00000000010000010000000100010011;
ROM[445] <= 32'b00000000010100010010000000100011;
ROM[446] <= 32'b00000000010000010000000100010011;
ROM[447] <= 32'b00000000011000010010000000100011;
ROM[448] <= 32'b00000000010000010000000100010011;
ROM[449] <= 32'b00000001010000000000001110010011;
ROM[450] <= 32'b00000000100000111000001110010011;
ROM[451] <= 32'b01000000011100010000001110110011;
ROM[452] <= 32'b00000000011100000000001000110011;
ROM[453] <= 32'b00000000001000000000000110110011;
ROM[454] <= 32'b01001001010000101001000011101111;
ROM[455] <= 32'b00000110010100000000001110010011;
ROM[456] <= 32'b00000000011100010010000000100011;
ROM[457] <= 32'b00000000010000010000000100010011;
ROM[458] <= 32'b00000000000000000000001110110111;
ROM[459] <= 32'b01110111010000111000001110010011;
ROM[460] <= 32'b00000000111000111000001110110011;
ROM[461] <= 32'b00000000011100010010000000100011;
ROM[462] <= 32'b00000000010000010000000100010011;
ROM[463] <= 32'b00000000001100010010000000100011;
ROM[464] <= 32'b00000000010000010000000100010011;
ROM[465] <= 32'b00000000010000010010000000100011;
ROM[466] <= 32'b00000000010000010000000100010011;
ROM[467] <= 32'b00000000010100010010000000100011;
ROM[468] <= 32'b00000000010000010000000100010011;
ROM[469] <= 32'b00000000011000010010000000100011;
ROM[470] <= 32'b00000000010000010000000100010011;
ROM[471] <= 32'b00000001010000000000001110010011;
ROM[472] <= 32'b00000000100000111000001110010011;
ROM[473] <= 32'b01000000011100010000001110110011;
ROM[474] <= 32'b00000000011100000000001000110011;
ROM[475] <= 32'b00000000001000000000000110110011;
ROM[476] <= 32'b01000011110000101001000011101111;
ROM[477] <= 32'b00000111001000000000001110010011;
ROM[478] <= 32'b00000000011100010010000000100011;
ROM[479] <= 32'b00000000010000010000000100010011;
ROM[480] <= 32'b00000000000000000000001110110111;
ROM[481] <= 32'b01111100110000111000001110010011;
ROM[482] <= 32'b00000000111000111000001110110011;
ROM[483] <= 32'b00000000011100010010000000100011;
ROM[484] <= 32'b00000000010000010000000100010011;
ROM[485] <= 32'b00000000001100010010000000100011;
ROM[486] <= 32'b00000000010000010000000100010011;
ROM[487] <= 32'b00000000010000010010000000100011;
ROM[488] <= 32'b00000000010000010000000100010011;
ROM[489] <= 32'b00000000010100010010000000100011;
ROM[490] <= 32'b00000000010000010000000100010011;
ROM[491] <= 32'b00000000011000010010000000100011;
ROM[492] <= 32'b00000000010000010000000100010011;
ROM[493] <= 32'b00000001010000000000001110010011;
ROM[494] <= 32'b00000000100000111000001110010011;
ROM[495] <= 32'b01000000011100010000001110110011;
ROM[496] <= 32'b00000000011100000000001000110011;
ROM[497] <= 32'b00000000001000000000000110110011;
ROM[498] <= 32'b00111110010000101001000011101111;
ROM[499] <= 32'b00000010000000000000001110010011;
ROM[500] <= 32'b00000000011100010010000000100011;
ROM[501] <= 32'b00000000010000010000000100010011;
ROM[502] <= 32'b00000000000000000001001110110111;
ROM[503] <= 32'b10000010010000111000001110010011;
ROM[504] <= 32'b00000000111000111000001110110011;
ROM[505] <= 32'b00000000011100010010000000100011;
ROM[506] <= 32'b00000000010000010000000100010011;
ROM[507] <= 32'b00000000001100010010000000100011;
ROM[508] <= 32'b00000000010000010000000100010011;
ROM[509] <= 32'b00000000010000010010000000100011;
ROM[510] <= 32'b00000000010000010000000100010011;
ROM[511] <= 32'b00000000010100010010000000100011;
ROM[512] <= 32'b00000000010000010000000100010011;
ROM[513] <= 32'b00000000011000010010000000100011;
ROM[514] <= 32'b00000000010000010000000100010011;
ROM[515] <= 32'b00000001010000000000001110010011;
ROM[516] <= 32'b00000000100000111000001110010011;
ROM[517] <= 32'b01000000011100010000001110110011;
ROM[518] <= 32'b00000000011100000000001000110011;
ROM[519] <= 32'b00000000001000000000000110110011;
ROM[520] <= 32'b00111000110000101001000011101111;
ROM[521] <= 32'b00000110111100000000001110010011;
ROM[522] <= 32'b00000000011100010010000000100011;
ROM[523] <= 32'b00000000010000010000000100010011;
ROM[524] <= 32'b00000000000000000001001110110111;
ROM[525] <= 32'b10000111110000111000001110010011;
ROM[526] <= 32'b00000000111000111000001110110011;
ROM[527] <= 32'b00000000011100010010000000100011;
ROM[528] <= 32'b00000000010000010000000100010011;
ROM[529] <= 32'b00000000001100010010000000100011;
ROM[530] <= 32'b00000000010000010000000100010011;
ROM[531] <= 32'b00000000010000010010000000100011;
ROM[532] <= 32'b00000000010000010000000100010011;
ROM[533] <= 32'b00000000010100010010000000100011;
ROM[534] <= 32'b00000000010000010000000100010011;
ROM[535] <= 32'b00000000011000010010000000100011;
ROM[536] <= 32'b00000000010000010000000100010011;
ROM[537] <= 32'b00000001010000000000001110010011;
ROM[538] <= 32'b00000000100000111000001110010011;
ROM[539] <= 32'b01000000011100010000001110110011;
ROM[540] <= 32'b00000000011100000000001000110011;
ROM[541] <= 32'b00000000001000000000000110110011;
ROM[542] <= 32'b00110011010000101001000011101111;
ROM[543] <= 32'b00000110011000000000001110010011;
ROM[544] <= 32'b00000000011100010010000000100011;
ROM[545] <= 32'b00000000010000010000000100010011;
ROM[546] <= 32'b00000000000000000001001110110111;
ROM[547] <= 32'b10001101010000111000001110010011;
ROM[548] <= 32'b00000000111000111000001110110011;
ROM[549] <= 32'b00000000011100010010000000100011;
ROM[550] <= 32'b00000000010000010000000100010011;
ROM[551] <= 32'b00000000001100010010000000100011;
ROM[552] <= 32'b00000000010000010000000100010011;
ROM[553] <= 32'b00000000010000010010000000100011;
ROM[554] <= 32'b00000000010000010000000100010011;
ROM[555] <= 32'b00000000010100010010000000100011;
ROM[556] <= 32'b00000000010000010000000100010011;
ROM[557] <= 32'b00000000011000010010000000100011;
ROM[558] <= 32'b00000000010000010000000100010011;
ROM[559] <= 32'b00000001010000000000001110010011;
ROM[560] <= 32'b00000000100000111000001110010011;
ROM[561] <= 32'b01000000011100010000001110110011;
ROM[562] <= 32'b00000000011100000000001000110011;
ROM[563] <= 32'b00000000001000000000000110110011;
ROM[564] <= 32'b00101101110000101001000011101111;
ROM[565] <= 32'b00000010000000000000001110010011;
ROM[566] <= 32'b00000000011100010010000000100011;
ROM[567] <= 32'b00000000010000010000000100010011;
ROM[568] <= 32'b00000000000000000001001110110111;
ROM[569] <= 32'b10010010110000111000001110010011;
ROM[570] <= 32'b00000000111000111000001110110011;
ROM[571] <= 32'b00000000011100010010000000100011;
ROM[572] <= 32'b00000000010000010000000100010011;
ROM[573] <= 32'b00000000001100010010000000100011;
ROM[574] <= 32'b00000000010000010000000100010011;
ROM[575] <= 32'b00000000010000010010000000100011;
ROM[576] <= 32'b00000000010000010000000100010011;
ROM[577] <= 32'b00000000010100010010000000100011;
ROM[578] <= 32'b00000000010000010000000100010011;
ROM[579] <= 32'b00000000011000010010000000100011;
ROM[580] <= 32'b00000000010000010000000100010011;
ROM[581] <= 32'b00000001010000000000001110010011;
ROM[582] <= 32'b00000000100000111000001110010011;
ROM[583] <= 32'b01000000011100010000001110110011;
ROM[584] <= 32'b00000000011100000000001000110011;
ROM[585] <= 32'b00000000001000000000000110110011;
ROM[586] <= 32'b00101000010000101001000011101111;
ROM[587] <= 32'b00000100011000000000001110010011;
ROM[588] <= 32'b00000000011100010010000000100011;
ROM[589] <= 32'b00000000010000010000000100010011;
ROM[590] <= 32'b00000000000000000001001110110111;
ROM[591] <= 32'b10011000010000111000001110010011;
ROM[592] <= 32'b00000000111000111000001110110011;
ROM[593] <= 32'b00000000011100010010000000100011;
ROM[594] <= 32'b00000000010000010000000100010011;
ROM[595] <= 32'b00000000001100010010000000100011;
ROM[596] <= 32'b00000000010000010000000100010011;
ROM[597] <= 32'b00000000010000010010000000100011;
ROM[598] <= 32'b00000000010000010000000100010011;
ROM[599] <= 32'b00000000010100010010000000100011;
ROM[600] <= 32'b00000000010000010000000100010011;
ROM[601] <= 32'b00000000011000010010000000100011;
ROM[602] <= 32'b00000000010000010000000100010011;
ROM[603] <= 32'b00000001010000000000001110010011;
ROM[604] <= 32'b00000000100000111000001110010011;
ROM[605] <= 32'b01000000011100010000001110110011;
ROM[606] <= 32'b00000000011100000000001000110011;
ROM[607] <= 32'b00000000001000000000000110110011;
ROM[608] <= 32'b00100010110000101001000011101111;
ROM[609] <= 32'b00000110100100000000001110010011;
ROM[610] <= 32'b00000000011100010010000000100011;
ROM[611] <= 32'b00000000010000010000000100010011;
ROM[612] <= 32'b00000000000000000001001110110111;
ROM[613] <= 32'b10011101110000111000001110010011;
ROM[614] <= 32'b00000000111000111000001110110011;
ROM[615] <= 32'b00000000011100010010000000100011;
ROM[616] <= 32'b00000000010000010000000100010011;
ROM[617] <= 32'b00000000001100010010000000100011;
ROM[618] <= 32'b00000000010000010000000100010011;
ROM[619] <= 32'b00000000010000010010000000100011;
ROM[620] <= 32'b00000000010000010000000100010011;
ROM[621] <= 32'b00000000010100010010000000100011;
ROM[622] <= 32'b00000000010000010000000100010011;
ROM[623] <= 32'b00000000011000010010000000100011;
ROM[624] <= 32'b00000000010000010000000100010011;
ROM[625] <= 32'b00000001010000000000001110010011;
ROM[626] <= 32'b00000000100000111000001110010011;
ROM[627] <= 32'b01000000011100010000001110110011;
ROM[628] <= 32'b00000000011100000000001000110011;
ROM[629] <= 32'b00000000001000000000000110110011;
ROM[630] <= 32'b00011101010000101001000011101111;
ROM[631] <= 32'b00000110001000000000001110010011;
ROM[632] <= 32'b00000000011100010010000000100011;
ROM[633] <= 32'b00000000010000010000000100010011;
ROM[634] <= 32'b00000000000000000001001110110111;
ROM[635] <= 32'b10100011010000111000001110010011;
ROM[636] <= 32'b00000000111000111000001110110011;
ROM[637] <= 32'b00000000011100010010000000100011;
ROM[638] <= 32'b00000000010000010000000100010011;
ROM[639] <= 32'b00000000001100010010000000100011;
ROM[640] <= 32'b00000000010000010000000100010011;
ROM[641] <= 32'b00000000010000010010000000100011;
ROM[642] <= 32'b00000000010000010000000100010011;
ROM[643] <= 32'b00000000010100010010000000100011;
ROM[644] <= 32'b00000000010000010000000100010011;
ROM[645] <= 32'b00000000011000010010000000100011;
ROM[646] <= 32'b00000000010000010000000100010011;
ROM[647] <= 32'b00000001010000000000001110010011;
ROM[648] <= 32'b00000000100000111000001110010011;
ROM[649] <= 32'b01000000011100010000001110110011;
ROM[650] <= 32'b00000000011100000000001000110011;
ROM[651] <= 32'b00000000001000000000000110110011;
ROM[652] <= 32'b00010111110000101001000011101111;
ROM[653] <= 32'b00000110111100000000001110010011;
ROM[654] <= 32'b00000000011100010010000000100011;
ROM[655] <= 32'b00000000010000010000000100010011;
ROM[656] <= 32'b00000000000000000001001110110111;
ROM[657] <= 32'b10101000110000111000001110010011;
ROM[658] <= 32'b00000000111000111000001110110011;
ROM[659] <= 32'b00000000011100010010000000100011;
ROM[660] <= 32'b00000000010000010000000100010011;
ROM[661] <= 32'b00000000001100010010000000100011;
ROM[662] <= 32'b00000000010000010000000100010011;
ROM[663] <= 32'b00000000010000010010000000100011;
ROM[664] <= 32'b00000000010000010000000100010011;
ROM[665] <= 32'b00000000010100010010000000100011;
ROM[666] <= 32'b00000000010000010000000100010011;
ROM[667] <= 32'b00000000011000010010000000100011;
ROM[668] <= 32'b00000000010000010000000100010011;
ROM[669] <= 32'b00000001010000000000001110010011;
ROM[670] <= 32'b00000000100000111000001110010011;
ROM[671] <= 32'b01000000011100010000001110110011;
ROM[672] <= 32'b00000000011100000000001000110011;
ROM[673] <= 32'b00000000001000000000000110110011;
ROM[674] <= 32'b00010010010000101001000011101111;
ROM[675] <= 32'b00000110111000000000001110010011;
ROM[676] <= 32'b00000000011100010010000000100011;
ROM[677] <= 32'b00000000010000010000000100010011;
ROM[678] <= 32'b00000000000000000001001110110111;
ROM[679] <= 32'b10101110010000111000001110010011;
ROM[680] <= 32'b00000000111000111000001110110011;
ROM[681] <= 32'b00000000011100010010000000100011;
ROM[682] <= 32'b00000000010000010000000100010011;
ROM[683] <= 32'b00000000001100010010000000100011;
ROM[684] <= 32'b00000000010000010000000100010011;
ROM[685] <= 32'b00000000010000010010000000100011;
ROM[686] <= 32'b00000000010000010000000100010011;
ROM[687] <= 32'b00000000010100010010000000100011;
ROM[688] <= 32'b00000000010000010000000100010011;
ROM[689] <= 32'b00000000011000010010000000100011;
ROM[690] <= 32'b00000000010000010000000100010011;
ROM[691] <= 32'b00000001010000000000001110010011;
ROM[692] <= 32'b00000000100000111000001110010011;
ROM[693] <= 32'b01000000011100010000001110110011;
ROM[694] <= 32'b00000000011100000000001000110011;
ROM[695] <= 32'b00000000001000000000000110110011;
ROM[696] <= 32'b00001100110000101001000011101111;
ROM[697] <= 32'b00000110000100000000001110010011;
ROM[698] <= 32'b00000000011100010010000000100011;
ROM[699] <= 32'b00000000010000010000000100010011;
ROM[700] <= 32'b00000000000000000001001110110111;
ROM[701] <= 32'b10110011110000111000001110010011;
ROM[702] <= 32'b00000000111000111000001110110011;
ROM[703] <= 32'b00000000011100010010000000100011;
ROM[704] <= 32'b00000000010000010000000100010011;
ROM[705] <= 32'b00000000001100010010000000100011;
ROM[706] <= 32'b00000000010000010000000100010011;
ROM[707] <= 32'b00000000010000010010000000100011;
ROM[708] <= 32'b00000000010000010000000100010011;
ROM[709] <= 32'b00000000010100010010000000100011;
ROM[710] <= 32'b00000000010000010000000100010011;
ROM[711] <= 32'b00000000011000010010000000100011;
ROM[712] <= 32'b00000000010000010000000100010011;
ROM[713] <= 32'b00000001010000000000001110010011;
ROM[714] <= 32'b00000000100000111000001110010011;
ROM[715] <= 32'b01000000011100010000001110110011;
ROM[716] <= 32'b00000000011100000000001000110011;
ROM[717] <= 32'b00000000001000000000000110110011;
ROM[718] <= 32'b00000111010000101001000011101111;
ROM[719] <= 32'b00000110001100000000001110010011;
ROM[720] <= 32'b00000000011100010010000000100011;
ROM[721] <= 32'b00000000010000010000000100010011;
ROM[722] <= 32'b00000000000000000001001110110111;
ROM[723] <= 32'b10111001010000111000001110010011;
ROM[724] <= 32'b00000000111000111000001110110011;
ROM[725] <= 32'b00000000011100010010000000100011;
ROM[726] <= 32'b00000000010000010000000100010011;
ROM[727] <= 32'b00000000001100010010000000100011;
ROM[728] <= 32'b00000000010000010000000100010011;
ROM[729] <= 32'b00000000010000010010000000100011;
ROM[730] <= 32'b00000000010000010000000100010011;
ROM[731] <= 32'b00000000010100010010000000100011;
ROM[732] <= 32'b00000000010000010000000100010011;
ROM[733] <= 32'b00000000011000010010000000100011;
ROM[734] <= 32'b00000000010000010000000100010011;
ROM[735] <= 32'b00000001010000000000001110010011;
ROM[736] <= 32'b00000000100000111000001110010011;
ROM[737] <= 32'b01000000011100010000001110110011;
ROM[738] <= 32'b00000000011100000000001000110011;
ROM[739] <= 32'b00000000001000000000000110110011;
ROM[740] <= 32'b00000001110000101001000011101111;
ROM[741] <= 32'b00000110001100000000001110010011;
ROM[742] <= 32'b00000000011100010010000000100011;
ROM[743] <= 32'b00000000010000010000000100010011;
ROM[744] <= 32'b00000000000000000001001110110111;
ROM[745] <= 32'b10111110110000111000001110010011;
ROM[746] <= 32'b00000000111000111000001110110011;
ROM[747] <= 32'b00000000011100010010000000100011;
ROM[748] <= 32'b00000000010000010000000100010011;
ROM[749] <= 32'b00000000001100010010000000100011;
ROM[750] <= 32'b00000000010000010000000100010011;
ROM[751] <= 32'b00000000010000010010000000100011;
ROM[752] <= 32'b00000000010000010000000100010011;
ROM[753] <= 32'b00000000010100010010000000100011;
ROM[754] <= 32'b00000000010000010000000100010011;
ROM[755] <= 32'b00000000011000010010000000100011;
ROM[756] <= 32'b00000000010000010000000100010011;
ROM[757] <= 32'b00000001010000000000001110010011;
ROM[758] <= 32'b00000000100000111000001110010011;
ROM[759] <= 32'b01000000011100010000001110110011;
ROM[760] <= 32'b00000000011100000000001000110011;
ROM[761] <= 32'b00000000001000000000000110110011;
ROM[762] <= 32'b01111100010100101000000011101111;
ROM[763] <= 32'b00000110100100000000001110010011;
ROM[764] <= 32'b00000000011100010010000000100011;
ROM[765] <= 32'b00000000010000010000000100010011;
ROM[766] <= 32'b00000000000000000001001110110111;
ROM[767] <= 32'b11000100010000111000001110010011;
ROM[768] <= 32'b00000000111000111000001110110011;
ROM[769] <= 32'b00000000011100010010000000100011;
ROM[770] <= 32'b00000000010000010000000100010011;
ROM[771] <= 32'b00000000001100010010000000100011;
ROM[772] <= 32'b00000000010000010000000100010011;
ROM[773] <= 32'b00000000010000010010000000100011;
ROM[774] <= 32'b00000000010000010000000100010011;
ROM[775] <= 32'b00000000010100010010000000100011;
ROM[776] <= 32'b00000000010000010000000100010011;
ROM[777] <= 32'b00000000011000010010000000100011;
ROM[778] <= 32'b00000000010000010000000100010011;
ROM[779] <= 32'b00000001010000000000001110010011;
ROM[780] <= 32'b00000000100000111000001110010011;
ROM[781] <= 32'b01000000011100010000001110110011;
ROM[782] <= 32'b00000000011100000000001000110011;
ROM[783] <= 32'b00000000001000000000000110110011;
ROM[784] <= 32'b01110110110100101000000011101111;
ROM[785] <= 32'b00000010000000000000001110010011;
ROM[786] <= 32'b00000000011100010010000000100011;
ROM[787] <= 32'b00000000010000010000000100010011;
ROM[788] <= 32'b00000000000000000001001110110111;
ROM[789] <= 32'b11001001110000111000001110010011;
ROM[790] <= 32'b00000000111000111000001110110011;
ROM[791] <= 32'b00000000011100010010000000100011;
ROM[792] <= 32'b00000000010000010000000100010011;
ROM[793] <= 32'b00000000001100010010000000100011;
ROM[794] <= 32'b00000000010000010000000100010011;
ROM[795] <= 32'b00000000010000010010000000100011;
ROM[796] <= 32'b00000000010000010000000100010011;
ROM[797] <= 32'b00000000010100010010000000100011;
ROM[798] <= 32'b00000000010000010000000100010011;
ROM[799] <= 32'b00000000011000010010000000100011;
ROM[800] <= 32'b00000000010000010000000100010011;
ROM[801] <= 32'b00000001010000000000001110010011;
ROM[802] <= 32'b00000000100000111000001110010011;
ROM[803] <= 32'b01000000011100010000001110110011;
ROM[804] <= 32'b00000000011100000000001000110011;
ROM[805] <= 32'b00000000001000000000000110110011;
ROM[806] <= 32'b01110001010100101000000011101111;
ROM[807] <= 32'b00000110111000000000001110010011;
ROM[808] <= 32'b00000000011100010010000000100011;
ROM[809] <= 32'b00000000010000010000000100010011;
ROM[810] <= 32'b00000000000000000001001110110111;
ROM[811] <= 32'b11001111010000111000001110010011;
ROM[812] <= 32'b00000000111000111000001110110011;
ROM[813] <= 32'b00000000011100010010000000100011;
ROM[814] <= 32'b00000000010000010000000100010011;
ROM[815] <= 32'b00000000001100010010000000100011;
ROM[816] <= 32'b00000000010000010000000100010011;
ROM[817] <= 32'b00000000010000010010000000100011;
ROM[818] <= 32'b00000000010000010000000100010011;
ROM[819] <= 32'b00000000010100010010000000100011;
ROM[820] <= 32'b00000000010000010000000100010011;
ROM[821] <= 32'b00000000011000010010000000100011;
ROM[822] <= 32'b00000000010000010000000100010011;
ROM[823] <= 32'b00000001010000000000001110010011;
ROM[824] <= 32'b00000000100000111000001110010011;
ROM[825] <= 32'b01000000011100010000001110110011;
ROM[826] <= 32'b00000000011100000000001000110011;
ROM[827] <= 32'b00000000001000000000000110110011;
ROM[828] <= 32'b01101011110100101000000011101111;
ROM[829] <= 32'b00000111010100000000001110010011;
ROM[830] <= 32'b00000000011100010010000000100011;
ROM[831] <= 32'b00000000010000010000000100010011;
ROM[832] <= 32'b00000000000000000001001110110111;
ROM[833] <= 32'b11010100110000111000001110010011;
ROM[834] <= 32'b00000000111000111000001110110011;
ROM[835] <= 32'b00000000011100010010000000100011;
ROM[836] <= 32'b00000000010000010000000100010011;
ROM[837] <= 32'b00000000001100010010000000100011;
ROM[838] <= 32'b00000000010000010000000100010011;
ROM[839] <= 32'b00000000010000010010000000100011;
ROM[840] <= 32'b00000000010000010000000100010011;
ROM[841] <= 32'b00000000010100010010000000100011;
ROM[842] <= 32'b00000000010000010000000100010011;
ROM[843] <= 32'b00000000011000010010000000100011;
ROM[844] <= 32'b00000000010000010000000100010011;
ROM[845] <= 32'b00000001010000000000001110010011;
ROM[846] <= 32'b00000000100000111000001110010011;
ROM[847] <= 32'b01000000011100010000001110110011;
ROM[848] <= 32'b00000000011100000000001000110011;
ROM[849] <= 32'b00000000001000000000000110110011;
ROM[850] <= 32'b01100110010100101000000011101111;
ROM[851] <= 32'b00000110110100000000001110010011;
ROM[852] <= 32'b00000000011100010010000000100011;
ROM[853] <= 32'b00000000010000010000000100010011;
ROM[854] <= 32'b00000000000000000001001110110111;
ROM[855] <= 32'b11011010010000111000001110010011;
ROM[856] <= 32'b00000000111000111000001110110011;
ROM[857] <= 32'b00000000011100010010000000100011;
ROM[858] <= 32'b00000000010000010000000100010011;
ROM[859] <= 32'b00000000001100010010000000100011;
ROM[860] <= 32'b00000000010000010000000100010011;
ROM[861] <= 32'b00000000010000010010000000100011;
ROM[862] <= 32'b00000000010000010000000100010011;
ROM[863] <= 32'b00000000010100010010000000100011;
ROM[864] <= 32'b00000000010000010000000100010011;
ROM[865] <= 32'b00000000011000010010000000100011;
ROM[866] <= 32'b00000000010000010000000100010011;
ROM[867] <= 32'b00000001010000000000001110010011;
ROM[868] <= 32'b00000000100000111000001110010011;
ROM[869] <= 32'b01000000011100010000001110110011;
ROM[870] <= 32'b00000000011100000000001000110011;
ROM[871] <= 32'b00000000001000000000000110110011;
ROM[872] <= 32'b01100000110100101000000011101111;
ROM[873] <= 32'b00000110001000000000001110010011;
ROM[874] <= 32'b00000000011100010010000000100011;
ROM[875] <= 32'b00000000010000010000000100010011;
ROM[876] <= 32'b00000000000000000001001110110111;
ROM[877] <= 32'b11011111110000111000001110010011;
ROM[878] <= 32'b00000000111000111000001110110011;
ROM[879] <= 32'b00000000011100010010000000100011;
ROM[880] <= 32'b00000000010000010000000100010011;
ROM[881] <= 32'b00000000001100010010000000100011;
ROM[882] <= 32'b00000000010000010000000100010011;
ROM[883] <= 32'b00000000010000010010000000100011;
ROM[884] <= 32'b00000000010000010000000100010011;
ROM[885] <= 32'b00000000010100010010000000100011;
ROM[886] <= 32'b00000000010000010000000100010011;
ROM[887] <= 32'b00000000011000010010000000100011;
ROM[888] <= 32'b00000000010000010000000100010011;
ROM[889] <= 32'b00000001010000000000001110010011;
ROM[890] <= 32'b00000000100000111000001110010011;
ROM[891] <= 32'b01000000011100010000001110110011;
ROM[892] <= 32'b00000000011100000000001000110011;
ROM[893] <= 32'b00000000001000000000000110110011;
ROM[894] <= 32'b01011011010100101000000011101111;
ROM[895] <= 32'b00000110010100000000001110010011;
ROM[896] <= 32'b00000000011100010010000000100011;
ROM[897] <= 32'b00000000010000010000000100010011;
ROM[898] <= 32'b00000000000000000001001110110111;
ROM[899] <= 32'b11100101010000111000001110010011;
ROM[900] <= 32'b00000000111000111000001110110011;
ROM[901] <= 32'b00000000011100010010000000100011;
ROM[902] <= 32'b00000000010000010000000100010011;
ROM[903] <= 32'b00000000001100010010000000100011;
ROM[904] <= 32'b00000000010000010000000100010011;
ROM[905] <= 32'b00000000010000010010000000100011;
ROM[906] <= 32'b00000000010000010000000100010011;
ROM[907] <= 32'b00000000010100010010000000100011;
ROM[908] <= 32'b00000000010000010000000100010011;
ROM[909] <= 32'b00000000011000010010000000100011;
ROM[910] <= 32'b00000000010000010000000100010011;
ROM[911] <= 32'b00000001010000000000001110010011;
ROM[912] <= 32'b00000000100000111000001110010011;
ROM[913] <= 32'b01000000011100010000001110110011;
ROM[914] <= 32'b00000000011100000000001000110011;
ROM[915] <= 32'b00000000001000000000000110110011;
ROM[916] <= 32'b01010101110100101000000011101111;
ROM[917] <= 32'b00000111001000000000001110010011;
ROM[918] <= 32'b00000000011100010010000000100011;
ROM[919] <= 32'b00000000010000010000000100010011;
ROM[920] <= 32'b00000000000000000001001110110111;
ROM[921] <= 32'b11101010110000111000001110010011;
ROM[922] <= 32'b00000000111000111000001110110011;
ROM[923] <= 32'b00000000011100010010000000100011;
ROM[924] <= 32'b00000000010000010000000100010011;
ROM[925] <= 32'b00000000001100010010000000100011;
ROM[926] <= 32'b00000000010000010000000100010011;
ROM[927] <= 32'b00000000010000010010000000100011;
ROM[928] <= 32'b00000000010000010000000100010011;
ROM[929] <= 32'b00000000010100010010000000100011;
ROM[930] <= 32'b00000000010000010000000100010011;
ROM[931] <= 32'b00000000011000010010000000100011;
ROM[932] <= 32'b00000000010000010000000100010011;
ROM[933] <= 32'b00000001010000000000001110010011;
ROM[934] <= 32'b00000000100000111000001110010011;
ROM[935] <= 32'b01000000011100010000001110110011;
ROM[936] <= 32'b00000000011100000000001000110011;
ROM[937] <= 32'b00000000001000000000000110110011;
ROM[938] <= 32'b01010000010100101000000011101111;
ROM[939] <= 32'b00000111001100000000001110010011;
ROM[940] <= 32'b00000000011100010010000000100011;
ROM[941] <= 32'b00000000010000010000000100010011;
ROM[942] <= 32'b00000000000000000001001110110111;
ROM[943] <= 32'b11110000010000111000001110010011;
ROM[944] <= 32'b00000000111000111000001110110011;
ROM[945] <= 32'b00000000011100010010000000100011;
ROM[946] <= 32'b00000000010000010000000100010011;
ROM[947] <= 32'b00000000001100010010000000100011;
ROM[948] <= 32'b00000000010000010000000100010011;
ROM[949] <= 32'b00000000010000010010000000100011;
ROM[950] <= 32'b00000000010000010000000100010011;
ROM[951] <= 32'b00000000010100010010000000100011;
ROM[952] <= 32'b00000000010000010000000100010011;
ROM[953] <= 32'b00000000011000010010000000100011;
ROM[954] <= 32'b00000000010000010000000100010011;
ROM[955] <= 32'b00000001010000000000001110010011;
ROM[956] <= 32'b00000000100000111000001110010011;
ROM[957] <= 32'b01000000011100010000001110110011;
ROM[958] <= 32'b00000000011100000000001000110011;
ROM[959] <= 32'b00000000001000000000000110110011;
ROM[960] <= 32'b01001010110100101000000011101111;
ROM[961] <= 32'b00000010000000000000001110010011;
ROM[962] <= 32'b00000000011100010010000000100011;
ROM[963] <= 32'b00000000010000010000000100010011;
ROM[964] <= 32'b00000000000000000001001110110111;
ROM[965] <= 32'b11110101110000111000001110010011;
ROM[966] <= 32'b00000000111000111000001110110011;
ROM[967] <= 32'b00000000011100010010000000100011;
ROM[968] <= 32'b00000000010000010000000100010011;
ROM[969] <= 32'b00000000001100010010000000100011;
ROM[970] <= 32'b00000000010000010000000100010011;
ROM[971] <= 32'b00000000010000010010000000100011;
ROM[972] <= 32'b00000000010000010000000100010011;
ROM[973] <= 32'b00000000010100010010000000100011;
ROM[974] <= 32'b00000000010000010000000100010011;
ROM[975] <= 32'b00000000011000010010000000100011;
ROM[976] <= 32'b00000000010000010000000100010011;
ROM[977] <= 32'b00000001010000000000001110010011;
ROM[978] <= 32'b00000000100000111000001110010011;
ROM[979] <= 32'b01000000011100010000001110110011;
ROM[980] <= 32'b00000000011100000000001000110011;
ROM[981] <= 32'b00000000001000000000000110110011;
ROM[982] <= 32'b01000101010100101000000011101111;
ROM[983] <= 32'b00000111010000000000001110010011;
ROM[984] <= 32'b00000000011100010010000000100011;
ROM[985] <= 32'b00000000010000010000000100010011;
ROM[986] <= 32'b00000000000000000001001110110111;
ROM[987] <= 32'b11111011010000111000001110010011;
ROM[988] <= 32'b00000000111000111000001110110011;
ROM[989] <= 32'b00000000011100010010000000100011;
ROM[990] <= 32'b00000000010000010000000100010011;
ROM[991] <= 32'b00000000001100010010000000100011;
ROM[992] <= 32'b00000000010000010000000100010011;
ROM[993] <= 32'b00000000010000010010000000100011;
ROM[994] <= 32'b00000000010000010000000100010011;
ROM[995] <= 32'b00000000010100010010000000100011;
ROM[996] <= 32'b00000000010000010000000100010011;
ROM[997] <= 32'b00000000011000010010000000100011;
ROM[998] <= 32'b00000000010000010000000100010011;
ROM[999] <= 32'b00000001010000000000001110010011;
ROM[1000] <= 32'b00000000100000111000001110010011;
ROM[1001] <= 32'b01000000011100010000001110110011;
ROM[1002] <= 32'b00000000011100000000001000110011;
ROM[1003] <= 32'b00000000001000000000000110110011;
ROM[1004] <= 32'b00111111110100101000000011101111;
ROM[1005] <= 32'b00000110111100000000001110010011;
ROM[1006] <= 32'b00000000011100010010000000100011;
ROM[1007] <= 32'b00000000010000010000000100010011;
ROM[1008] <= 32'b00000000000000000001001110110111;
ROM[1009] <= 32'b00000000110000111000001110010011;
ROM[1010] <= 32'b00000000111000111000001110110011;
ROM[1011] <= 32'b00000000011100010010000000100011;
ROM[1012] <= 32'b00000000010000010000000100010011;
ROM[1013] <= 32'b00000000001100010010000000100011;
ROM[1014] <= 32'b00000000010000010000000100010011;
ROM[1015] <= 32'b00000000010000010010000000100011;
ROM[1016] <= 32'b00000000010000010000000100010011;
ROM[1017] <= 32'b00000000010100010010000000100011;
ROM[1018] <= 32'b00000000010000010000000100010011;
ROM[1019] <= 32'b00000000011000010010000000100011;
ROM[1020] <= 32'b00000000010000010000000100010011;
ROM[1021] <= 32'b00000001010000000000001110010011;
ROM[1022] <= 32'b00000000100000111000001110010011;
ROM[1023] <= 32'b01000000011100010000001110110011;
ROM[1024] <= 32'b00000000011100000000001000110011;
ROM[1025] <= 32'b00000000001000000000000110110011;
ROM[1026] <= 32'b00111010010100101000000011101111;
ROM[1027] <= 32'b00000010000000000000001110010011;
ROM[1028] <= 32'b00000000011100010010000000100011;
ROM[1029] <= 32'b00000000010000010000000100010011;
ROM[1030] <= 32'b00000000000000000001001110110111;
ROM[1031] <= 32'b00000110010000111000001110010011;
ROM[1032] <= 32'b00000000111000111000001110110011;
ROM[1033] <= 32'b00000000011100010010000000100011;
ROM[1034] <= 32'b00000000010000010000000100010011;
ROM[1035] <= 32'b00000000001100010010000000100011;
ROM[1036] <= 32'b00000000010000010000000100010011;
ROM[1037] <= 32'b00000000010000010010000000100011;
ROM[1038] <= 32'b00000000010000010000000100010011;
ROM[1039] <= 32'b00000000010100010010000000100011;
ROM[1040] <= 32'b00000000010000010000000100010011;
ROM[1041] <= 32'b00000000011000010010000000100011;
ROM[1042] <= 32'b00000000010000010000000100010011;
ROM[1043] <= 32'b00000001010000000000001110010011;
ROM[1044] <= 32'b00000000100000111000001110010011;
ROM[1045] <= 32'b01000000011100010000001110110011;
ROM[1046] <= 32'b00000000011100000000001000110011;
ROM[1047] <= 32'b00000000001000000000000110110011;
ROM[1048] <= 32'b00110100110100101000000011101111;
ROM[1049] <= 32'b00000111000000000000001110010011;
ROM[1050] <= 32'b00000000011100010010000000100011;
ROM[1051] <= 32'b00000000010000010000000100010011;
ROM[1052] <= 32'b00000000000000000001001110110111;
ROM[1053] <= 32'b00001011110000111000001110010011;
ROM[1054] <= 32'b00000000111000111000001110110011;
ROM[1055] <= 32'b00000000011100010010000000100011;
ROM[1056] <= 32'b00000000010000010000000100010011;
ROM[1057] <= 32'b00000000001100010010000000100011;
ROM[1058] <= 32'b00000000010000010000000100010011;
ROM[1059] <= 32'b00000000010000010010000000100011;
ROM[1060] <= 32'b00000000010000010000000100010011;
ROM[1061] <= 32'b00000000010100010010000000100011;
ROM[1062] <= 32'b00000000010000010000000100010011;
ROM[1063] <= 32'b00000000011000010010000000100011;
ROM[1064] <= 32'b00000000010000010000000100010011;
ROM[1065] <= 32'b00000001010000000000001110010011;
ROM[1066] <= 32'b00000000100000111000001110010011;
ROM[1067] <= 32'b01000000011100010000001110110011;
ROM[1068] <= 32'b00000000011100000000001000110011;
ROM[1069] <= 32'b00000000001000000000000110110011;
ROM[1070] <= 32'b00101111010100101000000011101111;
ROM[1071] <= 32'b00000111001000000000001110010011;
ROM[1072] <= 32'b00000000011100010010000000100011;
ROM[1073] <= 32'b00000000010000010000000100010011;
ROM[1074] <= 32'b00000000000000000001001110110111;
ROM[1075] <= 32'b00010001010000111000001110010011;
ROM[1076] <= 32'b00000000111000111000001110110011;
ROM[1077] <= 32'b00000000011100010010000000100011;
ROM[1078] <= 32'b00000000010000010000000100010011;
ROM[1079] <= 32'b00000000001100010010000000100011;
ROM[1080] <= 32'b00000000010000010000000100010011;
ROM[1081] <= 32'b00000000010000010010000000100011;
ROM[1082] <= 32'b00000000010000010000000100010011;
ROM[1083] <= 32'b00000000010100010010000000100011;
ROM[1084] <= 32'b00000000010000010000000100010011;
ROM[1085] <= 32'b00000000011000010010000000100011;
ROM[1086] <= 32'b00000000010000010000000100010011;
ROM[1087] <= 32'b00000001010000000000001110010011;
ROM[1088] <= 32'b00000000100000111000001110010011;
ROM[1089] <= 32'b01000000011100010000001110110011;
ROM[1090] <= 32'b00000000011100000000001000110011;
ROM[1091] <= 32'b00000000001000000000000110110011;
ROM[1092] <= 32'b00101001110100101000000011101111;
ROM[1093] <= 32'b00000110100100000000001110010011;
ROM[1094] <= 32'b00000000011100010010000000100011;
ROM[1095] <= 32'b00000000010000010000000100010011;
ROM[1096] <= 32'b00000000000000000001001110110111;
ROM[1097] <= 32'b00010110110000111000001110010011;
ROM[1098] <= 32'b00000000111000111000001110110011;
ROM[1099] <= 32'b00000000011100010010000000100011;
ROM[1100] <= 32'b00000000010000010000000100010011;
ROM[1101] <= 32'b00000000001100010010000000100011;
ROM[1102] <= 32'b00000000010000010000000100010011;
ROM[1103] <= 32'b00000000010000010010000000100011;
ROM[1104] <= 32'b00000000010000010000000100010011;
ROM[1105] <= 32'b00000000010100010010000000100011;
ROM[1106] <= 32'b00000000010000010000000100010011;
ROM[1107] <= 32'b00000000011000010010000000100011;
ROM[1108] <= 32'b00000000010000010000000100010011;
ROM[1109] <= 32'b00000001010000000000001110010011;
ROM[1110] <= 32'b00000000100000111000001110010011;
ROM[1111] <= 32'b01000000011100010000001110110011;
ROM[1112] <= 32'b00000000011100000000001000110011;
ROM[1113] <= 32'b00000000001000000000000110110011;
ROM[1114] <= 32'b00100100010100101000000011101111;
ROM[1115] <= 32'b00000110111000000000001110010011;
ROM[1116] <= 32'b00000000011100010010000000100011;
ROM[1117] <= 32'b00000000010000010000000100010011;
ROM[1118] <= 32'b00000000000000000001001110110111;
ROM[1119] <= 32'b00011100010000111000001110010011;
ROM[1120] <= 32'b00000000111000111000001110110011;
ROM[1121] <= 32'b00000000011100010010000000100011;
ROM[1122] <= 32'b00000000010000010000000100010011;
ROM[1123] <= 32'b00000000001100010010000000100011;
ROM[1124] <= 32'b00000000010000010000000100010011;
ROM[1125] <= 32'b00000000010000010010000000100011;
ROM[1126] <= 32'b00000000010000010000000100010011;
ROM[1127] <= 32'b00000000010100010010000000100011;
ROM[1128] <= 32'b00000000010000010000000100010011;
ROM[1129] <= 32'b00000000011000010010000000100011;
ROM[1130] <= 32'b00000000010000010000000100010011;
ROM[1131] <= 32'b00000001010000000000001110010011;
ROM[1132] <= 32'b00000000100000111000001110010011;
ROM[1133] <= 32'b01000000011100010000001110110011;
ROM[1134] <= 32'b00000000011100000000001000110011;
ROM[1135] <= 32'b00000000001000000000000110110011;
ROM[1136] <= 32'b00011110110100101000000011101111;
ROM[1137] <= 32'b00000111010000000000001110010011;
ROM[1138] <= 32'b00000000011100010010000000100011;
ROM[1139] <= 32'b00000000010000010000000100010011;
ROM[1140] <= 32'b00000000000000000001001110110111;
ROM[1141] <= 32'b00100001110000111000001110010011;
ROM[1142] <= 32'b00000000111000111000001110110011;
ROM[1143] <= 32'b00000000011100010010000000100011;
ROM[1144] <= 32'b00000000010000010000000100010011;
ROM[1145] <= 32'b00000000001100010010000000100011;
ROM[1146] <= 32'b00000000010000010000000100010011;
ROM[1147] <= 32'b00000000010000010010000000100011;
ROM[1148] <= 32'b00000000010000010000000100010011;
ROM[1149] <= 32'b00000000010100010010000000100011;
ROM[1150] <= 32'b00000000010000010000000100010011;
ROM[1151] <= 32'b00000000011000010010000000100011;
ROM[1152] <= 32'b00000000010000010000000100010011;
ROM[1153] <= 32'b00000001010000000000001110010011;
ROM[1154] <= 32'b00000000100000111000001110010011;
ROM[1155] <= 32'b01000000011100010000001110110011;
ROM[1156] <= 32'b00000000011100000000001000110011;
ROM[1157] <= 32'b00000000001000000000000110110011;
ROM[1158] <= 32'b00011001010100101000000011101111;
ROM[1159] <= 32'b00000011101000000000001110010011;
ROM[1160] <= 32'b00000000011100010010000000100011;
ROM[1161] <= 32'b00000000010000010000000100010011;
ROM[1162] <= 32'b00000000000000000001001110110111;
ROM[1163] <= 32'b00100111010000111000001110010011;
ROM[1164] <= 32'b00000000111000111000001110110011;
ROM[1165] <= 32'b00000000011100010010000000100011;
ROM[1166] <= 32'b00000000010000010000000100010011;
ROM[1167] <= 32'b00000000001100010010000000100011;
ROM[1168] <= 32'b00000000010000010000000100010011;
ROM[1169] <= 32'b00000000010000010010000000100011;
ROM[1170] <= 32'b00000000010000010000000100010011;
ROM[1171] <= 32'b00000000010100010010000000100011;
ROM[1172] <= 32'b00000000010000010000000100010011;
ROM[1173] <= 32'b00000000011000010010000000100011;
ROM[1174] <= 32'b00000000010000010000000100010011;
ROM[1175] <= 32'b00000001010000000000001110010011;
ROM[1176] <= 32'b00000000100000111000001110010011;
ROM[1177] <= 32'b01000000011100010000001110110011;
ROM[1178] <= 32'b00000000011100000000001000110011;
ROM[1179] <= 32'b00000000001000000000000110110011;
ROM[1180] <= 32'b00010011110100101000000011101111;
ROM[1181] <= 32'b00000010000000000000001110010011;
ROM[1182] <= 32'b00000000011100010010000000100011;
ROM[1183] <= 32'b00000000010000010000000100010011;
ROM[1184] <= 32'b00000000000000000001001110110111;
ROM[1185] <= 32'b00101100110000111000001110010011;
ROM[1186] <= 32'b00000000111000111000001110110011;
ROM[1187] <= 32'b00000000011100010010000000100011;
ROM[1188] <= 32'b00000000010000010000000100010011;
ROM[1189] <= 32'b00000000001100010010000000100011;
ROM[1190] <= 32'b00000000010000010000000100010011;
ROM[1191] <= 32'b00000000010000010010000000100011;
ROM[1192] <= 32'b00000000010000010000000100010011;
ROM[1193] <= 32'b00000000010100010010000000100011;
ROM[1194] <= 32'b00000000010000010000000100010011;
ROM[1195] <= 32'b00000000011000010010000000100011;
ROM[1196] <= 32'b00000000010000010000000100010011;
ROM[1197] <= 32'b00000001010000000000001110010011;
ROM[1198] <= 32'b00000000100000111000001110010011;
ROM[1199] <= 32'b01000000011100010000001110110011;
ROM[1200] <= 32'b00000000011100000000001000110011;
ROM[1201] <= 32'b00000000001000000000000110110011;
ROM[1202] <= 32'b00001110010100101000000011101111;
ROM[1203] <= 32'b00000000000000000001001110110111;
ROM[1204] <= 32'b00110001100000111000001110010011;
ROM[1205] <= 32'b00000000111000111000001110110011;
ROM[1206] <= 32'b00000000011100010010000000100011;
ROM[1207] <= 32'b00000000010000010000000100010011;
ROM[1208] <= 32'b00000000001100010010000000100011;
ROM[1209] <= 32'b00000000010000010000000100010011;
ROM[1210] <= 32'b00000000010000010010000000100011;
ROM[1211] <= 32'b00000000010000010000000100010011;
ROM[1212] <= 32'b00000000010100010010000000100011;
ROM[1213] <= 32'b00000000010000010000000100010011;
ROM[1214] <= 32'b00000000011000010010000000100011;
ROM[1215] <= 32'b00000000010000010000000100010011;
ROM[1216] <= 32'b00000001010000000000001110010011;
ROM[1217] <= 32'b00000000010000111000001110010011;
ROM[1218] <= 32'b01000000011100010000001110110011;
ROM[1219] <= 32'b00000000011100000000001000110011;
ROM[1220] <= 32'b00000000001000000000000110110011;
ROM[1221] <= 32'b01011011010100001100000011101111;
ROM[1222] <= 32'b11111111110000010000000100010011;
ROM[1223] <= 32'b00000000000000010010001110000011;
ROM[1224] <= 32'b00000000011100011010000000100011;
ROM[1225] <= 32'b00000000000000000000001110010011;
ROM[1226] <= 32'b00000000011100010010000000100011;
ROM[1227] <= 32'b00000000010000010000000100010011;
ROM[1228] <= 32'b11111111110000010000000100010011;
ROM[1229] <= 32'b00000000000000010010001110000011;
ROM[1230] <= 32'b00000000011100011010001000100011;
ROM[1231] <= 32'b00000000000100000000001110010011;
ROM[1232] <= 32'b00000000011100010010000000100011;
ROM[1233] <= 32'b00000000010000010000000100010011;
ROM[1234] <= 32'b11111111110000010000000100010011;
ROM[1235] <= 32'b00000000000000010010001110000011;
ROM[1236] <= 32'b00000000011100011010010000100011;
ROM[1237] <= 32'b00000000101000000000001110010011;
ROM[1238] <= 32'b00000000011100010010000000100011;
ROM[1239] <= 32'b00000000010000010000000100010011;
ROM[1240] <= 32'b00000000000000000001001110110111;
ROM[1241] <= 32'b00111010110000111000001110010011;
ROM[1242] <= 32'b00000000111000111000001110110011;
ROM[1243] <= 32'b00000000011100010010000000100011;
ROM[1244] <= 32'b00000000010000010000000100010011;
ROM[1245] <= 32'b00000000001100010010000000100011;
ROM[1246] <= 32'b00000000010000010000000100010011;
ROM[1247] <= 32'b00000000010000010010000000100011;
ROM[1248] <= 32'b00000000010000010000000100010011;
ROM[1249] <= 32'b00000000010100010010000000100011;
ROM[1250] <= 32'b00000000010000010000000100010011;
ROM[1251] <= 32'b00000000011000010010000000100011;
ROM[1252] <= 32'b00000000010000010000000100010011;
ROM[1253] <= 32'b00000001010000000000001110010011;
ROM[1254] <= 32'b00000000010000111000001110010011;
ROM[1255] <= 32'b01000000011100010000001110110011;
ROM[1256] <= 32'b00000000011100000000001000110011;
ROM[1257] <= 32'b00000000001000000000000110110011;
ROM[1258] <= 32'b00111001010000101000000011101111;
ROM[1259] <= 32'b00000101010000000000001110010011;
ROM[1260] <= 32'b00000000011100010010000000100011;
ROM[1261] <= 32'b00000000010000010000000100010011;
ROM[1262] <= 32'b00000000000000000001001110110111;
ROM[1263] <= 32'b01000000010000111000001110010011;
ROM[1264] <= 32'b00000000111000111000001110110011;
ROM[1265] <= 32'b00000000011100010010000000100011;
ROM[1266] <= 32'b00000000010000010000000100010011;
ROM[1267] <= 32'b00000000001100010010000000100011;
ROM[1268] <= 32'b00000000010000010000000100010011;
ROM[1269] <= 32'b00000000010000010010000000100011;
ROM[1270] <= 32'b00000000010000010000000100010011;
ROM[1271] <= 32'b00000000010100010010000000100011;
ROM[1272] <= 32'b00000000010000010000000100010011;
ROM[1273] <= 32'b00000000011000010010000000100011;
ROM[1274] <= 32'b00000000010000010000000100010011;
ROM[1275] <= 32'b00000001010000000000001110010011;
ROM[1276] <= 32'b00000000100000111000001110010011;
ROM[1277] <= 32'b01000000011100010000001110110011;
ROM[1278] <= 32'b00000000011100000000001000110011;
ROM[1279] <= 32'b00000000001000000000000110110011;
ROM[1280] <= 32'b01111010110000101000000011101111;
ROM[1281] <= 32'b00000110100000000000001110010011;
ROM[1282] <= 32'b00000000011100010010000000100011;
ROM[1283] <= 32'b00000000010000010000000100010011;
ROM[1284] <= 32'b00000000000000000001001110110111;
ROM[1285] <= 32'b01000101110000111000001110010011;
ROM[1286] <= 32'b00000000111000111000001110110011;
ROM[1287] <= 32'b00000000011100010010000000100011;
ROM[1288] <= 32'b00000000010000010000000100010011;
ROM[1289] <= 32'b00000000001100010010000000100011;
ROM[1290] <= 32'b00000000010000010000000100010011;
ROM[1291] <= 32'b00000000010000010010000000100011;
ROM[1292] <= 32'b00000000010000010000000100010011;
ROM[1293] <= 32'b00000000010100010010000000100011;
ROM[1294] <= 32'b00000000010000010000000100010011;
ROM[1295] <= 32'b00000000011000010010000000100011;
ROM[1296] <= 32'b00000000010000010000000100010011;
ROM[1297] <= 32'b00000001010000000000001110010011;
ROM[1298] <= 32'b00000000100000111000001110010011;
ROM[1299] <= 32'b01000000011100010000001110110011;
ROM[1300] <= 32'b00000000011100000000001000110011;
ROM[1301] <= 32'b00000000001000000000000110110011;
ROM[1302] <= 32'b01110101010000101000000011101111;
ROM[1303] <= 32'b00000110010100000000001110010011;
ROM[1304] <= 32'b00000000011100010010000000100011;
ROM[1305] <= 32'b00000000010000010000000100010011;
ROM[1306] <= 32'b00000000000000000001001110110111;
ROM[1307] <= 32'b01001011010000111000001110010011;
ROM[1308] <= 32'b00000000111000111000001110110011;
ROM[1309] <= 32'b00000000011100010010000000100011;
ROM[1310] <= 32'b00000000010000010000000100010011;
ROM[1311] <= 32'b00000000001100010010000000100011;
ROM[1312] <= 32'b00000000010000010000000100010011;
ROM[1313] <= 32'b00000000010000010010000000100011;
ROM[1314] <= 32'b00000000010000010000000100010011;
ROM[1315] <= 32'b00000000010100010010000000100011;
ROM[1316] <= 32'b00000000010000010000000100010011;
ROM[1317] <= 32'b00000000011000010010000000100011;
ROM[1318] <= 32'b00000000010000010000000100010011;
ROM[1319] <= 32'b00000001010000000000001110010011;
ROM[1320] <= 32'b00000000100000111000001110010011;
ROM[1321] <= 32'b01000000011100010000001110110011;
ROM[1322] <= 32'b00000000011100000000001000110011;
ROM[1323] <= 32'b00000000001000000000000110110011;
ROM[1324] <= 32'b01101111110000101000000011101111;
ROM[1325] <= 32'b00000010000000000000001110010011;
ROM[1326] <= 32'b00000000011100010010000000100011;
ROM[1327] <= 32'b00000000010000010000000100010011;
ROM[1328] <= 32'b00000000000000000001001110110111;
ROM[1329] <= 32'b01010000110000111000001110010011;
ROM[1330] <= 32'b00000000111000111000001110110011;
ROM[1331] <= 32'b00000000011100010010000000100011;
ROM[1332] <= 32'b00000000010000010000000100010011;
ROM[1333] <= 32'b00000000001100010010000000100011;
ROM[1334] <= 32'b00000000010000010000000100010011;
ROM[1335] <= 32'b00000000010000010010000000100011;
ROM[1336] <= 32'b00000000010000010000000100010011;
ROM[1337] <= 32'b00000000010100010010000000100011;
ROM[1338] <= 32'b00000000010000010000000100010011;
ROM[1339] <= 32'b00000000011000010010000000100011;
ROM[1340] <= 32'b00000000010000010000000100010011;
ROM[1341] <= 32'b00000001010000000000001110010011;
ROM[1342] <= 32'b00000000100000111000001110010011;
ROM[1343] <= 32'b01000000011100010000001110110011;
ROM[1344] <= 32'b00000000011100000000001000110011;
ROM[1345] <= 32'b00000000001000000000000110110011;
ROM[1346] <= 32'b01101010010000101000000011101111;
ROM[1347] <= 32'b00000110011000000000001110010011;
ROM[1348] <= 32'b00000000011100010010000000100011;
ROM[1349] <= 32'b00000000010000010000000100010011;
ROM[1350] <= 32'b00000000000000000001001110110111;
ROM[1351] <= 32'b01010110010000111000001110010011;
ROM[1352] <= 32'b00000000111000111000001110110011;
ROM[1353] <= 32'b00000000011100010010000000100011;
ROM[1354] <= 32'b00000000010000010000000100010011;
ROM[1355] <= 32'b00000000001100010010000000100011;
ROM[1356] <= 32'b00000000010000010000000100010011;
ROM[1357] <= 32'b00000000010000010010000000100011;
ROM[1358] <= 32'b00000000010000010000000100010011;
ROM[1359] <= 32'b00000000010100010010000000100011;
ROM[1360] <= 32'b00000000010000010000000100010011;
ROM[1361] <= 32'b00000000011000010010000000100011;
ROM[1362] <= 32'b00000000010000010000000100010011;
ROM[1363] <= 32'b00000001010000000000001110010011;
ROM[1364] <= 32'b00000000100000111000001110010011;
ROM[1365] <= 32'b01000000011100010000001110110011;
ROM[1366] <= 32'b00000000011100000000001000110011;
ROM[1367] <= 32'b00000000001000000000000110110011;
ROM[1368] <= 32'b01100100110000101000000011101111;
ROM[1369] <= 32'b00000110100100000000001110010011;
ROM[1370] <= 32'b00000000011100010010000000100011;
ROM[1371] <= 32'b00000000010000010000000100010011;
ROM[1372] <= 32'b00000000000000000001001110110111;
ROM[1373] <= 32'b01011011110000111000001110010011;
ROM[1374] <= 32'b00000000111000111000001110110011;
ROM[1375] <= 32'b00000000011100010010000000100011;
ROM[1376] <= 32'b00000000010000010000000100010011;
ROM[1377] <= 32'b00000000001100010010000000100011;
ROM[1378] <= 32'b00000000010000010000000100010011;
ROM[1379] <= 32'b00000000010000010010000000100011;
ROM[1380] <= 32'b00000000010000010000000100010011;
ROM[1381] <= 32'b00000000010100010010000000100011;
ROM[1382] <= 32'b00000000010000010000000100010011;
ROM[1383] <= 32'b00000000011000010010000000100011;
ROM[1384] <= 32'b00000000010000010000000100010011;
ROM[1385] <= 32'b00000001010000000000001110010011;
ROM[1386] <= 32'b00000000100000111000001110010011;
ROM[1387] <= 32'b01000000011100010000001110110011;
ROM[1388] <= 32'b00000000011100000000001000110011;
ROM[1389] <= 32'b00000000001000000000000110110011;
ROM[1390] <= 32'b01011111010000101000000011101111;
ROM[1391] <= 32'b00000111001000000000001110010011;
ROM[1392] <= 32'b00000000011100010010000000100011;
ROM[1393] <= 32'b00000000010000010000000100010011;
ROM[1394] <= 32'b00000000000000000001001110110111;
ROM[1395] <= 32'b01100001010000111000001110010011;
ROM[1396] <= 32'b00000000111000111000001110110011;
ROM[1397] <= 32'b00000000011100010010000000100011;
ROM[1398] <= 32'b00000000010000010000000100010011;
ROM[1399] <= 32'b00000000001100010010000000100011;
ROM[1400] <= 32'b00000000010000010000000100010011;
ROM[1401] <= 32'b00000000010000010010000000100011;
ROM[1402] <= 32'b00000000010000010000000100010011;
ROM[1403] <= 32'b00000000010100010010000000100011;
ROM[1404] <= 32'b00000000010000010000000100010011;
ROM[1405] <= 32'b00000000011000010010000000100011;
ROM[1406] <= 32'b00000000010000010000000100010011;
ROM[1407] <= 32'b00000001010000000000001110010011;
ROM[1408] <= 32'b00000000100000111000001110010011;
ROM[1409] <= 32'b01000000011100010000001110110011;
ROM[1410] <= 32'b00000000011100000000001000110011;
ROM[1411] <= 32'b00000000001000000000000110110011;
ROM[1412] <= 32'b01011001110000101000000011101111;
ROM[1413] <= 32'b00000111001100000000001110010011;
ROM[1414] <= 32'b00000000011100010010000000100011;
ROM[1415] <= 32'b00000000010000010000000100010011;
ROM[1416] <= 32'b00000000000000000001001110110111;
ROM[1417] <= 32'b01100110110000111000001110010011;
ROM[1418] <= 32'b00000000111000111000001110110011;
ROM[1419] <= 32'b00000000011100010010000000100011;
ROM[1420] <= 32'b00000000010000010000000100010011;
ROM[1421] <= 32'b00000000001100010010000000100011;
ROM[1422] <= 32'b00000000010000010000000100010011;
ROM[1423] <= 32'b00000000010000010010000000100011;
ROM[1424] <= 32'b00000000010000010000000100010011;
ROM[1425] <= 32'b00000000010100010010000000100011;
ROM[1426] <= 32'b00000000010000010000000100010011;
ROM[1427] <= 32'b00000000011000010010000000100011;
ROM[1428] <= 32'b00000000010000010000000100010011;
ROM[1429] <= 32'b00000001010000000000001110010011;
ROM[1430] <= 32'b00000000100000111000001110010011;
ROM[1431] <= 32'b01000000011100010000001110110011;
ROM[1432] <= 32'b00000000011100000000001000110011;
ROM[1433] <= 32'b00000000001000000000000110110011;
ROM[1434] <= 32'b01010100010000101000000011101111;
ROM[1435] <= 32'b00000111010000000000001110010011;
ROM[1436] <= 32'b00000000011100010010000000100011;
ROM[1437] <= 32'b00000000010000010000000100010011;
ROM[1438] <= 32'b00000000000000000001001110110111;
ROM[1439] <= 32'b01101100010000111000001110010011;
ROM[1440] <= 32'b00000000111000111000001110110011;
ROM[1441] <= 32'b00000000011100010010000000100011;
ROM[1442] <= 32'b00000000010000010000000100010011;
ROM[1443] <= 32'b00000000001100010010000000100011;
ROM[1444] <= 32'b00000000010000010000000100010011;
ROM[1445] <= 32'b00000000010000010010000000100011;
ROM[1446] <= 32'b00000000010000010000000100010011;
ROM[1447] <= 32'b00000000010100010010000000100011;
ROM[1448] <= 32'b00000000010000010000000100010011;
ROM[1449] <= 32'b00000000011000010010000000100011;
ROM[1450] <= 32'b00000000010000010000000100010011;
ROM[1451] <= 32'b00000001010000000000001110010011;
ROM[1452] <= 32'b00000000100000111000001110010011;
ROM[1453] <= 32'b01000000011100010000001110110011;
ROM[1454] <= 32'b00000000011100000000001000110011;
ROM[1455] <= 32'b00000000001000000000000110110011;
ROM[1456] <= 32'b01001110110000101000000011101111;
ROM[1457] <= 32'b00000010000000000000001110010011;
ROM[1458] <= 32'b00000000011100010010000000100011;
ROM[1459] <= 32'b00000000010000010000000100010011;
ROM[1460] <= 32'b00000000000000000001001110110111;
ROM[1461] <= 32'b01110001110000111000001110010011;
ROM[1462] <= 32'b00000000111000111000001110110011;
ROM[1463] <= 32'b00000000011100010010000000100011;
ROM[1464] <= 32'b00000000010000010000000100010011;
ROM[1465] <= 32'b00000000001100010010000000100011;
ROM[1466] <= 32'b00000000010000010000000100010011;
ROM[1467] <= 32'b00000000010000010010000000100011;
ROM[1468] <= 32'b00000000010000010000000100010011;
ROM[1469] <= 32'b00000000010100010010000000100011;
ROM[1470] <= 32'b00000000010000010000000100010011;
ROM[1471] <= 32'b00000000011000010010000000100011;
ROM[1472] <= 32'b00000000010000010000000100010011;
ROM[1473] <= 32'b00000001010000000000001110010011;
ROM[1474] <= 32'b00000000100000111000001110010011;
ROM[1475] <= 32'b01000000011100010000001110110011;
ROM[1476] <= 32'b00000000011100000000001000110011;
ROM[1477] <= 32'b00000000001000000000000110110011;
ROM[1478] <= 32'b01001001010000101000000011101111;
ROM[1479] <= 32'b00000000000000000001001110110111;
ROM[1480] <= 32'b01110110100000111000001110010011;
ROM[1481] <= 32'b00000000111000111000001110110011;
ROM[1482] <= 32'b00000000011100010010000000100011;
ROM[1483] <= 32'b00000000010000010000000100010011;
ROM[1484] <= 32'b00000000001100010010000000100011;
ROM[1485] <= 32'b00000000010000010000000100010011;
ROM[1486] <= 32'b00000000010000010010000000100011;
ROM[1487] <= 32'b00000000010000010000000100010011;
ROM[1488] <= 32'b00000000010100010010000000100011;
ROM[1489] <= 32'b00000000010000010000000100010011;
ROM[1490] <= 32'b00000000011000010010000000100011;
ROM[1491] <= 32'b00000000010000010000000100010011;
ROM[1492] <= 32'b00000001010000000000001110010011;
ROM[1493] <= 32'b00000000010000111000001110010011;
ROM[1494] <= 32'b01000000011100010000001110110011;
ROM[1495] <= 32'b00000000011100000000001000110011;
ROM[1496] <= 32'b00000000001000000000000110110011;
ROM[1497] <= 32'b00000000010100010101000011101111;
ROM[1498] <= 32'b11111111110000010000000100010011;
ROM[1499] <= 32'b00000000000000010010001110000011;
ROM[1500] <= 32'b00000000011101100010000000100011;
ROM[1501] <= 32'b00000000000000011010001110000011;
ROM[1502] <= 32'b00000000011100010010000000100011;
ROM[1503] <= 32'b00000000010000010000000100010011;
ROM[1504] <= 32'b00000000000000000001001110110111;
ROM[1505] <= 32'b01111100110000111000001110010011;
ROM[1506] <= 32'b00000000111000111000001110110011;
ROM[1507] <= 32'b00000000011100010010000000100011;
ROM[1508] <= 32'b00000000010000010000000100010011;
ROM[1509] <= 32'b00000000001100010010000000100011;
ROM[1510] <= 32'b00000000010000010000000100010011;
ROM[1511] <= 32'b00000000010000010010000000100011;
ROM[1512] <= 32'b00000000010000010000000100010011;
ROM[1513] <= 32'b00000000010100010010000000100011;
ROM[1514] <= 32'b00000000010000010000000100010011;
ROM[1515] <= 32'b00000000011000010010000000100011;
ROM[1516] <= 32'b00000000010000010000000100010011;
ROM[1517] <= 32'b00000001010000000000001110010011;
ROM[1518] <= 32'b00000000010000111000001110010011;
ROM[1519] <= 32'b01000000011100010000001110110011;
ROM[1520] <= 32'b00000000011100000000001000110011;
ROM[1521] <= 32'b00000000001000000000000110110011;
ROM[1522] <= 32'b00011011100100010101000011101111;
ROM[1523] <= 32'b11111111110000010000000100010011;
ROM[1524] <= 32'b00000000000000010010001110000011;
ROM[1525] <= 32'b00000000011101100010000000100011;
ROM[1526] <= 32'b00000001100000000000001110010011;
ROM[1527] <= 32'b00000000011100010010000000100011;
ROM[1528] <= 32'b00000000010000010000000100010011;
ROM[1529] <= 32'b00000000000000000010001110110111;
ROM[1530] <= 32'b10000011000000111000001110010011;
ROM[1531] <= 32'b00000000111000111000001110110011;
ROM[1532] <= 32'b00000000011100010010000000100011;
ROM[1533] <= 32'b00000000010000010000000100010011;
ROM[1534] <= 32'b00000000001100010010000000100011;
ROM[1535] <= 32'b00000000010000010000000100010011;
ROM[1536] <= 32'b00000000010000010010000000100011;
ROM[1537] <= 32'b00000000010000010000000100010011;
ROM[1538] <= 32'b00000000010100010010000000100011;
ROM[1539] <= 32'b00000000010000010000000100010011;
ROM[1540] <= 32'b00000000011000010010000000100011;
ROM[1541] <= 32'b00000000010000010000000100010011;
ROM[1542] <= 32'b00000001010000000000001110010011;
ROM[1543] <= 32'b00000000010000111000001110010011;
ROM[1544] <= 32'b01000000011100010000001110110011;
ROM[1545] <= 32'b00000000011100000000001000110011;
ROM[1546] <= 32'b00000000001000000000000110110011;
ROM[1547] <= 32'b01110001000100100111000011101111;
ROM[1548] <= 32'b00000010000000000000001110010011;
ROM[1549] <= 32'b00000000011100010010000000100011;
ROM[1550] <= 32'b00000000010000010000000100010011;
ROM[1551] <= 32'b00000000000000000010001110110111;
ROM[1552] <= 32'b10001000100000111000001110010011;
ROM[1553] <= 32'b00000000111000111000001110110011;
ROM[1554] <= 32'b00000000011100010010000000100011;
ROM[1555] <= 32'b00000000010000010000000100010011;
ROM[1556] <= 32'b00000000001100010010000000100011;
ROM[1557] <= 32'b00000000010000010000000100010011;
ROM[1558] <= 32'b00000000010000010010000000100011;
ROM[1559] <= 32'b00000000010000010000000100010011;
ROM[1560] <= 32'b00000000010100010010000000100011;
ROM[1561] <= 32'b00000000010000010000000100010011;
ROM[1562] <= 32'b00000000011000010010000000100011;
ROM[1563] <= 32'b00000000010000010000000100010011;
ROM[1564] <= 32'b00000001010000000000001110010011;
ROM[1565] <= 32'b00000000100000111000001110010011;
ROM[1566] <= 32'b01000000011100010000001110110011;
ROM[1567] <= 32'b00000000011100000000001000110011;
ROM[1568] <= 32'b00000000001000000000000110110011;
ROM[1569] <= 32'b00110010100000101000000011101111;
ROM[1570] <= 32'b00000100011000000000001110010011;
ROM[1571] <= 32'b00000000011100010010000000100011;
ROM[1572] <= 32'b00000000010000010000000100010011;
ROM[1573] <= 32'b00000000000000000010001110110111;
ROM[1574] <= 32'b10001110000000111000001110010011;
ROM[1575] <= 32'b00000000111000111000001110110011;
ROM[1576] <= 32'b00000000011100010010000000100011;
ROM[1577] <= 32'b00000000010000010000000100010011;
ROM[1578] <= 32'b00000000001100010010000000100011;
ROM[1579] <= 32'b00000000010000010000000100010011;
ROM[1580] <= 32'b00000000010000010010000000100011;
ROM[1581] <= 32'b00000000010000010000000100010011;
ROM[1582] <= 32'b00000000010100010010000000100011;
ROM[1583] <= 32'b00000000010000010000000100010011;
ROM[1584] <= 32'b00000000011000010010000000100011;
ROM[1585] <= 32'b00000000010000010000000100010011;
ROM[1586] <= 32'b00000001010000000000001110010011;
ROM[1587] <= 32'b00000000100000111000001110010011;
ROM[1588] <= 32'b01000000011100010000001110110011;
ROM[1589] <= 32'b00000000011100000000001000110011;
ROM[1590] <= 32'b00000000001000000000000110110011;
ROM[1591] <= 32'b00101101000000101000000011101111;
ROM[1592] <= 32'b00000110100100000000001110010011;
ROM[1593] <= 32'b00000000011100010010000000100011;
ROM[1594] <= 32'b00000000010000010000000100010011;
ROM[1595] <= 32'b00000000000000000010001110110111;
ROM[1596] <= 32'b10010011100000111000001110010011;
ROM[1597] <= 32'b00000000111000111000001110110011;
ROM[1598] <= 32'b00000000011100010010000000100011;
ROM[1599] <= 32'b00000000010000010000000100010011;
ROM[1600] <= 32'b00000000001100010010000000100011;
ROM[1601] <= 32'b00000000010000010000000100010011;
ROM[1602] <= 32'b00000000010000010010000000100011;
ROM[1603] <= 32'b00000000010000010000000100010011;
ROM[1604] <= 32'b00000000010100010010000000100011;
ROM[1605] <= 32'b00000000010000010000000100010011;
ROM[1606] <= 32'b00000000011000010010000000100011;
ROM[1607] <= 32'b00000000010000010000000100010011;
ROM[1608] <= 32'b00000001010000000000001110010011;
ROM[1609] <= 32'b00000000100000111000001110010011;
ROM[1610] <= 32'b01000000011100010000001110110011;
ROM[1611] <= 32'b00000000011100000000001000110011;
ROM[1612] <= 32'b00000000001000000000000110110011;
ROM[1613] <= 32'b00100111100000101000000011101111;
ROM[1614] <= 32'b00000110001000000000001110010011;
ROM[1615] <= 32'b00000000011100010010000000100011;
ROM[1616] <= 32'b00000000010000010000000100010011;
ROM[1617] <= 32'b00000000000000000010001110110111;
ROM[1618] <= 32'b10011001000000111000001110010011;
ROM[1619] <= 32'b00000000111000111000001110110011;
ROM[1620] <= 32'b00000000011100010010000000100011;
ROM[1621] <= 32'b00000000010000010000000100010011;
ROM[1622] <= 32'b00000000001100010010000000100011;
ROM[1623] <= 32'b00000000010000010000000100010011;
ROM[1624] <= 32'b00000000010000010010000000100011;
ROM[1625] <= 32'b00000000010000010000000100010011;
ROM[1626] <= 32'b00000000010100010010000000100011;
ROM[1627] <= 32'b00000000010000010000000100010011;
ROM[1628] <= 32'b00000000011000010010000000100011;
ROM[1629] <= 32'b00000000010000010000000100010011;
ROM[1630] <= 32'b00000001010000000000001110010011;
ROM[1631] <= 32'b00000000100000111000001110010011;
ROM[1632] <= 32'b01000000011100010000001110110011;
ROM[1633] <= 32'b00000000011100000000001000110011;
ROM[1634] <= 32'b00000000001000000000000110110011;
ROM[1635] <= 32'b00100010000000101000000011101111;
ROM[1636] <= 32'b00000110111100000000001110010011;
ROM[1637] <= 32'b00000000011100010010000000100011;
ROM[1638] <= 32'b00000000010000010000000100010011;
ROM[1639] <= 32'b00000000000000000010001110110111;
ROM[1640] <= 32'b10011110100000111000001110010011;
ROM[1641] <= 32'b00000000111000111000001110110011;
ROM[1642] <= 32'b00000000011100010010000000100011;
ROM[1643] <= 32'b00000000010000010000000100010011;
ROM[1644] <= 32'b00000000001100010010000000100011;
ROM[1645] <= 32'b00000000010000010000000100010011;
ROM[1646] <= 32'b00000000010000010010000000100011;
ROM[1647] <= 32'b00000000010000010000000100010011;
ROM[1648] <= 32'b00000000010100010010000000100011;
ROM[1649] <= 32'b00000000010000010000000100010011;
ROM[1650] <= 32'b00000000011000010010000000100011;
ROM[1651] <= 32'b00000000010000010000000100010011;
ROM[1652] <= 32'b00000001010000000000001110010011;
ROM[1653] <= 32'b00000000100000111000001110010011;
ROM[1654] <= 32'b01000000011100010000001110110011;
ROM[1655] <= 32'b00000000011100000000001000110011;
ROM[1656] <= 32'b00000000001000000000000110110011;
ROM[1657] <= 32'b00011100100000101000000011101111;
ROM[1658] <= 32'b00000110111000000000001110010011;
ROM[1659] <= 32'b00000000011100010010000000100011;
ROM[1660] <= 32'b00000000010000010000000100010011;
ROM[1661] <= 32'b00000000000000000010001110110111;
ROM[1662] <= 32'b10100100000000111000001110010011;
ROM[1663] <= 32'b00000000111000111000001110110011;
ROM[1664] <= 32'b00000000011100010010000000100011;
ROM[1665] <= 32'b00000000010000010000000100010011;
ROM[1666] <= 32'b00000000001100010010000000100011;
ROM[1667] <= 32'b00000000010000010000000100010011;
ROM[1668] <= 32'b00000000010000010010000000100011;
ROM[1669] <= 32'b00000000010000010000000100010011;
ROM[1670] <= 32'b00000000010100010010000000100011;
ROM[1671] <= 32'b00000000010000010000000100010011;
ROM[1672] <= 32'b00000000011000010010000000100011;
ROM[1673] <= 32'b00000000010000010000000100010011;
ROM[1674] <= 32'b00000001010000000000001110010011;
ROM[1675] <= 32'b00000000100000111000001110010011;
ROM[1676] <= 32'b01000000011100010000001110110011;
ROM[1677] <= 32'b00000000011100000000001000110011;
ROM[1678] <= 32'b00000000001000000000000110110011;
ROM[1679] <= 32'b00010111000000101000000011101111;
ROM[1680] <= 32'b00000110000100000000001110010011;
ROM[1681] <= 32'b00000000011100010010000000100011;
ROM[1682] <= 32'b00000000010000010000000100010011;
ROM[1683] <= 32'b00000000000000000010001110110111;
ROM[1684] <= 32'b10101001100000111000001110010011;
ROM[1685] <= 32'b00000000111000111000001110110011;
ROM[1686] <= 32'b00000000011100010010000000100011;
ROM[1687] <= 32'b00000000010000010000000100010011;
ROM[1688] <= 32'b00000000001100010010000000100011;
ROM[1689] <= 32'b00000000010000010000000100010011;
ROM[1690] <= 32'b00000000010000010010000000100011;
ROM[1691] <= 32'b00000000010000010000000100010011;
ROM[1692] <= 32'b00000000010100010010000000100011;
ROM[1693] <= 32'b00000000010000010000000100010011;
ROM[1694] <= 32'b00000000011000010010000000100011;
ROM[1695] <= 32'b00000000010000010000000100010011;
ROM[1696] <= 32'b00000001010000000000001110010011;
ROM[1697] <= 32'b00000000100000111000001110010011;
ROM[1698] <= 32'b01000000011100010000001110110011;
ROM[1699] <= 32'b00000000011100000000001000110011;
ROM[1700] <= 32'b00000000001000000000000110110011;
ROM[1701] <= 32'b00010001100000101000000011101111;
ROM[1702] <= 32'b00000110001100000000001110010011;
ROM[1703] <= 32'b00000000011100010010000000100011;
ROM[1704] <= 32'b00000000010000010000000100010011;
ROM[1705] <= 32'b00000000000000000010001110110111;
ROM[1706] <= 32'b10101111000000111000001110010011;
ROM[1707] <= 32'b00000000111000111000001110110011;
ROM[1708] <= 32'b00000000011100010010000000100011;
ROM[1709] <= 32'b00000000010000010000000100010011;
ROM[1710] <= 32'b00000000001100010010000000100011;
ROM[1711] <= 32'b00000000010000010000000100010011;
ROM[1712] <= 32'b00000000010000010010000000100011;
ROM[1713] <= 32'b00000000010000010000000100010011;
ROM[1714] <= 32'b00000000010100010010000000100011;
ROM[1715] <= 32'b00000000010000010000000100010011;
ROM[1716] <= 32'b00000000011000010010000000100011;
ROM[1717] <= 32'b00000000010000010000000100010011;
ROM[1718] <= 32'b00000001010000000000001110010011;
ROM[1719] <= 32'b00000000100000111000001110010011;
ROM[1720] <= 32'b01000000011100010000001110110011;
ROM[1721] <= 32'b00000000011100000000001000110011;
ROM[1722] <= 32'b00000000001000000000000110110011;
ROM[1723] <= 32'b00001100000000101000000011101111;
ROM[1724] <= 32'b00000110001100000000001110010011;
ROM[1725] <= 32'b00000000011100010010000000100011;
ROM[1726] <= 32'b00000000010000010000000100010011;
ROM[1727] <= 32'b00000000000000000010001110110111;
ROM[1728] <= 32'b10110100100000111000001110010011;
ROM[1729] <= 32'b00000000111000111000001110110011;
ROM[1730] <= 32'b00000000011100010010000000100011;
ROM[1731] <= 32'b00000000010000010000000100010011;
ROM[1732] <= 32'b00000000001100010010000000100011;
ROM[1733] <= 32'b00000000010000010000000100010011;
ROM[1734] <= 32'b00000000010000010010000000100011;
ROM[1735] <= 32'b00000000010000010000000100010011;
ROM[1736] <= 32'b00000000010100010010000000100011;
ROM[1737] <= 32'b00000000010000010000000100010011;
ROM[1738] <= 32'b00000000011000010010000000100011;
ROM[1739] <= 32'b00000000010000010000000100010011;
ROM[1740] <= 32'b00000001010000000000001110010011;
ROM[1741] <= 32'b00000000100000111000001110010011;
ROM[1742] <= 32'b01000000011100010000001110110011;
ROM[1743] <= 32'b00000000011100000000001000110011;
ROM[1744] <= 32'b00000000001000000000000110110011;
ROM[1745] <= 32'b00000110100000101000000011101111;
ROM[1746] <= 32'b00000110100100000000001110010011;
ROM[1747] <= 32'b00000000011100010010000000100011;
ROM[1748] <= 32'b00000000010000010000000100010011;
ROM[1749] <= 32'b00000000000000000010001110110111;
ROM[1750] <= 32'b10111010000000111000001110010011;
ROM[1751] <= 32'b00000000111000111000001110110011;
ROM[1752] <= 32'b00000000011100010010000000100011;
ROM[1753] <= 32'b00000000010000010000000100010011;
ROM[1754] <= 32'b00000000001100010010000000100011;
ROM[1755] <= 32'b00000000010000010000000100010011;
ROM[1756] <= 32'b00000000010000010010000000100011;
ROM[1757] <= 32'b00000000010000010000000100010011;
ROM[1758] <= 32'b00000000010100010010000000100011;
ROM[1759] <= 32'b00000000010000010000000100010011;
ROM[1760] <= 32'b00000000011000010010000000100011;
ROM[1761] <= 32'b00000000010000010000000100010011;
ROM[1762] <= 32'b00000001010000000000001110010011;
ROM[1763] <= 32'b00000000100000111000001110010011;
ROM[1764] <= 32'b01000000011100010000001110110011;
ROM[1765] <= 32'b00000000011100000000001000110011;
ROM[1766] <= 32'b00000000001000000000000110110011;
ROM[1767] <= 32'b00000001000000101000000011101111;
ROM[1768] <= 32'b00000010000000000000001110010011;
ROM[1769] <= 32'b00000000011100010010000000100011;
ROM[1770] <= 32'b00000000010000010000000100010011;
ROM[1771] <= 32'b00000000000000000010001110110111;
ROM[1772] <= 32'b10111111100000111000001110010011;
ROM[1773] <= 32'b00000000111000111000001110110011;
ROM[1774] <= 32'b00000000011100010010000000100011;
ROM[1775] <= 32'b00000000010000010000000100010011;
ROM[1776] <= 32'b00000000001100010010000000100011;
ROM[1777] <= 32'b00000000010000010000000100010011;
ROM[1778] <= 32'b00000000010000010010000000100011;
ROM[1779] <= 32'b00000000010000010000000100010011;
ROM[1780] <= 32'b00000000010100010010000000100011;
ROM[1781] <= 32'b00000000010000010000000100010011;
ROM[1782] <= 32'b00000000011000010010000000100011;
ROM[1783] <= 32'b00000000010000010000000100010011;
ROM[1784] <= 32'b00000001010000000000001110010011;
ROM[1785] <= 32'b00000000100000111000001110010011;
ROM[1786] <= 32'b01000000011100010000001110110011;
ROM[1787] <= 32'b00000000011100000000001000110011;
ROM[1788] <= 32'b00000000001000000000000110110011;
ROM[1789] <= 32'b01111011100100100111000011101111;
ROM[1790] <= 32'b00000110111000000000001110010011;
ROM[1791] <= 32'b00000000011100010010000000100011;
ROM[1792] <= 32'b00000000010000010000000100010011;
ROM[1793] <= 32'b00000000000000000010001110110111;
ROM[1794] <= 32'b11000101000000111000001110010011;
ROM[1795] <= 32'b00000000111000111000001110110011;
ROM[1796] <= 32'b00000000011100010010000000100011;
ROM[1797] <= 32'b00000000010000010000000100010011;
ROM[1798] <= 32'b00000000001100010010000000100011;
ROM[1799] <= 32'b00000000010000010000000100010011;
ROM[1800] <= 32'b00000000010000010010000000100011;
ROM[1801] <= 32'b00000000010000010000000100010011;
ROM[1802] <= 32'b00000000010100010010000000100011;
ROM[1803] <= 32'b00000000010000010000000100010011;
ROM[1804] <= 32'b00000000011000010010000000100011;
ROM[1805] <= 32'b00000000010000010000000100010011;
ROM[1806] <= 32'b00000001010000000000001110010011;
ROM[1807] <= 32'b00000000100000111000001110010011;
ROM[1808] <= 32'b01000000011100010000001110110011;
ROM[1809] <= 32'b00000000011100000000001000110011;
ROM[1810] <= 32'b00000000001000000000000110110011;
ROM[1811] <= 32'b01110110000100100111000011101111;
ROM[1812] <= 32'b00000111010100000000001110010011;
ROM[1813] <= 32'b00000000011100010010000000100011;
ROM[1814] <= 32'b00000000010000010000000100010011;
ROM[1815] <= 32'b00000000000000000010001110110111;
ROM[1816] <= 32'b11001010100000111000001110010011;
ROM[1817] <= 32'b00000000111000111000001110110011;
ROM[1818] <= 32'b00000000011100010010000000100011;
ROM[1819] <= 32'b00000000010000010000000100010011;
ROM[1820] <= 32'b00000000001100010010000000100011;
ROM[1821] <= 32'b00000000010000010000000100010011;
ROM[1822] <= 32'b00000000010000010010000000100011;
ROM[1823] <= 32'b00000000010000010000000100010011;
ROM[1824] <= 32'b00000000010100010010000000100011;
ROM[1825] <= 32'b00000000010000010000000100010011;
ROM[1826] <= 32'b00000000011000010010000000100011;
ROM[1827] <= 32'b00000000010000010000000100010011;
ROM[1828] <= 32'b00000001010000000000001110010011;
ROM[1829] <= 32'b00000000100000111000001110010011;
ROM[1830] <= 32'b01000000011100010000001110110011;
ROM[1831] <= 32'b00000000011100000000001000110011;
ROM[1832] <= 32'b00000000001000000000000110110011;
ROM[1833] <= 32'b01110000100100100111000011101111;
ROM[1834] <= 32'b00000110110100000000001110010011;
ROM[1835] <= 32'b00000000011100010010000000100011;
ROM[1836] <= 32'b00000000010000010000000100010011;
ROM[1837] <= 32'b00000000000000000010001110110111;
ROM[1838] <= 32'b11010000000000111000001110010011;
ROM[1839] <= 32'b00000000111000111000001110110011;
ROM[1840] <= 32'b00000000011100010010000000100011;
ROM[1841] <= 32'b00000000010000010000000100010011;
ROM[1842] <= 32'b00000000001100010010000000100011;
ROM[1843] <= 32'b00000000010000010000000100010011;
ROM[1844] <= 32'b00000000010000010010000000100011;
ROM[1845] <= 32'b00000000010000010000000100010011;
ROM[1846] <= 32'b00000000010100010010000000100011;
ROM[1847] <= 32'b00000000010000010000000100010011;
ROM[1848] <= 32'b00000000011000010010000000100011;
ROM[1849] <= 32'b00000000010000010000000100010011;
ROM[1850] <= 32'b00000001010000000000001110010011;
ROM[1851] <= 32'b00000000100000111000001110010011;
ROM[1852] <= 32'b01000000011100010000001110110011;
ROM[1853] <= 32'b00000000011100000000001000110011;
ROM[1854] <= 32'b00000000001000000000000110110011;
ROM[1855] <= 32'b01101011000100100111000011101111;
ROM[1856] <= 32'b00000110001000000000001110010011;
ROM[1857] <= 32'b00000000011100010010000000100011;
ROM[1858] <= 32'b00000000010000010000000100010011;
ROM[1859] <= 32'b00000000000000000010001110110111;
ROM[1860] <= 32'b11010101100000111000001110010011;
ROM[1861] <= 32'b00000000111000111000001110110011;
ROM[1862] <= 32'b00000000011100010010000000100011;
ROM[1863] <= 32'b00000000010000010000000100010011;
ROM[1864] <= 32'b00000000001100010010000000100011;
ROM[1865] <= 32'b00000000010000010000000100010011;
ROM[1866] <= 32'b00000000010000010010000000100011;
ROM[1867] <= 32'b00000000010000010000000100010011;
ROM[1868] <= 32'b00000000010100010010000000100011;
ROM[1869] <= 32'b00000000010000010000000100010011;
ROM[1870] <= 32'b00000000011000010010000000100011;
ROM[1871] <= 32'b00000000010000010000000100010011;
ROM[1872] <= 32'b00000001010000000000001110010011;
ROM[1873] <= 32'b00000000100000111000001110010011;
ROM[1874] <= 32'b01000000011100010000001110110011;
ROM[1875] <= 32'b00000000011100000000001000110011;
ROM[1876] <= 32'b00000000001000000000000110110011;
ROM[1877] <= 32'b01100101100100100111000011101111;
ROM[1878] <= 32'b00000110010100000000001110010011;
ROM[1879] <= 32'b00000000011100010010000000100011;
ROM[1880] <= 32'b00000000010000010000000100010011;
ROM[1881] <= 32'b00000000000000000010001110110111;
ROM[1882] <= 32'b11011011000000111000001110010011;
ROM[1883] <= 32'b00000000111000111000001110110011;
ROM[1884] <= 32'b00000000011100010010000000100011;
ROM[1885] <= 32'b00000000010000010000000100010011;
ROM[1886] <= 32'b00000000001100010010000000100011;
ROM[1887] <= 32'b00000000010000010000000100010011;
ROM[1888] <= 32'b00000000010000010010000000100011;
ROM[1889] <= 32'b00000000010000010000000100010011;
ROM[1890] <= 32'b00000000010100010010000000100011;
ROM[1891] <= 32'b00000000010000010000000100010011;
ROM[1892] <= 32'b00000000011000010010000000100011;
ROM[1893] <= 32'b00000000010000010000000100010011;
ROM[1894] <= 32'b00000001010000000000001110010011;
ROM[1895] <= 32'b00000000100000111000001110010011;
ROM[1896] <= 32'b01000000011100010000001110110011;
ROM[1897] <= 32'b00000000011100000000001000110011;
ROM[1898] <= 32'b00000000001000000000000110110011;
ROM[1899] <= 32'b01100000000100100111000011101111;
ROM[1900] <= 32'b00000111001000000000001110010011;
ROM[1901] <= 32'b00000000011100010010000000100011;
ROM[1902] <= 32'b00000000010000010000000100010011;
ROM[1903] <= 32'b00000000000000000010001110110111;
ROM[1904] <= 32'b11100000100000111000001110010011;
ROM[1905] <= 32'b00000000111000111000001110110011;
ROM[1906] <= 32'b00000000011100010010000000100011;
ROM[1907] <= 32'b00000000010000010000000100010011;
ROM[1908] <= 32'b00000000001100010010000000100011;
ROM[1909] <= 32'b00000000010000010000000100010011;
ROM[1910] <= 32'b00000000010000010010000000100011;
ROM[1911] <= 32'b00000000010000010000000100010011;
ROM[1912] <= 32'b00000000010100010010000000100011;
ROM[1913] <= 32'b00000000010000010000000100010011;
ROM[1914] <= 32'b00000000011000010010000000100011;
ROM[1915] <= 32'b00000000010000010000000100010011;
ROM[1916] <= 32'b00000001010000000000001110010011;
ROM[1917] <= 32'b00000000100000111000001110010011;
ROM[1918] <= 32'b01000000011100010000001110110011;
ROM[1919] <= 32'b00000000011100000000001000110011;
ROM[1920] <= 32'b00000000001000000000000110110011;
ROM[1921] <= 32'b01011010100100100111000011101111;
ROM[1922] <= 32'b00000111001100000000001110010011;
ROM[1923] <= 32'b00000000011100010010000000100011;
ROM[1924] <= 32'b00000000010000010000000100010011;
ROM[1925] <= 32'b00000000000000000010001110110111;
ROM[1926] <= 32'b11100110000000111000001110010011;
ROM[1927] <= 32'b00000000111000111000001110110011;
ROM[1928] <= 32'b00000000011100010010000000100011;
ROM[1929] <= 32'b00000000010000010000000100010011;
ROM[1930] <= 32'b00000000001100010010000000100011;
ROM[1931] <= 32'b00000000010000010000000100010011;
ROM[1932] <= 32'b00000000010000010010000000100011;
ROM[1933] <= 32'b00000000010000010000000100010011;
ROM[1934] <= 32'b00000000010100010010000000100011;
ROM[1935] <= 32'b00000000010000010000000100010011;
ROM[1936] <= 32'b00000000011000010010000000100011;
ROM[1937] <= 32'b00000000010000010000000100010011;
ROM[1938] <= 32'b00000001010000000000001110010011;
ROM[1939] <= 32'b00000000100000111000001110010011;
ROM[1940] <= 32'b01000000011100010000001110110011;
ROM[1941] <= 32'b00000000011100000000001000110011;
ROM[1942] <= 32'b00000000001000000000000110110011;
ROM[1943] <= 32'b01010101000100100111000011101111;
ROM[1944] <= 32'b00000010000000000000001110010011;
ROM[1945] <= 32'b00000000011100010010000000100011;
ROM[1946] <= 32'b00000000010000010000000100010011;
ROM[1947] <= 32'b00000000000000000010001110110111;
ROM[1948] <= 32'b11101011100000111000001110010011;
ROM[1949] <= 32'b00000000111000111000001110110011;
ROM[1950] <= 32'b00000000011100010010000000100011;
ROM[1951] <= 32'b00000000010000010000000100010011;
ROM[1952] <= 32'b00000000001100010010000000100011;
ROM[1953] <= 32'b00000000010000010000000100010011;
ROM[1954] <= 32'b00000000010000010010000000100011;
ROM[1955] <= 32'b00000000010000010000000100010011;
ROM[1956] <= 32'b00000000010100010010000000100011;
ROM[1957] <= 32'b00000000010000010000000100010011;
ROM[1958] <= 32'b00000000011000010010000000100011;
ROM[1959] <= 32'b00000000010000010000000100010011;
ROM[1960] <= 32'b00000001010000000000001110010011;
ROM[1961] <= 32'b00000000100000111000001110010011;
ROM[1962] <= 32'b01000000011100010000001110110011;
ROM[1963] <= 32'b00000000011100000000001000110011;
ROM[1964] <= 32'b00000000001000000000000110110011;
ROM[1965] <= 32'b01001111100100100111000011101111;
ROM[1966] <= 32'b00000110000100000000001110010011;
ROM[1967] <= 32'b00000000011100010010000000100011;
ROM[1968] <= 32'b00000000010000010000000100010011;
ROM[1969] <= 32'b00000000000000000010001110110111;
ROM[1970] <= 32'b11110001000000111000001110010011;
ROM[1971] <= 32'b00000000111000111000001110110011;
ROM[1972] <= 32'b00000000011100010010000000100011;
ROM[1973] <= 32'b00000000010000010000000100010011;
ROM[1974] <= 32'b00000000001100010010000000100011;
ROM[1975] <= 32'b00000000010000010000000100010011;
ROM[1976] <= 32'b00000000010000010010000000100011;
ROM[1977] <= 32'b00000000010000010000000100010011;
ROM[1978] <= 32'b00000000010100010010000000100011;
ROM[1979] <= 32'b00000000010000010000000100010011;
ROM[1980] <= 32'b00000000011000010010000000100011;
ROM[1981] <= 32'b00000000010000010000000100010011;
ROM[1982] <= 32'b00000001010000000000001110010011;
ROM[1983] <= 32'b00000000100000111000001110010011;
ROM[1984] <= 32'b01000000011100010000001110110011;
ROM[1985] <= 32'b00000000011100000000001000110011;
ROM[1986] <= 32'b00000000001000000000000110110011;
ROM[1987] <= 32'b01001010000100100111000011101111;
ROM[1988] <= 32'b00000111001000000000001110010011;
ROM[1989] <= 32'b00000000011100010010000000100011;
ROM[1990] <= 32'b00000000010000010000000100010011;
ROM[1991] <= 32'b00000000000000000010001110110111;
ROM[1992] <= 32'b11110110100000111000001110010011;
ROM[1993] <= 32'b00000000111000111000001110110011;
ROM[1994] <= 32'b00000000011100010010000000100011;
ROM[1995] <= 32'b00000000010000010000000100010011;
ROM[1996] <= 32'b00000000001100010010000000100011;
ROM[1997] <= 32'b00000000010000010000000100010011;
ROM[1998] <= 32'b00000000010000010010000000100011;
ROM[1999] <= 32'b00000000010000010000000100010011;
ROM[2000] <= 32'b00000000010100010010000000100011;
ROM[2001] <= 32'b00000000010000010000000100010011;
ROM[2002] <= 32'b00000000011000010010000000100011;
ROM[2003] <= 32'b00000000010000010000000100010011;
ROM[2004] <= 32'b00000001010000000000001110010011;
ROM[2005] <= 32'b00000000100000111000001110010011;
ROM[2006] <= 32'b01000000011100010000001110110011;
ROM[2007] <= 32'b00000000011100000000001000110011;
ROM[2008] <= 32'b00000000001000000000000110110011;
ROM[2009] <= 32'b01000100100100100111000011101111;
ROM[2010] <= 32'b00000110010100000000001110010011;
ROM[2011] <= 32'b00000000011100010010000000100011;
ROM[2012] <= 32'b00000000010000010000000100010011;
ROM[2013] <= 32'b00000000000000000010001110110111;
ROM[2014] <= 32'b11111100000000111000001110010011;
ROM[2015] <= 32'b00000000111000111000001110110011;
ROM[2016] <= 32'b00000000011100010010000000100011;
ROM[2017] <= 32'b00000000010000010000000100010011;
ROM[2018] <= 32'b00000000001100010010000000100011;
ROM[2019] <= 32'b00000000010000010000000100010011;
ROM[2020] <= 32'b00000000010000010010000000100011;
ROM[2021] <= 32'b00000000010000010000000100010011;
ROM[2022] <= 32'b00000000010100010010000000100011;
ROM[2023] <= 32'b00000000010000010000000100010011;
ROM[2024] <= 32'b00000000011000010010000000100011;
ROM[2025] <= 32'b00000000010000010000000100010011;
ROM[2026] <= 32'b00000001010000000000001110010011;
ROM[2027] <= 32'b00000000100000111000001110010011;
ROM[2028] <= 32'b01000000011100010000001110110011;
ROM[2029] <= 32'b00000000011100000000001000110011;
ROM[2030] <= 32'b00000000001000000000000110110011;
ROM[2031] <= 32'b00111111000100100111000011101111;
ROM[2032] <= 32'b00000011101000000000001110010011;
ROM[2033] <= 32'b00000000011100010010000000100011;
ROM[2034] <= 32'b00000000010000010000000100010011;
ROM[2035] <= 32'b00000000000000000010001110110111;
ROM[2036] <= 32'b00000001100000111000001110010011;
ROM[2037] <= 32'b00000000111000111000001110110011;
ROM[2038] <= 32'b00000000011100010010000000100011;
ROM[2039] <= 32'b00000000010000010000000100010011;
ROM[2040] <= 32'b00000000001100010010000000100011;
ROM[2041] <= 32'b00000000010000010000000100010011;
ROM[2042] <= 32'b00000000010000010010000000100011;
ROM[2043] <= 32'b00000000010000010000000100010011;
ROM[2044] <= 32'b00000000010100010010000000100011;
ROM[2045] <= 32'b00000000010000010000000100010011;
ROM[2046] <= 32'b00000000011000010010000000100011;
ROM[2047] <= 32'b00000000010000010000000100010011;
ROM[2048] <= 32'b00000001010000000000001110010011;
ROM[2049] <= 32'b00000000100000111000001110010011;
ROM[2050] <= 32'b01000000011100010000001110110011;
ROM[2051] <= 32'b00000000011100000000001000110011;
ROM[2052] <= 32'b00000000001000000000000110110011;
ROM[2053] <= 32'b00111001100100100111000011101111;
ROM[2054] <= 32'b00000010000000000000001110010011;
ROM[2055] <= 32'b00000000011100010010000000100011;
ROM[2056] <= 32'b00000000010000010000000100010011;
ROM[2057] <= 32'b00000000000000000010001110110111;
ROM[2058] <= 32'b00000111000000111000001110010011;
ROM[2059] <= 32'b00000000111000111000001110110011;
ROM[2060] <= 32'b00000000011100010010000000100011;
ROM[2061] <= 32'b00000000010000010000000100010011;
ROM[2062] <= 32'b00000000001100010010000000100011;
ROM[2063] <= 32'b00000000010000010000000100010011;
ROM[2064] <= 32'b00000000010000010010000000100011;
ROM[2065] <= 32'b00000000010000010000000100010011;
ROM[2066] <= 32'b00000000010100010010000000100011;
ROM[2067] <= 32'b00000000010000010000000100010011;
ROM[2068] <= 32'b00000000011000010010000000100011;
ROM[2069] <= 32'b00000000010000010000000100010011;
ROM[2070] <= 32'b00000001010000000000001110010011;
ROM[2071] <= 32'b00000000100000111000001110010011;
ROM[2072] <= 32'b01000000011100010000001110110011;
ROM[2073] <= 32'b00000000011100000000001000110011;
ROM[2074] <= 32'b00000000001000000000000110110011;
ROM[2075] <= 32'b00110100000100100111000011101111;
ROM[2076] <= 32'b00000000000000000010001110110111;
ROM[2077] <= 32'b00001011110000111000001110010011;
ROM[2078] <= 32'b00000000111000111000001110110011;
ROM[2079] <= 32'b00000000011100010010000000100011;
ROM[2080] <= 32'b00000000010000010000000100010011;
ROM[2081] <= 32'b00000000001100010010000000100011;
ROM[2082] <= 32'b00000000010000010000000100010011;
ROM[2083] <= 32'b00000000010000010010000000100011;
ROM[2084] <= 32'b00000000010000010000000100010011;
ROM[2085] <= 32'b00000000010100010010000000100011;
ROM[2086] <= 32'b00000000010000010000000100010011;
ROM[2087] <= 32'b00000000011000010010000000100011;
ROM[2088] <= 32'b00000000010000010000000100010011;
ROM[2089] <= 32'b00000001010000000000001110010011;
ROM[2090] <= 32'b00000000010000111000001110010011;
ROM[2091] <= 32'b01000000011100010000001110110011;
ROM[2092] <= 32'b00000000011100000000001000110011;
ROM[2093] <= 32'b00000000001000000000000110110011;
ROM[2094] <= 32'b01101011000100010100000011101111;
ROM[2095] <= 32'b11111111110000010000000100010011;
ROM[2096] <= 32'b00000000000000010010001110000011;
ROM[2097] <= 32'b00000000011101100010000000100011;
ROM[2098] <= 32'b00000000010000011010001110000011;
ROM[2099] <= 32'b00000000011100010010000000100011;
ROM[2100] <= 32'b00000000010000010000000100010011;
ROM[2101] <= 32'b00000000000000000010001110110111;
ROM[2102] <= 32'b00010010000000111000001110010011;
ROM[2103] <= 32'b00000000111000111000001110110011;
ROM[2104] <= 32'b00000000011100010010000000100011;
ROM[2105] <= 32'b00000000010000010000000100010011;
ROM[2106] <= 32'b00000000001100010010000000100011;
ROM[2107] <= 32'b00000000010000010000000100010011;
ROM[2108] <= 32'b00000000010000010010000000100011;
ROM[2109] <= 32'b00000000010000010000000100010011;
ROM[2110] <= 32'b00000000010100010010000000100011;
ROM[2111] <= 32'b00000000010000010000000100010011;
ROM[2112] <= 32'b00000000011000010010000000100011;
ROM[2113] <= 32'b00000000010000010000000100010011;
ROM[2114] <= 32'b00000001010000000000001110010011;
ROM[2115] <= 32'b00000000010000111000001110010011;
ROM[2116] <= 32'b01000000011100010000001110110011;
ROM[2117] <= 32'b00000000011100000000001000110011;
ROM[2118] <= 32'b00000000001000000000000110110011;
ROM[2119] <= 32'b00000110010000010101000011101111;
ROM[2120] <= 32'b11111111110000010000000100010011;
ROM[2121] <= 32'b00000000000000010010001110000011;
ROM[2122] <= 32'b00000000011101100010000000100011;
ROM[2123] <= 32'b00000000000000011010001110000011;
ROM[2124] <= 32'b00000000011100010010000000100011;
ROM[2125] <= 32'b00000000010000010000000100010011;
ROM[2126] <= 32'b00000000000100000000001110010011;
ROM[2127] <= 32'b00000000011100010010000000100011;
ROM[2128] <= 32'b00000000010000010000000100010011;
ROM[2129] <= 32'b11111111110000010000000100010011;
ROM[2130] <= 32'b00000000000000010010001110000011;
ROM[2131] <= 32'b11111111110000010000000100010011;
ROM[2132] <= 32'b00000000000000010010010000000011;
ROM[2133] <= 32'b00000000100000111010001110110011;
ROM[2134] <= 32'b00000000011100010010000000100011;
ROM[2135] <= 32'b00000000010000010000000100010011;
ROM[2136] <= 32'b11111111110000010000000100010011;
ROM[2137] <= 32'b00000000000000010010001110000011;
ROM[2138] <= 32'b00000000000000111000101001100011;
ROM[2139] <= 32'b00000000000000000010001110110111;
ROM[2140] <= 32'b00011000000000111000001110010011;
ROM[2141] <= 32'b00000000111000111000001110110011;
ROM[2142] <= 32'b00000000000000111000000011100111;
ROM[2143] <= 32'b00011100100000000000000011101111;
ROM[2144] <= 32'b00000000001000000000001110010011;
ROM[2145] <= 32'b00000000011100010010000000100011;
ROM[2146] <= 32'b00000000010000010000000100010011;
ROM[2147] <= 32'b00000000000000000010001110110111;
ROM[2148] <= 32'b00011101100000111000001110010011;
ROM[2149] <= 32'b00000000111000111000001110110011;
ROM[2150] <= 32'b00000000011100010010000000100011;
ROM[2151] <= 32'b00000000010000010000000100010011;
ROM[2152] <= 32'b00000000001100010010000000100011;
ROM[2153] <= 32'b00000000010000010000000100010011;
ROM[2154] <= 32'b00000000010000010010000000100011;
ROM[2155] <= 32'b00000000010000010000000100010011;
ROM[2156] <= 32'b00000000010100010010000000100011;
ROM[2157] <= 32'b00000000010000010000000100010011;
ROM[2158] <= 32'b00000000011000010010000000100011;
ROM[2159] <= 32'b00000000010000010000000100010011;
ROM[2160] <= 32'b00000001010000000000001110010011;
ROM[2161] <= 32'b00000000010000111000001110010011;
ROM[2162] <= 32'b01000000011100010000001110110011;
ROM[2163] <= 32'b00000000011100000000001000110011;
ROM[2164] <= 32'b00000000001000000000000110110011;
ROM[2165] <= 32'b01010110100000100111000011101111;
ROM[2166] <= 32'b00000010110000000000001110010011;
ROM[2167] <= 32'b00000000011100010010000000100011;
ROM[2168] <= 32'b00000000010000010000000100010011;
ROM[2169] <= 32'b00000000000000000010001110110111;
ROM[2170] <= 32'b00100011000000111000001110010011;
ROM[2171] <= 32'b00000000111000111000001110110011;
ROM[2172] <= 32'b00000000011100010010000000100011;
ROM[2173] <= 32'b00000000010000010000000100010011;
ROM[2174] <= 32'b00000000001100010010000000100011;
ROM[2175] <= 32'b00000000010000010000000100010011;
ROM[2176] <= 32'b00000000010000010010000000100011;
ROM[2177] <= 32'b00000000010000010000000100010011;
ROM[2178] <= 32'b00000000010100010010000000100011;
ROM[2179] <= 32'b00000000010000010000000100010011;
ROM[2180] <= 32'b00000000011000010010000000100011;
ROM[2181] <= 32'b00000000010000010000000100010011;
ROM[2182] <= 32'b00000001010000000000001110010011;
ROM[2183] <= 32'b00000000100000111000001110010011;
ROM[2184] <= 32'b01000000011100010000001110110011;
ROM[2185] <= 32'b00000000011100000000001000110011;
ROM[2186] <= 32'b00000000001000000000000110110011;
ROM[2187] <= 32'b00011000000100100111000011101111;
ROM[2188] <= 32'b00000010000000000000001110010011;
ROM[2189] <= 32'b00000000011100010010000000100011;
ROM[2190] <= 32'b00000000010000010000000100010011;
ROM[2191] <= 32'b00000000000000000010001110110111;
ROM[2192] <= 32'b00101000100000111000001110010011;
ROM[2193] <= 32'b00000000111000111000001110110011;
ROM[2194] <= 32'b00000000011100010010000000100011;
ROM[2195] <= 32'b00000000010000010000000100010011;
ROM[2196] <= 32'b00000000001100010010000000100011;
ROM[2197] <= 32'b00000000010000010000000100010011;
ROM[2198] <= 32'b00000000010000010010000000100011;
ROM[2199] <= 32'b00000000010000010000000100010011;
ROM[2200] <= 32'b00000000010100010010000000100011;
ROM[2201] <= 32'b00000000010000010000000100010011;
ROM[2202] <= 32'b00000000011000010010000000100011;
ROM[2203] <= 32'b00000000010000010000000100010011;
ROM[2204] <= 32'b00000001010000000000001110010011;
ROM[2205] <= 32'b00000000100000111000001110010011;
ROM[2206] <= 32'b01000000011100010000001110110011;
ROM[2207] <= 32'b00000000011100000000001000110011;
ROM[2208] <= 32'b00000000001000000000000110110011;
ROM[2209] <= 32'b00010010100100100111000011101111;
ROM[2210] <= 32'b00000000000000000010001110110111;
ROM[2211] <= 32'b00101101010000111000001110010011;
ROM[2212] <= 32'b00000000111000111000001110110011;
ROM[2213] <= 32'b00000000011100010010000000100011;
ROM[2214] <= 32'b00000000010000010000000100010011;
ROM[2215] <= 32'b00000000001100010010000000100011;
ROM[2216] <= 32'b00000000010000010000000100010011;
ROM[2217] <= 32'b00000000010000010010000000100011;
ROM[2218] <= 32'b00000000010000010000000100010011;
ROM[2219] <= 32'b00000000010100010010000000100011;
ROM[2220] <= 32'b00000000010000010000000100010011;
ROM[2221] <= 32'b00000000011000010010000000100011;
ROM[2222] <= 32'b00000000010000010000000100010011;
ROM[2223] <= 32'b00000001010000000000001110010011;
ROM[2224] <= 32'b00000000010000111000001110010011;
ROM[2225] <= 32'b01000000011100010000001110110011;
ROM[2226] <= 32'b00000000011100000000001000110011;
ROM[2227] <= 32'b00000000001000000000000110110011;
ROM[2228] <= 32'b01001001100100010100000011101111;
ROM[2229] <= 32'b11111111110000010000000100010011;
ROM[2230] <= 32'b00000000000000010010001110000011;
ROM[2231] <= 32'b00000000011101100010000000100011;
ROM[2232] <= 32'b00000000100000011010001110000011;
ROM[2233] <= 32'b00000000011100010010000000100011;
ROM[2234] <= 32'b00000000010000010000000100010011;
ROM[2235] <= 32'b00000000000000000010001110110111;
ROM[2236] <= 32'b00110011100000111000001110010011;
ROM[2237] <= 32'b00000000111000111000001110110011;
ROM[2238] <= 32'b00000000011100010010000000100011;
ROM[2239] <= 32'b00000000010000010000000100010011;
ROM[2240] <= 32'b00000000001100010010000000100011;
ROM[2241] <= 32'b00000000010000010000000100010011;
ROM[2242] <= 32'b00000000010000010010000000100011;
ROM[2243] <= 32'b00000000010000010000000100010011;
ROM[2244] <= 32'b00000000010100010010000000100011;
ROM[2245] <= 32'b00000000010000010000000100010011;
ROM[2246] <= 32'b00000000011000010010000000100011;
ROM[2247] <= 32'b00000000010000010000000100010011;
ROM[2248] <= 32'b00000001010000000000001110010011;
ROM[2249] <= 32'b00000000010000111000001110010011;
ROM[2250] <= 32'b01000000011100010000001110110011;
ROM[2251] <= 32'b00000000011100000000001000110011;
ROM[2252] <= 32'b00000000001000000000000110110011;
ROM[2253] <= 32'b01100100110100010100000011101111;
ROM[2254] <= 32'b11111111110000010000000100010011;
ROM[2255] <= 32'b00000000000000010010001110000011;
ROM[2256] <= 32'b00000000011101100010000000100011;
ROM[2257] <= 32'b00000000001000000000001110010011;
ROM[2258] <= 32'b00000000011100010010000000100011;
ROM[2259] <= 32'b00000000010000010000000100010011;
ROM[2260] <= 32'b11111111110000010000000100010011;
ROM[2261] <= 32'b00000000000000010010001110000011;
ROM[2262] <= 32'b00000000011100011010100000100011;
ROM[2263] <= 32'b00000001000000011010001110000011;
ROM[2264] <= 32'b00000000011100010010000000100011;
ROM[2265] <= 32'b00000000010000010000000100010011;
ROM[2266] <= 32'b00000000000000011010001110000011;
ROM[2267] <= 32'b00000000011100010010000000100011;
ROM[2268] <= 32'b00000000010000010000000100010011;
ROM[2269] <= 32'b11111111110000010000000100010011;
ROM[2270] <= 32'b00000000000000010010001110000011;
ROM[2271] <= 32'b11111111110000010000000100010011;
ROM[2272] <= 32'b00000000000000010010010000000011;
ROM[2273] <= 32'b00000000011101000010001110110011;
ROM[2274] <= 32'b00000000011100010010000000100011;
ROM[2275] <= 32'b00000000010000010000000100010011;
ROM[2276] <= 32'b11111111110000010000000100010011;
ROM[2277] <= 32'b00000000000000010010001110000011;
ROM[2278] <= 32'b01000000011100000000001110110011;
ROM[2279] <= 32'b00000000000100111000001110010011;
ROM[2280] <= 32'b00000000011100010010000000100011;
ROM[2281] <= 32'b00000000010000010000000100010011;
ROM[2282] <= 32'b11111111110000010000000100010011;
ROM[2283] <= 32'b00000000000000010010001110000011;
ROM[2284] <= 32'b00000000000000111000101001100011;
ROM[2285] <= 32'b00000000000000000010001110110111;
ROM[2286] <= 32'b01100011110000111000001110010011;
ROM[2287] <= 32'b00000000111000111000001110110011;
ROM[2288] <= 32'b00000000000000111000000011100111;
ROM[2289] <= 32'b00000000010000011010001110000011;
ROM[2290] <= 32'b00000000011100010010000000100011;
ROM[2291] <= 32'b00000000010000010000000100010011;
ROM[2292] <= 32'b00000000100000011010001110000011;
ROM[2293] <= 32'b00000000011100010010000000100011;
ROM[2294] <= 32'b00000000010000010000000100010011;
ROM[2295] <= 32'b11111111110000010000000100010011;
ROM[2296] <= 32'b00000000000000010010001110000011;
ROM[2297] <= 32'b11111111110000010000000100010011;
ROM[2298] <= 32'b00000000000000010010010000000011;
ROM[2299] <= 32'b00000000011101000000001110110011;
ROM[2300] <= 32'b00000000011100010010000000100011;
ROM[2301] <= 32'b00000000010000010000000100010011;
ROM[2302] <= 32'b11111111110000010000000100010011;
ROM[2303] <= 32'b00000000000000010010001110000011;
ROM[2304] <= 32'b00000000011100011010011000100011;
ROM[2305] <= 32'b00000000001000000000001110010011;
ROM[2306] <= 32'b00000000011100010010000000100011;
ROM[2307] <= 32'b00000000010000010000000100010011;
ROM[2308] <= 32'b00000000000000000010001110110111;
ROM[2309] <= 32'b01000101110000111000001110010011;
ROM[2310] <= 32'b00000000111000111000001110110011;
ROM[2311] <= 32'b00000000011100010010000000100011;
ROM[2312] <= 32'b00000000010000010000000100010011;
ROM[2313] <= 32'b00000000001100010010000000100011;
ROM[2314] <= 32'b00000000010000010000000100010011;
ROM[2315] <= 32'b00000000010000010010000000100011;
ROM[2316] <= 32'b00000000010000010000000100010011;
ROM[2317] <= 32'b00000000010100010010000000100011;
ROM[2318] <= 32'b00000000010000010000000100010011;
ROM[2319] <= 32'b00000000011000010010000000100011;
ROM[2320] <= 32'b00000000010000010000000100010011;
ROM[2321] <= 32'b00000001010000000000001110010011;
ROM[2322] <= 32'b00000000010000111000001110010011;
ROM[2323] <= 32'b01000000011100010000001110110011;
ROM[2324] <= 32'b00000000011100000000001000110011;
ROM[2325] <= 32'b00000000001000000000000110110011;
ROM[2326] <= 32'b00101110010000100111000011101111;
ROM[2327] <= 32'b00000010110000000000001110010011;
ROM[2328] <= 32'b00000000011100010010000000100011;
ROM[2329] <= 32'b00000000010000010000000100010011;
ROM[2330] <= 32'b00000000000000000010001110110111;
ROM[2331] <= 32'b01001011010000111000001110010011;
ROM[2332] <= 32'b00000000111000111000001110110011;
ROM[2333] <= 32'b00000000011100010010000000100011;
ROM[2334] <= 32'b00000000010000010000000100010011;
ROM[2335] <= 32'b00000000001100010010000000100011;
ROM[2336] <= 32'b00000000010000010000000100010011;
ROM[2337] <= 32'b00000000010000010010000000100011;
ROM[2338] <= 32'b00000000010000010000000100010011;
ROM[2339] <= 32'b00000000010100010010000000100011;
ROM[2340] <= 32'b00000000010000010000000100010011;
ROM[2341] <= 32'b00000000011000010010000000100011;
ROM[2342] <= 32'b00000000010000010000000100010011;
ROM[2343] <= 32'b00000001010000000000001110010011;
ROM[2344] <= 32'b00000000100000111000001110010011;
ROM[2345] <= 32'b01000000011100010000001110110011;
ROM[2346] <= 32'b00000000011100000000001000110011;
ROM[2347] <= 32'b00000000001000000000000110110011;
ROM[2348] <= 32'b01101111110000100111000011101111;
ROM[2349] <= 32'b00000010000000000000001110010011;
ROM[2350] <= 32'b00000000011100010010000000100011;
ROM[2351] <= 32'b00000000010000010000000100010011;
ROM[2352] <= 32'b00000000000000000010001110110111;
ROM[2353] <= 32'b01010000110000111000001110010011;
ROM[2354] <= 32'b00000000111000111000001110110011;
ROM[2355] <= 32'b00000000011100010010000000100011;
ROM[2356] <= 32'b00000000010000010000000100010011;
ROM[2357] <= 32'b00000000001100010010000000100011;
ROM[2358] <= 32'b00000000010000010000000100010011;
ROM[2359] <= 32'b00000000010000010010000000100011;
ROM[2360] <= 32'b00000000010000010000000100010011;
ROM[2361] <= 32'b00000000010100010010000000100011;
ROM[2362] <= 32'b00000000010000010000000100010011;
ROM[2363] <= 32'b00000000011000010010000000100011;
ROM[2364] <= 32'b00000000010000010000000100010011;
ROM[2365] <= 32'b00000001010000000000001110010011;
ROM[2366] <= 32'b00000000100000111000001110010011;
ROM[2367] <= 32'b01000000011100010000001110110011;
ROM[2368] <= 32'b00000000011100000000001000110011;
ROM[2369] <= 32'b00000000001000000000000110110011;
ROM[2370] <= 32'b01101010010000100111000011101111;
ROM[2371] <= 32'b00000000000000000010001110110111;
ROM[2372] <= 32'b01010101100000111000001110010011;
ROM[2373] <= 32'b00000000111000111000001110110011;
ROM[2374] <= 32'b00000000011100010010000000100011;
ROM[2375] <= 32'b00000000010000010000000100010011;
ROM[2376] <= 32'b00000000001100010010000000100011;
ROM[2377] <= 32'b00000000010000010000000100010011;
ROM[2378] <= 32'b00000000010000010010000000100011;
ROM[2379] <= 32'b00000000010000010000000100010011;
ROM[2380] <= 32'b00000000010100010010000000100011;
ROM[2381] <= 32'b00000000010000010000000100010011;
ROM[2382] <= 32'b00000000011000010010000000100011;
ROM[2383] <= 32'b00000000010000010000000100010011;
ROM[2384] <= 32'b00000001010000000000001110010011;
ROM[2385] <= 32'b00000000010000111000001110010011;
ROM[2386] <= 32'b01000000011100010000001110110011;
ROM[2387] <= 32'b00000000011100000000001000110011;
ROM[2388] <= 32'b00000000001000000000000110110011;
ROM[2389] <= 32'b00100001010100010100000011101111;
ROM[2390] <= 32'b11111111110000010000000100010011;
ROM[2391] <= 32'b00000000000000010010001110000011;
ROM[2392] <= 32'b00000000011101100010000000100011;
ROM[2393] <= 32'b00000000110000011010001110000011;
ROM[2394] <= 32'b00000000011100010010000000100011;
ROM[2395] <= 32'b00000000010000010000000100010011;
ROM[2396] <= 32'b00000000000000000010001110110111;
ROM[2397] <= 32'b01011011110000111000001110010011;
ROM[2398] <= 32'b00000000111000111000001110110011;
ROM[2399] <= 32'b00000000011100010010000000100011;
ROM[2400] <= 32'b00000000010000010000000100010011;
ROM[2401] <= 32'b00000000001100010010000000100011;
ROM[2402] <= 32'b00000000010000010000000100010011;
ROM[2403] <= 32'b00000000010000010010000000100011;
ROM[2404] <= 32'b00000000010000010000000100010011;
ROM[2405] <= 32'b00000000010100010010000000100011;
ROM[2406] <= 32'b00000000010000010000000100010011;
ROM[2407] <= 32'b00000000011000010010000000100011;
ROM[2408] <= 32'b00000000010000010000000100010011;
ROM[2409] <= 32'b00000001010000000000001110010011;
ROM[2410] <= 32'b00000000010000111000001110010011;
ROM[2411] <= 32'b01000000011100010000001110110011;
ROM[2412] <= 32'b00000000011100000000001000110011;
ROM[2413] <= 32'b00000000001000000000000110110011;
ROM[2414] <= 32'b00111100100100010100000011101111;
ROM[2415] <= 32'b11111111110000010000000100010011;
ROM[2416] <= 32'b00000000000000010010001110000011;
ROM[2417] <= 32'b00000000011101100010000000100011;
ROM[2418] <= 32'b00000000100000011010001110000011;
ROM[2419] <= 32'b00000000011100010010000000100011;
ROM[2420] <= 32'b00000000010000010000000100010011;
ROM[2421] <= 32'b11111111110000010000000100010011;
ROM[2422] <= 32'b00000000000000010010001110000011;
ROM[2423] <= 32'b00000000011100011010001000100011;
ROM[2424] <= 32'b00000000110000011010001110000011;
ROM[2425] <= 32'b00000000011100010010000000100011;
ROM[2426] <= 32'b00000000010000010000000100010011;
ROM[2427] <= 32'b11111111110000010000000100010011;
ROM[2428] <= 32'b00000000000000010010001110000011;
ROM[2429] <= 32'b00000000011100011010010000100011;
ROM[2430] <= 32'b00000001000000011010001110000011;
ROM[2431] <= 32'b00000000011100010010000000100011;
ROM[2432] <= 32'b00000000010000010000000100010011;
ROM[2433] <= 32'b00000000000100000000001110010011;
ROM[2434] <= 32'b00000000011100010010000000100011;
ROM[2435] <= 32'b00000000010000010000000100010011;
ROM[2436] <= 32'b11111111110000010000000100010011;
ROM[2437] <= 32'b00000000000000010010001110000011;
ROM[2438] <= 32'b11111111110000010000000100010011;
ROM[2439] <= 32'b00000000000000010010010000000011;
ROM[2440] <= 32'b00000000011101000000001110110011;
ROM[2441] <= 32'b00000000011100010010000000100011;
ROM[2442] <= 32'b00000000010000010000000100010011;
ROM[2443] <= 32'b11111111110000010000000100010011;
ROM[2444] <= 32'b00000000000000010010001110000011;
ROM[2445] <= 32'b00000000011100011010100000100011;
ROM[2446] <= 32'b11010010010111111111000011101111;
ROM[2447] <= 32'b00000000000000000000001110010011;
ROM[2448] <= 32'b00000000011100010010000000100011;
ROM[2449] <= 32'b00000000010000010000000100010011;
ROM[2450] <= 32'b00000001010000000000001110010011;
ROM[2451] <= 32'b01000000011100011000001110110011;
ROM[2452] <= 32'b00000000000000111010000010000011;
ROM[2453] <= 32'b11111111110000010000000100010011;
ROM[2454] <= 32'b00000000000000010010001110000011;
ROM[2455] <= 32'b00000000011100100010000000100011;
ROM[2456] <= 32'b00000000010000100000000100010011;
ROM[2457] <= 32'b00000001010000000000001110010011;
ROM[2458] <= 32'b01000000011100011000001110110011;
ROM[2459] <= 32'b00000000010000111010000110000011;
ROM[2460] <= 32'b00000000100000111010001000000011;
ROM[2461] <= 32'b00000000110000111010001010000011;
ROM[2462] <= 32'b00000001000000111010001100000011;
ROM[2463] <= 32'b00000000000000001000000011100111;
ROM[2464] <= 32'b00000000000000010010000000100011;
ROM[2465] <= 32'b00000000010000010000000100010011;
ROM[2466] <= 32'b00000000000000010010000000100011;
ROM[2467] <= 32'b00000000010000010000000100010011;
ROM[2468] <= 32'b00000000000100000000001110010011;
ROM[2469] <= 32'b00000000011100010010000000100011;
ROM[2470] <= 32'b00000000010000010000000100010011;
ROM[2471] <= 32'b11111111110000010000000100010011;
ROM[2472] <= 32'b00000000000000010010001110000011;
ROM[2473] <= 32'b00000000011100011010000000100011;
ROM[2474] <= 32'b00000000000000000010001110110111;
ROM[2475] <= 32'b01101111010000111000001110010011;
ROM[2476] <= 32'b00000000111000111000001110110011;
ROM[2477] <= 32'b00000000011100010010000000100011;
ROM[2478] <= 32'b00000000010000010000000100010011;
ROM[2479] <= 32'b00000000001100010010000000100011;
ROM[2480] <= 32'b00000000010000010000000100010011;
ROM[2481] <= 32'b00000000010000010010000000100011;
ROM[2482] <= 32'b00000000010000010000000100010011;
ROM[2483] <= 32'b00000000010100010010000000100011;
ROM[2484] <= 32'b00000000010000010000000100010011;
ROM[2485] <= 32'b00000000011000010010000000100011;
ROM[2486] <= 32'b00000000010000010000000100010011;
ROM[2487] <= 32'b00000001010000000000001110010011;
ROM[2488] <= 32'b00000000000000111000001110010011;
ROM[2489] <= 32'b01000000011100010000001110110011;
ROM[2490] <= 32'b00000000011100000000001000110011;
ROM[2491] <= 32'b00000000001000000000000110110011;
ROM[2492] <= 32'b10101101110111111101000011101111;
ROM[2493] <= 32'b11111111110000010000000100010011;
ROM[2494] <= 32'b00000000000000010010001110000011;
ROM[2495] <= 32'b00000000011101100010000000100011;
ROM[2496] <= 32'b00000000000000011010001110000011;
ROM[2497] <= 32'b00000000011100010010000000100011;
ROM[2498] <= 32'b00000000010000010000000100010011;
ROM[2499] <= 32'b00000000000100000000001110010011;
ROM[2500] <= 32'b00000000011100010010000000100011;
ROM[2501] <= 32'b00000000010000010000000100010011;
ROM[2502] <= 32'b11111111110000010000000100010011;
ROM[2503] <= 32'b00000000000000010010001110000011;
ROM[2504] <= 32'b11111111110000010000000100010011;
ROM[2505] <= 32'b00000000000000010010010000000011;
ROM[2506] <= 32'b00000000011101000010010010110011;
ROM[2507] <= 32'b00000000100000111010010100110011;
ROM[2508] <= 32'b00000000101001001000001110110011;
ROM[2509] <= 32'b00000000000100111000001110010011;
ROM[2510] <= 32'b00000000000100111111001110010011;
ROM[2511] <= 32'b00000000011100010010000000100011;
ROM[2512] <= 32'b00000000010000010000000100010011;
ROM[2513] <= 32'b11111111110000010000000100010011;
ROM[2514] <= 32'b00000000000000010010001110000011;
ROM[2515] <= 32'b01000000011100000000001110110011;
ROM[2516] <= 32'b00000000000100111000001110010011;
ROM[2517] <= 32'b00000000011100010010000000100011;
ROM[2518] <= 32'b00000000010000010000000100010011;
ROM[2519] <= 32'b11111111110000010000000100010011;
ROM[2520] <= 32'b00000000000000010010001110000011;
ROM[2521] <= 32'b00000000000000111000101001100011;
ROM[2522] <= 32'b00000000000000000100001110110111;
ROM[2523] <= 32'b11001111000000111000001110010011;
ROM[2524] <= 32'b00000000111000111000001110110011;
ROM[2525] <= 32'b00000000000000111000000011100111;
ROM[2526] <= 32'b00000000000000000010001110110111;
ROM[2527] <= 32'b01111100010000111000001110010011;
ROM[2528] <= 32'b00000000111000111000001110110011;
ROM[2529] <= 32'b00000000011100010010000000100011;
ROM[2530] <= 32'b00000000010000010000000100010011;
ROM[2531] <= 32'b00000000001100010010000000100011;
ROM[2532] <= 32'b00000000010000010000000100010011;
ROM[2533] <= 32'b00000000010000010010000000100011;
ROM[2534] <= 32'b00000000010000010000000100010011;
ROM[2535] <= 32'b00000000010100010010000000100011;
ROM[2536] <= 32'b00000000010000010000000100010011;
ROM[2537] <= 32'b00000000011000010010000000100011;
ROM[2538] <= 32'b00000000010000010000000100010011;
ROM[2539] <= 32'b00000001010000000000001110010011;
ROM[2540] <= 32'b00000000000000111000001110010011;
ROM[2541] <= 32'b01000000011100010000001110110011;
ROM[2542] <= 32'b00000000011100000000001000110011;
ROM[2543] <= 32'b00000000001000000000000110110011;
ROM[2544] <= 32'b00111010100100010100000011101111;
ROM[2545] <= 32'b11111111110000010000000100010011;
ROM[2546] <= 32'b00000000000000010010001110000011;
ROM[2547] <= 32'b00000000011101100010000000100011;
ROM[2548] <= 32'b00000010100100000000001110010011;
ROM[2549] <= 32'b00000000011100010010000000100011;
ROM[2550] <= 32'b00000000010000010000000100010011;
ROM[2551] <= 32'b00000000000000000011001110110111;
ROM[2552] <= 32'b10000010100000111000001110010011;
ROM[2553] <= 32'b00000000111000111000001110110011;
ROM[2554] <= 32'b00000000011100010010000000100011;
ROM[2555] <= 32'b00000000010000010000000100010011;
ROM[2556] <= 32'b00000000001100010010000000100011;
ROM[2557] <= 32'b00000000010000010000000100010011;
ROM[2558] <= 32'b00000000010000010010000000100011;
ROM[2559] <= 32'b00000000010000010000000100010011;
ROM[2560] <= 32'b00000000010100010010000000100011;
ROM[2561] <= 32'b00000000010000010000000100010011;
ROM[2562] <= 32'b00000000011000010010000000100011;
ROM[2563] <= 32'b00000000010000010000000100010011;
ROM[2564] <= 32'b00000001010000000000001110010011;
ROM[2565] <= 32'b00000000010000111000001110010011;
ROM[2566] <= 32'b01000000011100010000001110110011;
ROM[2567] <= 32'b00000000011100000000001000110011;
ROM[2568] <= 32'b00000000001000000000000110110011;
ROM[2569] <= 32'b01110001100100100110000011101111;
ROM[2570] <= 32'b00000100010000000000001110010011;
ROM[2571] <= 32'b00000000011100010010000000100011;
ROM[2572] <= 32'b00000000010000010000000100010011;
ROM[2573] <= 32'b00000000000000000011001110110111;
ROM[2574] <= 32'b10001000000000111000001110010011;
ROM[2575] <= 32'b00000000111000111000001110110011;
ROM[2576] <= 32'b00000000011100010010000000100011;
ROM[2577] <= 32'b00000000010000010000000100010011;
ROM[2578] <= 32'b00000000001100010010000000100011;
ROM[2579] <= 32'b00000000010000010000000100010011;
ROM[2580] <= 32'b00000000010000010010000000100011;
ROM[2581] <= 32'b00000000010000010000000100010011;
ROM[2582] <= 32'b00000000010100010010000000100011;
ROM[2583] <= 32'b00000000010000010000000100010011;
ROM[2584] <= 32'b00000000011000010010000000100011;
ROM[2585] <= 32'b00000000010000010000000100010011;
ROM[2586] <= 32'b00000001010000000000001110010011;
ROM[2587] <= 32'b00000000100000111000001110010011;
ROM[2588] <= 32'b01000000011100010000001110110011;
ROM[2589] <= 32'b00000000011100000000001000110011;
ROM[2590] <= 32'b00000000001000000000000110110011;
ROM[2591] <= 32'b00110011000000100111000011101111;
ROM[2592] <= 32'b00000110111100000000001110010011;
ROM[2593] <= 32'b00000000011100010010000000100011;
ROM[2594] <= 32'b00000000010000010000000100010011;
ROM[2595] <= 32'b00000000000000000011001110110111;
ROM[2596] <= 32'b10001101100000111000001110010011;
ROM[2597] <= 32'b00000000111000111000001110110011;
ROM[2598] <= 32'b00000000011100010010000000100011;
ROM[2599] <= 32'b00000000010000010000000100010011;
ROM[2600] <= 32'b00000000001100010010000000100011;
ROM[2601] <= 32'b00000000010000010000000100010011;
ROM[2602] <= 32'b00000000010000010010000000100011;
ROM[2603] <= 32'b00000000010000010000000100010011;
ROM[2604] <= 32'b00000000010100010010000000100011;
ROM[2605] <= 32'b00000000010000010000000100010011;
ROM[2606] <= 32'b00000000011000010010000000100011;
ROM[2607] <= 32'b00000000010000010000000100010011;
ROM[2608] <= 32'b00000001010000000000001110010011;
ROM[2609] <= 32'b00000000100000111000001110010011;
ROM[2610] <= 32'b01000000011100010000001110110011;
ROM[2611] <= 32'b00000000011100000000001000110011;
ROM[2612] <= 32'b00000000001000000000000110110011;
ROM[2613] <= 32'b00101101100000100111000011101111;
ROM[2614] <= 32'b00000010000000000000001110010011;
ROM[2615] <= 32'b00000000011100010010000000100011;
ROM[2616] <= 32'b00000000010000010000000100010011;
ROM[2617] <= 32'b00000000000000000011001110110111;
ROM[2618] <= 32'b10010011000000111000001110010011;
ROM[2619] <= 32'b00000000111000111000001110110011;
ROM[2620] <= 32'b00000000011100010010000000100011;
ROM[2621] <= 32'b00000000010000010000000100010011;
ROM[2622] <= 32'b00000000001100010010000000100011;
ROM[2623] <= 32'b00000000010000010000000100010011;
ROM[2624] <= 32'b00000000010000010010000000100011;
ROM[2625] <= 32'b00000000010000010000000100010011;
ROM[2626] <= 32'b00000000010100010010000000100011;
ROM[2627] <= 32'b00000000010000010000000100010011;
ROM[2628] <= 32'b00000000011000010010000000100011;
ROM[2629] <= 32'b00000000010000010000000100010011;
ROM[2630] <= 32'b00000001010000000000001110010011;
ROM[2631] <= 32'b00000000100000111000001110010011;
ROM[2632] <= 32'b01000000011100010000001110110011;
ROM[2633] <= 32'b00000000011100000000001000110011;
ROM[2634] <= 32'b00000000001000000000000110110011;
ROM[2635] <= 32'b00101000000000100111000011101111;
ROM[2636] <= 32'b00000111100100000000001110010011;
ROM[2637] <= 32'b00000000011100010010000000100011;
ROM[2638] <= 32'b00000000010000010000000100010011;
ROM[2639] <= 32'b00000000000000000011001110110111;
ROM[2640] <= 32'b10011000100000111000001110010011;
ROM[2641] <= 32'b00000000111000111000001110110011;
ROM[2642] <= 32'b00000000011100010010000000100011;
ROM[2643] <= 32'b00000000010000010000000100010011;
ROM[2644] <= 32'b00000000001100010010000000100011;
ROM[2645] <= 32'b00000000010000010000000100010011;
ROM[2646] <= 32'b00000000010000010010000000100011;
ROM[2647] <= 32'b00000000010000010000000100010011;
ROM[2648] <= 32'b00000000010100010010000000100011;
ROM[2649] <= 32'b00000000010000010000000100010011;
ROM[2650] <= 32'b00000000011000010010000000100011;
ROM[2651] <= 32'b00000000010000010000000100010011;
ROM[2652] <= 32'b00000001010000000000001110010011;
ROM[2653] <= 32'b00000000100000111000001110010011;
ROM[2654] <= 32'b01000000011100010000001110110011;
ROM[2655] <= 32'b00000000011100000000001000110011;
ROM[2656] <= 32'b00000000001000000000000110110011;
ROM[2657] <= 32'b00100010100000100111000011101111;
ROM[2658] <= 32'b00000110111100000000001110010011;
ROM[2659] <= 32'b00000000011100010010000000100011;
ROM[2660] <= 32'b00000000010000010000000100010011;
ROM[2661] <= 32'b00000000000000000011001110110111;
ROM[2662] <= 32'b10011110000000111000001110010011;
ROM[2663] <= 32'b00000000111000111000001110110011;
ROM[2664] <= 32'b00000000011100010010000000100011;
ROM[2665] <= 32'b00000000010000010000000100010011;
ROM[2666] <= 32'b00000000001100010010000000100011;
ROM[2667] <= 32'b00000000010000010000000100010011;
ROM[2668] <= 32'b00000000010000010010000000100011;
ROM[2669] <= 32'b00000000010000010000000100010011;
ROM[2670] <= 32'b00000000010100010010000000100011;
ROM[2671] <= 32'b00000000010000010000000100010011;
ROM[2672] <= 32'b00000000011000010010000000100011;
ROM[2673] <= 32'b00000000010000010000000100010011;
ROM[2674] <= 32'b00000001010000000000001110010011;
ROM[2675] <= 32'b00000000100000111000001110010011;
ROM[2676] <= 32'b01000000011100010000001110110011;
ROM[2677] <= 32'b00000000011100000000001000110011;
ROM[2678] <= 32'b00000000001000000000000110110011;
ROM[2679] <= 32'b00011101000000100111000011101111;
ROM[2680] <= 32'b00000111010100000000001110010011;
ROM[2681] <= 32'b00000000011100010010000000100011;
ROM[2682] <= 32'b00000000010000010000000100010011;
ROM[2683] <= 32'b00000000000000000011001110110111;
ROM[2684] <= 32'b10100011100000111000001110010011;
ROM[2685] <= 32'b00000000111000111000001110110011;
ROM[2686] <= 32'b00000000011100010010000000100011;
ROM[2687] <= 32'b00000000010000010000000100010011;
ROM[2688] <= 32'b00000000001100010010000000100011;
ROM[2689] <= 32'b00000000010000010000000100010011;
ROM[2690] <= 32'b00000000010000010010000000100011;
ROM[2691] <= 32'b00000000010000010000000100010011;
ROM[2692] <= 32'b00000000010100010010000000100011;
ROM[2693] <= 32'b00000000010000010000000100010011;
ROM[2694] <= 32'b00000000011000010010000000100011;
ROM[2695] <= 32'b00000000010000010000000100010011;
ROM[2696] <= 32'b00000001010000000000001110010011;
ROM[2697] <= 32'b00000000100000111000001110010011;
ROM[2698] <= 32'b01000000011100010000001110110011;
ROM[2699] <= 32'b00000000011100000000001000110011;
ROM[2700] <= 32'b00000000001000000000000110110011;
ROM[2701] <= 32'b00010111100000100111000011101111;
ROM[2702] <= 32'b00000010000000000000001110010011;
ROM[2703] <= 32'b00000000011100010010000000100011;
ROM[2704] <= 32'b00000000010000010000000100010011;
ROM[2705] <= 32'b00000000000000000011001110110111;
ROM[2706] <= 32'b10101001000000111000001110010011;
ROM[2707] <= 32'b00000000111000111000001110110011;
ROM[2708] <= 32'b00000000011100010010000000100011;
ROM[2709] <= 32'b00000000010000010000000100010011;
ROM[2710] <= 32'b00000000001100010010000000100011;
ROM[2711] <= 32'b00000000010000010000000100010011;
ROM[2712] <= 32'b00000000010000010010000000100011;
ROM[2713] <= 32'b00000000010000010000000100010011;
ROM[2714] <= 32'b00000000010100010010000000100011;
ROM[2715] <= 32'b00000000010000010000000100010011;
ROM[2716] <= 32'b00000000011000010010000000100011;
ROM[2717] <= 32'b00000000010000010000000100010011;
ROM[2718] <= 32'b00000001010000000000001110010011;
ROM[2719] <= 32'b00000000100000111000001110010011;
ROM[2720] <= 32'b01000000011100010000001110110011;
ROM[2721] <= 32'b00000000011100000000001000110011;
ROM[2722] <= 32'b00000000001000000000000110110011;
ROM[2723] <= 32'b00010010000000100111000011101111;
ROM[2724] <= 32'b00000111011100000000001110010011;
ROM[2725] <= 32'b00000000011100010010000000100011;
ROM[2726] <= 32'b00000000010000010000000100010011;
ROM[2727] <= 32'b00000000000000000011001110110111;
ROM[2728] <= 32'b10101110100000111000001110010011;
ROM[2729] <= 32'b00000000111000111000001110110011;
ROM[2730] <= 32'b00000000011100010010000000100011;
ROM[2731] <= 32'b00000000010000010000000100010011;
ROM[2732] <= 32'b00000000001100010010000000100011;
ROM[2733] <= 32'b00000000010000010000000100010011;
ROM[2734] <= 32'b00000000010000010010000000100011;
ROM[2735] <= 32'b00000000010000010000000100010011;
ROM[2736] <= 32'b00000000010100010010000000100011;
ROM[2737] <= 32'b00000000010000010000000100010011;
ROM[2738] <= 32'b00000000011000010010000000100011;
ROM[2739] <= 32'b00000000010000010000000100010011;
ROM[2740] <= 32'b00000001010000000000001110010011;
ROM[2741] <= 32'b00000000100000111000001110010011;
ROM[2742] <= 32'b01000000011100010000001110110011;
ROM[2743] <= 32'b00000000011100000000001000110011;
ROM[2744] <= 32'b00000000001000000000000110110011;
ROM[2745] <= 32'b00001100100000100111000011101111;
ROM[2746] <= 32'b00000110000100000000001110010011;
ROM[2747] <= 32'b00000000011100010010000000100011;
ROM[2748] <= 32'b00000000010000010000000100010011;
ROM[2749] <= 32'b00000000000000000011001110110111;
ROM[2750] <= 32'b10110100000000111000001110010011;
ROM[2751] <= 32'b00000000111000111000001110110011;
ROM[2752] <= 32'b00000000011100010010000000100011;
ROM[2753] <= 32'b00000000010000010000000100010011;
ROM[2754] <= 32'b00000000001100010010000000100011;
ROM[2755] <= 32'b00000000010000010000000100010011;
ROM[2756] <= 32'b00000000010000010010000000100011;
ROM[2757] <= 32'b00000000010000010000000100010011;
ROM[2758] <= 32'b00000000010100010010000000100011;
ROM[2759] <= 32'b00000000010000010000000100010011;
ROM[2760] <= 32'b00000000011000010010000000100011;
ROM[2761] <= 32'b00000000010000010000000100010011;
ROM[2762] <= 32'b00000001010000000000001110010011;
ROM[2763] <= 32'b00000000100000111000001110010011;
ROM[2764] <= 32'b01000000011100010000001110110011;
ROM[2765] <= 32'b00000000011100000000001000110011;
ROM[2766] <= 32'b00000000001000000000000110110011;
ROM[2767] <= 32'b00000111000000100111000011101111;
ROM[2768] <= 32'b00000110111000000000001110010011;
ROM[2769] <= 32'b00000000011100010010000000100011;
ROM[2770] <= 32'b00000000010000010000000100010011;
ROM[2771] <= 32'b00000000000000000011001110110111;
ROM[2772] <= 32'b10111001100000111000001110010011;
ROM[2773] <= 32'b00000000111000111000001110110011;
ROM[2774] <= 32'b00000000011100010010000000100011;
ROM[2775] <= 32'b00000000010000010000000100010011;
ROM[2776] <= 32'b00000000001100010010000000100011;
ROM[2777] <= 32'b00000000010000010000000100010011;
ROM[2778] <= 32'b00000000010000010010000000100011;
ROM[2779] <= 32'b00000000010000010000000100010011;
ROM[2780] <= 32'b00000000010100010010000000100011;
ROM[2781] <= 32'b00000000010000010000000100010011;
ROM[2782] <= 32'b00000000011000010010000000100011;
ROM[2783] <= 32'b00000000010000010000000100010011;
ROM[2784] <= 32'b00000001010000000000001110010011;
ROM[2785] <= 32'b00000000100000111000001110010011;
ROM[2786] <= 32'b01000000011100010000001110110011;
ROM[2787] <= 32'b00000000011100000000001000110011;
ROM[2788] <= 32'b00000000001000000000000110110011;
ROM[2789] <= 32'b00000001100000100111000011101111;
ROM[2790] <= 32'b00000111010000000000001110010011;
ROM[2791] <= 32'b00000000011100010010000000100011;
ROM[2792] <= 32'b00000000010000010000000100010011;
ROM[2793] <= 32'b00000000000000000011001110110111;
ROM[2794] <= 32'b10111111000000111000001110010011;
ROM[2795] <= 32'b00000000111000111000001110110011;
ROM[2796] <= 32'b00000000011100010010000000100011;
ROM[2797] <= 32'b00000000010000010000000100010011;
ROM[2798] <= 32'b00000000001100010010000000100011;
ROM[2799] <= 32'b00000000010000010000000100010011;
ROM[2800] <= 32'b00000000010000010010000000100011;
ROM[2801] <= 32'b00000000010000010000000100010011;
ROM[2802] <= 32'b00000000010100010010000000100011;
ROM[2803] <= 32'b00000000010000010000000100010011;
ROM[2804] <= 32'b00000000011000010010000000100011;
ROM[2805] <= 32'b00000000010000010000000100010011;
ROM[2806] <= 32'b00000001010000000000001110010011;
ROM[2807] <= 32'b00000000100000111000001110010011;
ROM[2808] <= 32'b01000000011100010000001110110011;
ROM[2809] <= 32'b00000000011100000000001000110011;
ROM[2810] <= 32'b00000000001000000000000110110011;
ROM[2811] <= 32'b01111100000100100110000011101111;
ROM[2812] <= 32'b00000010000000000000001110010011;
ROM[2813] <= 32'b00000000011100010010000000100011;
ROM[2814] <= 32'b00000000010000010000000100010011;
ROM[2815] <= 32'b00000000000000000011001110110111;
ROM[2816] <= 32'b11000100100000111000001110010011;
ROM[2817] <= 32'b00000000111000111000001110110011;
ROM[2818] <= 32'b00000000011100010010000000100011;
ROM[2819] <= 32'b00000000010000010000000100010011;
ROM[2820] <= 32'b00000000001100010010000000100011;
ROM[2821] <= 32'b00000000010000010000000100010011;
ROM[2822] <= 32'b00000000010000010010000000100011;
ROM[2823] <= 32'b00000000010000010000000100010011;
ROM[2824] <= 32'b00000000010100010010000000100011;
ROM[2825] <= 32'b00000000010000010000000100010011;
ROM[2826] <= 32'b00000000011000010010000000100011;
ROM[2827] <= 32'b00000000010000010000000100010011;
ROM[2828] <= 32'b00000001010000000000001110010011;
ROM[2829] <= 32'b00000000100000111000001110010011;
ROM[2830] <= 32'b01000000011100010000001110110011;
ROM[2831] <= 32'b00000000011100000000001000110011;
ROM[2832] <= 32'b00000000001000000000000110110011;
ROM[2833] <= 32'b01110110100100100110000011101111;
ROM[2834] <= 32'b00000111010000000000001110010011;
ROM[2835] <= 32'b00000000011100010010000000100011;
ROM[2836] <= 32'b00000000010000010000000100010011;
ROM[2837] <= 32'b00000000000000000011001110110111;
ROM[2838] <= 32'b11001010000000111000001110010011;
ROM[2839] <= 32'b00000000111000111000001110110011;
ROM[2840] <= 32'b00000000011100010010000000100011;
ROM[2841] <= 32'b00000000010000010000000100010011;
ROM[2842] <= 32'b00000000001100010010000000100011;
ROM[2843] <= 32'b00000000010000010000000100010011;
ROM[2844] <= 32'b00000000010000010010000000100011;
ROM[2845] <= 32'b00000000010000010000000100010011;
ROM[2846] <= 32'b00000000010100010010000000100011;
ROM[2847] <= 32'b00000000010000010000000100010011;
ROM[2848] <= 32'b00000000011000010010000000100011;
ROM[2849] <= 32'b00000000010000010000000100010011;
ROM[2850] <= 32'b00000001010000000000001110010011;
ROM[2851] <= 32'b00000000100000111000001110010011;
ROM[2852] <= 32'b01000000011100010000001110110011;
ROM[2853] <= 32'b00000000011100000000001000110011;
ROM[2854] <= 32'b00000000001000000000000110110011;
ROM[2855] <= 32'b01110001000100100110000011101111;
ROM[2856] <= 32'b00000110111100000000001110010011;
ROM[2857] <= 32'b00000000011100010010000000100011;
ROM[2858] <= 32'b00000000010000010000000100010011;
ROM[2859] <= 32'b00000000000000000011001110110111;
ROM[2860] <= 32'b11001111100000111000001110010011;
ROM[2861] <= 32'b00000000111000111000001110110011;
ROM[2862] <= 32'b00000000011100010010000000100011;
ROM[2863] <= 32'b00000000010000010000000100010011;
ROM[2864] <= 32'b00000000001100010010000000100011;
ROM[2865] <= 32'b00000000010000010000000100010011;
ROM[2866] <= 32'b00000000010000010010000000100011;
ROM[2867] <= 32'b00000000010000010000000100010011;
ROM[2868] <= 32'b00000000010100010010000000100011;
ROM[2869] <= 32'b00000000010000010000000100010011;
ROM[2870] <= 32'b00000000011000010010000000100011;
ROM[2871] <= 32'b00000000010000010000000100010011;
ROM[2872] <= 32'b00000001010000000000001110010011;
ROM[2873] <= 32'b00000000100000111000001110010011;
ROM[2874] <= 32'b01000000011100010000001110110011;
ROM[2875] <= 32'b00000000011100000000001000110011;
ROM[2876] <= 32'b00000000001000000000000110110011;
ROM[2877] <= 32'b01101011100100100110000011101111;
ROM[2878] <= 32'b00000010000000000000001110010011;
ROM[2879] <= 32'b00000000011100010010000000100011;
ROM[2880] <= 32'b00000000010000010000000100010011;
ROM[2881] <= 32'b00000000000000000011001110110111;
ROM[2882] <= 32'b11010101000000111000001110010011;
ROM[2883] <= 32'b00000000111000111000001110110011;
ROM[2884] <= 32'b00000000011100010010000000100011;
ROM[2885] <= 32'b00000000010000010000000100010011;
ROM[2886] <= 32'b00000000001100010010000000100011;
ROM[2887] <= 32'b00000000010000010000000100010011;
ROM[2888] <= 32'b00000000010000010010000000100011;
ROM[2889] <= 32'b00000000010000010000000100010011;
ROM[2890] <= 32'b00000000010100010010000000100011;
ROM[2891] <= 32'b00000000010000010000000100010011;
ROM[2892] <= 32'b00000000011000010010000000100011;
ROM[2893] <= 32'b00000000010000010000000100010011;
ROM[2894] <= 32'b00000001010000000000001110010011;
ROM[2895] <= 32'b00000000100000111000001110010011;
ROM[2896] <= 32'b01000000011100010000001110110011;
ROM[2897] <= 32'b00000000011100000000001000110011;
ROM[2898] <= 32'b00000000001000000000000110110011;
ROM[2899] <= 32'b01100110000100100110000011101111;
ROM[2900] <= 32'b00000110001100000000001110010011;
ROM[2901] <= 32'b00000000011100010010000000100011;
ROM[2902] <= 32'b00000000010000010000000100010011;
ROM[2903] <= 32'b00000000000000000011001110110111;
ROM[2904] <= 32'b11011010100000111000001110010011;
ROM[2905] <= 32'b00000000111000111000001110110011;
ROM[2906] <= 32'b00000000011100010010000000100011;
ROM[2907] <= 32'b00000000010000010000000100010011;
ROM[2908] <= 32'b00000000001100010010000000100011;
ROM[2909] <= 32'b00000000010000010000000100010011;
ROM[2910] <= 32'b00000000010000010010000000100011;
ROM[2911] <= 32'b00000000010000010000000100010011;
ROM[2912] <= 32'b00000000010100010010000000100011;
ROM[2913] <= 32'b00000000010000010000000100010011;
ROM[2914] <= 32'b00000000011000010010000000100011;
ROM[2915] <= 32'b00000000010000010000000100010011;
ROM[2916] <= 32'b00000001010000000000001110010011;
ROM[2917] <= 32'b00000000100000111000001110010011;
ROM[2918] <= 32'b01000000011100010000001110110011;
ROM[2919] <= 32'b00000000011100000000001000110011;
ROM[2920] <= 32'b00000000001000000000000110110011;
ROM[2921] <= 32'b01100000100100100110000011101111;
ROM[2922] <= 32'b00000110111100000000001110010011;
ROM[2923] <= 32'b00000000011100010010000000100011;
ROM[2924] <= 32'b00000000010000010000000100010011;
ROM[2925] <= 32'b00000000000000000011001110110111;
ROM[2926] <= 32'b11100000000000111000001110010011;
ROM[2927] <= 32'b00000000111000111000001110110011;
ROM[2928] <= 32'b00000000011100010010000000100011;
ROM[2929] <= 32'b00000000010000010000000100010011;
ROM[2930] <= 32'b00000000001100010010000000100011;
ROM[2931] <= 32'b00000000010000010000000100010011;
ROM[2932] <= 32'b00000000010000010010000000100011;
ROM[2933] <= 32'b00000000010000010000000100010011;
ROM[2934] <= 32'b00000000010100010010000000100011;
ROM[2935] <= 32'b00000000010000010000000100010011;
ROM[2936] <= 32'b00000000011000010010000000100011;
ROM[2937] <= 32'b00000000010000010000000100010011;
ROM[2938] <= 32'b00000001010000000000001110010011;
ROM[2939] <= 32'b00000000100000111000001110010011;
ROM[2940] <= 32'b01000000011100010000001110110011;
ROM[2941] <= 32'b00000000011100000000001000110011;
ROM[2942] <= 32'b00000000001000000000000110110011;
ROM[2943] <= 32'b01011011000100100110000011101111;
ROM[2944] <= 32'b00000110111000000000001110010011;
ROM[2945] <= 32'b00000000011100010010000000100011;
ROM[2946] <= 32'b00000000010000010000000100010011;
ROM[2947] <= 32'b00000000000000000011001110110111;
ROM[2948] <= 32'b11100101100000111000001110010011;
ROM[2949] <= 32'b00000000111000111000001110110011;
ROM[2950] <= 32'b00000000011100010010000000100011;
ROM[2951] <= 32'b00000000010000010000000100010011;
ROM[2952] <= 32'b00000000001100010010000000100011;
ROM[2953] <= 32'b00000000010000010000000100010011;
ROM[2954] <= 32'b00000000010000010010000000100011;
ROM[2955] <= 32'b00000000010000010000000100010011;
ROM[2956] <= 32'b00000000010100010010000000100011;
ROM[2957] <= 32'b00000000010000010000000100010011;
ROM[2958] <= 32'b00000000011000010010000000100011;
ROM[2959] <= 32'b00000000010000010000000100010011;
ROM[2960] <= 32'b00000001010000000000001110010011;
ROM[2961] <= 32'b00000000100000111000001110010011;
ROM[2962] <= 32'b01000000011100010000001110110011;
ROM[2963] <= 32'b00000000011100000000001000110011;
ROM[2964] <= 32'b00000000001000000000000110110011;
ROM[2965] <= 32'b01010101100100100110000011101111;
ROM[2966] <= 32'b00000111010000000000001110010011;
ROM[2967] <= 32'b00000000011100010010000000100011;
ROM[2968] <= 32'b00000000010000010000000100010011;
ROM[2969] <= 32'b00000000000000000011001110110111;
ROM[2970] <= 32'b11101011000000111000001110010011;
ROM[2971] <= 32'b00000000111000111000001110110011;
ROM[2972] <= 32'b00000000011100010010000000100011;
ROM[2973] <= 32'b00000000010000010000000100010011;
ROM[2974] <= 32'b00000000001100010010000000100011;
ROM[2975] <= 32'b00000000010000010000000100010011;
ROM[2976] <= 32'b00000000010000010010000000100011;
ROM[2977] <= 32'b00000000010000010000000100010011;
ROM[2978] <= 32'b00000000010100010010000000100011;
ROM[2979] <= 32'b00000000010000010000000100010011;
ROM[2980] <= 32'b00000000011000010010000000100011;
ROM[2981] <= 32'b00000000010000010000000100010011;
ROM[2982] <= 32'b00000001010000000000001110010011;
ROM[2983] <= 32'b00000000100000111000001110010011;
ROM[2984] <= 32'b01000000011100010000001110110011;
ROM[2985] <= 32'b00000000011100000000001000110011;
ROM[2986] <= 32'b00000000001000000000000110110011;
ROM[2987] <= 32'b01010000000100100110000011101111;
ROM[2988] <= 32'b00000110100100000000001110010011;
ROM[2989] <= 32'b00000000011100010010000000100011;
ROM[2990] <= 32'b00000000010000010000000100010011;
ROM[2991] <= 32'b00000000000000000011001110110111;
ROM[2992] <= 32'b11110000100000111000001110010011;
ROM[2993] <= 32'b00000000111000111000001110110011;
ROM[2994] <= 32'b00000000011100010010000000100011;
ROM[2995] <= 32'b00000000010000010000000100010011;
ROM[2996] <= 32'b00000000001100010010000000100011;
ROM[2997] <= 32'b00000000010000010000000100010011;
ROM[2998] <= 32'b00000000010000010010000000100011;
ROM[2999] <= 32'b00000000010000010000000100010011;
ROM[3000] <= 32'b00000000010100010010000000100011;
ROM[3001] <= 32'b00000000010000010000000100010011;
ROM[3002] <= 32'b00000000011000010010000000100011;
ROM[3003] <= 32'b00000000010000010000000100010011;
ROM[3004] <= 32'b00000001010000000000001110010011;
ROM[3005] <= 32'b00000000100000111000001110010011;
ROM[3006] <= 32'b01000000011100010000001110110011;
ROM[3007] <= 32'b00000000011100000000001000110011;
ROM[3008] <= 32'b00000000001000000000000110110011;
ROM[3009] <= 32'b01001010100100100110000011101111;
ROM[3010] <= 32'b00000110111000000000001110010011;
ROM[3011] <= 32'b00000000011100010010000000100011;
ROM[3012] <= 32'b00000000010000010000000100010011;
ROM[3013] <= 32'b00000000000000000011001110110111;
ROM[3014] <= 32'b11110110000000111000001110010011;
ROM[3015] <= 32'b00000000111000111000001110110011;
ROM[3016] <= 32'b00000000011100010010000000100011;
ROM[3017] <= 32'b00000000010000010000000100010011;
ROM[3018] <= 32'b00000000001100010010000000100011;
ROM[3019] <= 32'b00000000010000010000000100010011;
ROM[3020] <= 32'b00000000010000010010000000100011;
ROM[3021] <= 32'b00000000010000010000000100010011;
ROM[3022] <= 32'b00000000010100010010000000100011;
ROM[3023] <= 32'b00000000010000010000000100010011;
ROM[3024] <= 32'b00000000011000010010000000100011;
ROM[3025] <= 32'b00000000010000010000000100010011;
ROM[3026] <= 32'b00000001010000000000001110010011;
ROM[3027] <= 32'b00000000100000111000001110010011;
ROM[3028] <= 32'b01000000011100010000001110110011;
ROM[3029] <= 32'b00000000011100000000001000110011;
ROM[3030] <= 32'b00000000001000000000000110110011;
ROM[3031] <= 32'b01000101000100100110000011101111;
ROM[3032] <= 32'b00000111010100000000001110010011;
ROM[3033] <= 32'b00000000011100010010000000100011;
ROM[3034] <= 32'b00000000010000010000000100010011;
ROM[3035] <= 32'b00000000000000000011001110110111;
ROM[3036] <= 32'b11111011100000111000001110010011;
ROM[3037] <= 32'b00000000111000111000001110110011;
ROM[3038] <= 32'b00000000011100010010000000100011;
ROM[3039] <= 32'b00000000010000010000000100010011;
ROM[3040] <= 32'b00000000001100010010000000100011;
ROM[3041] <= 32'b00000000010000010000000100010011;
ROM[3042] <= 32'b00000000010000010010000000100011;
ROM[3043] <= 32'b00000000010000010000000100010011;
ROM[3044] <= 32'b00000000010100010010000000100011;
ROM[3045] <= 32'b00000000010000010000000100010011;
ROM[3046] <= 32'b00000000011000010010000000100011;
ROM[3047] <= 32'b00000000010000010000000100010011;
ROM[3048] <= 32'b00000001010000000000001110010011;
ROM[3049] <= 32'b00000000100000111000001110010011;
ROM[3050] <= 32'b01000000011100010000001110110011;
ROM[3051] <= 32'b00000000011100000000001000110011;
ROM[3052] <= 32'b00000000001000000000000110110011;
ROM[3053] <= 32'b00111111100100100110000011101111;
ROM[3054] <= 32'b00000110010100000000001110010011;
ROM[3055] <= 32'b00000000011100010010000000100011;
ROM[3056] <= 32'b00000000010000010000000100010011;
ROM[3057] <= 32'b00000000000000000011001110110111;
ROM[3058] <= 32'b00000001000000111000001110010011;
ROM[3059] <= 32'b00000000111000111000001110110011;
ROM[3060] <= 32'b00000000011100010010000000100011;
ROM[3061] <= 32'b00000000010000010000000100010011;
ROM[3062] <= 32'b00000000001100010010000000100011;
ROM[3063] <= 32'b00000000010000010000000100010011;
ROM[3064] <= 32'b00000000010000010010000000100011;
ROM[3065] <= 32'b00000000010000010000000100010011;
ROM[3066] <= 32'b00000000010100010010000000100011;
ROM[3067] <= 32'b00000000010000010000000100010011;
ROM[3068] <= 32'b00000000011000010010000000100011;
ROM[3069] <= 32'b00000000010000010000000100010011;
ROM[3070] <= 32'b00000001010000000000001110010011;
ROM[3071] <= 32'b00000000100000111000001110010011;
ROM[3072] <= 32'b01000000011100010000001110110011;
ROM[3073] <= 32'b00000000011100000000001000110011;
ROM[3074] <= 32'b00000000001000000000000110110011;
ROM[3075] <= 32'b00111010000100100110000011101111;
ROM[3076] <= 32'b00000011111100000000001110010011;
ROM[3077] <= 32'b00000000011100010010000000100011;
ROM[3078] <= 32'b00000000010000010000000100010011;
ROM[3079] <= 32'b00000000000000000011001110110111;
ROM[3080] <= 32'b00000110100000111000001110010011;
ROM[3081] <= 32'b00000000111000111000001110110011;
ROM[3082] <= 32'b00000000011100010010000000100011;
ROM[3083] <= 32'b00000000010000010000000100010011;
ROM[3084] <= 32'b00000000001100010010000000100011;
ROM[3085] <= 32'b00000000010000010000000100010011;
ROM[3086] <= 32'b00000000010000010010000000100011;
ROM[3087] <= 32'b00000000010000010000000100010011;
ROM[3088] <= 32'b00000000010100010010000000100011;
ROM[3089] <= 32'b00000000010000010000000100010011;
ROM[3090] <= 32'b00000000011000010010000000100011;
ROM[3091] <= 32'b00000000010000010000000100010011;
ROM[3092] <= 32'b00000001010000000000001110010011;
ROM[3093] <= 32'b00000000100000111000001110010011;
ROM[3094] <= 32'b01000000011100010000001110110011;
ROM[3095] <= 32'b00000000011100000000001000110011;
ROM[3096] <= 32'b00000000001000000000000110110011;
ROM[3097] <= 32'b00110100100100100110000011101111;
ROM[3098] <= 32'b00000010000000000000001110010011;
ROM[3099] <= 32'b00000000011100010010000000100011;
ROM[3100] <= 32'b00000000010000010000000100010011;
ROM[3101] <= 32'b00000000000000000011001110110111;
ROM[3102] <= 32'b00001100000000111000001110010011;
ROM[3103] <= 32'b00000000111000111000001110110011;
ROM[3104] <= 32'b00000000011100010010000000100011;
ROM[3105] <= 32'b00000000010000010000000100010011;
ROM[3106] <= 32'b00000000001100010010000000100011;
ROM[3107] <= 32'b00000000010000010000000100010011;
ROM[3108] <= 32'b00000000010000010010000000100011;
ROM[3109] <= 32'b00000000010000010000000100010011;
ROM[3110] <= 32'b00000000010100010010000000100011;
ROM[3111] <= 32'b00000000010000010000000100010011;
ROM[3112] <= 32'b00000000011000010010000000100011;
ROM[3113] <= 32'b00000000010000010000000100010011;
ROM[3114] <= 32'b00000001010000000000001110010011;
ROM[3115] <= 32'b00000000100000111000001110010011;
ROM[3116] <= 32'b01000000011100010000001110110011;
ROM[3117] <= 32'b00000000011100000000001000110011;
ROM[3118] <= 32'b00000000001000000000000110110011;
ROM[3119] <= 32'b00101111000100100110000011101111;
ROM[3120] <= 32'b00000010100000000000001110010011;
ROM[3121] <= 32'b00000000011100010010000000100011;
ROM[3122] <= 32'b00000000010000010000000100010011;
ROM[3123] <= 32'b00000000000000000011001110110111;
ROM[3124] <= 32'b00010001100000111000001110010011;
ROM[3125] <= 32'b00000000111000111000001110110011;
ROM[3126] <= 32'b00000000011100010010000000100011;
ROM[3127] <= 32'b00000000010000010000000100010011;
ROM[3128] <= 32'b00000000001100010010000000100011;
ROM[3129] <= 32'b00000000010000010000000100010011;
ROM[3130] <= 32'b00000000010000010010000000100011;
ROM[3131] <= 32'b00000000010000010000000100010011;
ROM[3132] <= 32'b00000000010100010010000000100011;
ROM[3133] <= 32'b00000000010000010000000100010011;
ROM[3134] <= 32'b00000000011000010010000000100011;
ROM[3135] <= 32'b00000000010000010000000100010011;
ROM[3136] <= 32'b00000001010000000000001110010011;
ROM[3137] <= 32'b00000000100000111000001110010011;
ROM[3138] <= 32'b01000000011100010000001110110011;
ROM[3139] <= 32'b00000000011100000000001000110011;
ROM[3140] <= 32'b00000000001000000000000110110011;
ROM[3141] <= 32'b00101001100100100110000011101111;
ROM[3142] <= 32'b00000111100100000000001110010011;
ROM[3143] <= 32'b00000000011100010010000000100011;
ROM[3144] <= 32'b00000000010000010000000100010011;
ROM[3145] <= 32'b00000000000000000011001110110111;
ROM[3146] <= 32'b00010111000000111000001110010011;
ROM[3147] <= 32'b00000000111000111000001110110011;
ROM[3148] <= 32'b00000000011100010010000000100011;
ROM[3149] <= 32'b00000000010000010000000100010011;
ROM[3150] <= 32'b00000000001100010010000000100011;
ROM[3151] <= 32'b00000000010000010000000100010011;
ROM[3152] <= 32'b00000000010000010010000000100011;
ROM[3153] <= 32'b00000000010000010000000100010011;
ROM[3154] <= 32'b00000000010100010010000000100011;
ROM[3155] <= 32'b00000000010000010000000100010011;
ROM[3156] <= 32'b00000000011000010010000000100011;
ROM[3157] <= 32'b00000000010000010000000100010011;
ROM[3158] <= 32'b00000001010000000000001110010011;
ROM[3159] <= 32'b00000000100000111000001110010011;
ROM[3160] <= 32'b01000000011100010000001110110011;
ROM[3161] <= 32'b00000000011100000000001000110011;
ROM[3162] <= 32'b00000000001000000000000110110011;
ROM[3163] <= 32'b00100100000100100110000011101111;
ROM[3164] <= 32'b00000110010100000000001110010011;
ROM[3165] <= 32'b00000000011100010010000000100011;
ROM[3166] <= 32'b00000000010000010000000100010011;
ROM[3167] <= 32'b00000000000000000011001110110111;
ROM[3168] <= 32'b00011100100000111000001110010011;
ROM[3169] <= 32'b00000000111000111000001110110011;
ROM[3170] <= 32'b00000000011100010010000000100011;
ROM[3171] <= 32'b00000000010000010000000100010011;
ROM[3172] <= 32'b00000000001100010010000000100011;
ROM[3173] <= 32'b00000000010000010000000100010011;
ROM[3174] <= 32'b00000000010000010010000000100011;
ROM[3175] <= 32'b00000000010000010000000100010011;
ROM[3176] <= 32'b00000000010100010010000000100011;
ROM[3177] <= 32'b00000000010000010000000100010011;
ROM[3178] <= 32'b00000000011000010010000000100011;
ROM[3179] <= 32'b00000000010000010000000100010011;
ROM[3180] <= 32'b00000001010000000000001110010011;
ROM[3181] <= 32'b00000000100000111000001110010011;
ROM[3182] <= 32'b01000000011100010000001110110011;
ROM[3183] <= 32'b00000000011100000000001000110011;
ROM[3184] <= 32'b00000000001000000000000110110011;
ROM[3185] <= 32'b00011110100100100110000011101111;
ROM[3186] <= 32'b00000111001100000000001110010011;
ROM[3187] <= 32'b00000000011100010010000000100011;
ROM[3188] <= 32'b00000000010000010000000100010011;
ROM[3189] <= 32'b00000000000000000011001110110111;
ROM[3190] <= 32'b00100010000000111000001110010011;
ROM[3191] <= 32'b00000000111000111000001110110011;
ROM[3192] <= 32'b00000000011100010010000000100011;
ROM[3193] <= 32'b00000000010000010000000100010011;
ROM[3194] <= 32'b00000000001100010010000000100011;
ROM[3195] <= 32'b00000000010000010000000100010011;
ROM[3196] <= 32'b00000000010000010010000000100011;
ROM[3197] <= 32'b00000000010000010000000100010011;
ROM[3198] <= 32'b00000000010100010010000000100011;
ROM[3199] <= 32'b00000000010000010000000100010011;
ROM[3200] <= 32'b00000000011000010010000000100011;
ROM[3201] <= 32'b00000000010000010000000100010011;
ROM[3202] <= 32'b00000001010000000000001110010011;
ROM[3203] <= 32'b00000000100000111000001110010011;
ROM[3204] <= 32'b01000000011100010000001110110011;
ROM[3205] <= 32'b00000000011100000000001000110011;
ROM[3206] <= 32'b00000000001000000000000110110011;
ROM[3207] <= 32'b00011001000100100110000011101111;
ROM[3208] <= 32'b00000010100000000000001110010011;
ROM[3209] <= 32'b00000000011100010010000000100011;
ROM[3210] <= 32'b00000000010000010000000100010011;
ROM[3211] <= 32'b00000000000000000011001110110111;
ROM[3212] <= 32'b00100111100000111000001110010011;
ROM[3213] <= 32'b00000000111000111000001110110011;
ROM[3214] <= 32'b00000000011100010010000000100011;
ROM[3215] <= 32'b00000000010000010000000100010011;
ROM[3216] <= 32'b00000000001100010010000000100011;
ROM[3217] <= 32'b00000000010000010000000100010011;
ROM[3218] <= 32'b00000000010000010010000000100011;
ROM[3219] <= 32'b00000000010000010000000100010011;
ROM[3220] <= 32'b00000000010100010010000000100011;
ROM[3221] <= 32'b00000000010000010000000100010011;
ROM[3222] <= 32'b00000000011000010010000000100011;
ROM[3223] <= 32'b00000000010000010000000100010011;
ROM[3224] <= 32'b00000001010000000000001110010011;
ROM[3225] <= 32'b00000000100000111000001110010011;
ROM[3226] <= 32'b01000000011100010000001110110011;
ROM[3227] <= 32'b00000000011100000000001000110011;
ROM[3228] <= 32'b00000000001000000000000110110011;
ROM[3229] <= 32'b00010011100100100110000011101111;
ROM[3230] <= 32'b00000011000100000000001110010011;
ROM[3231] <= 32'b00000000011100010010000000100011;
ROM[3232] <= 32'b00000000010000010000000100010011;
ROM[3233] <= 32'b00000000000000000011001110110111;
ROM[3234] <= 32'b00101101000000111000001110010011;
ROM[3235] <= 32'b00000000111000111000001110110011;
ROM[3236] <= 32'b00000000011100010010000000100011;
ROM[3237] <= 32'b00000000010000010000000100010011;
ROM[3238] <= 32'b00000000001100010010000000100011;
ROM[3239] <= 32'b00000000010000010000000100010011;
ROM[3240] <= 32'b00000000010000010010000000100011;
ROM[3241] <= 32'b00000000010000010000000100010011;
ROM[3242] <= 32'b00000000010100010010000000100011;
ROM[3243] <= 32'b00000000010000010000000100010011;
ROM[3244] <= 32'b00000000011000010010000000100011;
ROM[3245] <= 32'b00000000010000010000000100010011;
ROM[3246] <= 32'b00000001010000000000001110010011;
ROM[3247] <= 32'b00000000100000111000001110010011;
ROM[3248] <= 32'b01000000011100010000001110110011;
ROM[3249] <= 32'b00000000011100000000001000110011;
ROM[3250] <= 32'b00000000001000000000000110110011;
ROM[3251] <= 32'b00001110000100100110000011101111;
ROM[3252] <= 32'b00000010100100000000001110010011;
ROM[3253] <= 32'b00000000011100010010000000100011;
ROM[3254] <= 32'b00000000010000010000000100010011;
ROM[3255] <= 32'b00000000000000000011001110110111;
ROM[3256] <= 32'b00110010100000111000001110010011;
ROM[3257] <= 32'b00000000111000111000001110110011;
ROM[3258] <= 32'b00000000011100010010000000100011;
ROM[3259] <= 32'b00000000010000010000000100010011;
ROM[3260] <= 32'b00000000001100010010000000100011;
ROM[3261] <= 32'b00000000010000010000000100010011;
ROM[3262] <= 32'b00000000010000010010000000100011;
ROM[3263] <= 32'b00000000010000010000000100010011;
ROM[3264] <= 32'b00000000010100010010000000100011;
ROM[3265] <= 32'b00000000010000010000000100010011;
ROM[3266] <= 32'b00000000011000010010000000100011;
ROM[3267] <= 32'b00000000010000010000000100010011;
ROM[3268] <= 32'b00000001010000000000001110010011;
ROM[3269] <= 32'b00000000100000111000001110010011;
ROM[3270] <= 32'b01000000011100010000001110110011;
ROM[3271] <= 32'b00000000011100000000001000110011;
ROM[3272] <= 32'b00000000001000000000000110110011;
ROM[3273] <= 32'b00001000100100100110000011101111;
ROM[3274] <= 32'b00000010111100000000001110010011;
ROM[3275] <= 32'b00000000011100010010000000100011;
ROM[3276] <= 32'b00000000010000010000000100010011;
ROM[3277] <= 32'b00000000000000000011001110110111;
ROM[3278] <= 32'b00111000000000111000001110010011;
ROM[3279] <= 32'b00000000111000111000001110110011;
ROM[3280] <= 32'b00000000011100010010000000100011;
ROM[3281] <= 32'b00000000010000010000000100010011;
ROM[3282] <= 32'b00000000001100010010000000100011;
ROM[3283] <= 32'b00000000010000010000000100010011;
ROM[3284] <= 32'b00000000010000010010000000100011;
ROM[3285] <= 32'b00000000010000010000000100010011;
ROM[3286] <= 32'b00000000010100010010000000100011;
ROM[3287] <= 32'b00000000010000010000000100010011;
ROM[3288] <= 32'b00000000011000010010000000100011;
ROM[3289] <= 32'b00000000010000010000000100010011;
ROM[3290] <= 32'b00000001010000000000001110010011;
ROM[3291] <= 32'b00000000100000111000001110010011;
ROM[3292] <= 32'b01000000011100010000001110110011;
ROM[3293] <= 32'b00000000011100000000001000110011;
ROM[3294] <= 32'b00000000001000000000000110110011;
ROM[3295] <= 32'b00000011000100100110000011101111;
ROM[3296] <= 32'b00000110111000000000001110010011;
ROM[3297] <= 32'b00000000011100010010000000100011;
ROM[3298] <= 32'b00000000010000010000000100010011;
ROM[3299] <= 32'b00000000000000000011001110110111;
ROM[3300] <= 32'b00111101100000111000001110010011;
ROM[3301] <= 32'b00000000111000111000001110110011;
ROM[3302] <= 32'b00000000011100010010000000100011;
ROM[3303] <= 32'b00000000010000010000000100010011;
ROM[3304] <= 32'b00000000001100010010000000100011;
ROM[3305] <= 32'b00000000010000010000000100010011;
ROM[3306] <= 32'b00000000010000010010000000100011;
ROM[3307] <= 32'b00000000010000010000000100010011;
ROM[3308] <= 32'b00000000010100010010000000100011;
ROM[3309] <= 32'b00000000010000010000000100010011;
ROM[3310] <= 32'b00000000011000010010000000100011;
ROM[3311] <= 32'b00000000010000010000000100010011;
ROM[3312] <= 32'b00000001010000000000001110010011;
ROM[3313] <= 32'b00000000100000111000001110010011;
ROM[3314] <= 32'b01000000011100010000001110110011;
ROM[3315] <= 32'b00000000011100000000001000110011;
ROM[3316] <= 32'b00000000001000000000000110110011;
ROM[3317] <= 32'b01111101100000100110000011101111;
ROM[3318] <= 32'b00000110111100000000001110010011;
ROM[3319] <= 32'b00000000011100010010000000100011;
ROM[3320] <= 32'b00000000010000010000000100010011;
ROM[3321] <= 32'b00000000000000000011001110110111;
ROM[3322] <= 32'b01000011000000111000001110010011;
ROM[3323] <= 32'b00000000111000111000001110110011;
ROM[3324] <= 32'b00000000011100010010000000100011;
ROM[3325] <= 32'b00000000010000010000000100010011;
ROM[3326] <= 32'b00000000001100010010000000100011;
ROM[3327] <= 32'b00000000010000010000000100010011;
ROM[3328] <= 32'b00000000010000010010000000100011;
ROM[3329] <= 32'b00000000010000010000000100010011;
ROM[3330] <= 32'b00000000010100010010000000100011;
ROM[3331] <= 32'b00000000010000010000000100010011;
ROM[3332] <= 32'b00000000011000010010000000100011;
ROM[3333] <= 32'b00000000010000010000000100010011;
ROM[3334] <= 32'b00000001010000000000001110010011;
ROM[3335] <= 32'b00000000100000111000001110010011;
ROM[3336] <= 32'b01000000011100010000001110110011;
ROM[3337] <= 32'b00000000011100000000001000110011;
ROM[3338] <= 32'b00000000001000000000000110110011;
ROM[3339] <= 32'b01111000000000100110000011101111;
ROM[3340] <= 32'b00000010100000000000001110010011;
ROM[3341] <= 32'b00000000011100010010000000100011;
ROM[3342] <= 32'b00000000010000010000000100010011;
ROM[3343] <= 32'b00000000000000000011001110110111;
ROM[3344] <= 32'b01001000100000111000001110010011;
ROM[3345] <= 32'b00000000111000111000001110110011;
ROM[3346] <= 32'b00000000011100010010000000100011;
ROM[3347] <= 32'b00000000010000010000000100010011;
ROM[3348] <= 32'b00000000001100010010000000100011;
ROM[3349] <= 32'b00000000010000010000000100010011;
ROM[3350] <= 32'b00000000010000010010000000100011;
ROM[3351] <= 32'b00000000010000010000000100010011;
ROM[3352] <= 32'b00000000010100010010000000100011;
ROM[3353] <= 32'b00000000010000010000000100010011;
ROM[3354] <= 32'b00000000011000010010000000100011;
ROM[3355] <= 32'b00000000010000010000000100010011;
ROM[3356] <= 32'b00000001010000000000001110010011;
ROM[3357] <= 32'b00000000100000111000001110010011;
ROM[3358] <= 32'b01000000011100010000001110110011;
ROM[3359] <= 32'b00000000011100000000001000110011;
ROM[3360] <= 32'b00000000001000000000000110110011;
ROM[3361] <= 32'b01110010100000100110000011101111;
ROM[3362] <= 32'b00000011000000000000001110010011;
ROM[3363] <= 32'b00000000011100010010000000100011;
ROM[3364] <= 32'b00000000010000010000000100010011;
ROM[3365] <= 32'b00000000000000000011001110110111;
ROM[3366] <= 32'b01001110000000111000001110010011;
ROM[3367] <= 32'b00000000111000111000001110110011;
ROM[3368] <= 32'b00000000011100010010000000100011;
ROM[3369] <= 32'b00000000010000010000000100010011;
ROM[3370] <= 32'b00000000001100010010000000100011;
ROM[3371] <= 32'b00000000010000010000000100010011;
ROM[3372] <= 32'b00000000010000010010000000100011;
ROM[3373] <= 32'b00000000010000010000000100010011;
ROM[3374] <= 32'b00000000010100010010000000100011;
ROM[3375] <= 32'b00000000010000010000000100010011;
ROM[3376] <= 32'b00000000011000010010000000100011;
ROM[3377] <= 32'b00000000010000010000000100010011;
ROM[3378] <= 32'b00000001010000000000001110010011;
ROM[3379] <= 32'b00000000100000111000001110010011;
ROM[3380] <= 32'b01000000011100010000001110110011;
ROM[3381] <= 32'b00000000011100000000001000110011;
ROM[3382] <= 32'b00000000001000000000000110110011;
ROM[3383] <= 32'b01101101000000100110000011101111;
ROM[3384] <= 32'b00000010100100000000001110010011;
ROM[3385] <= 32'b00000000011100010010000000100011;
ROM[3386] <= 32'b00000000010000010000000100010011;
ROM[3387] <= 32'b00000000000000000011001110110111;
ROM[3388] <= 32'b01010011100000111000001110010011;
ROM[3389] <= 32'b00000000111000111000001110110011;
ROM[3390] <= 32'b00000000011100010010000000100011;
ROM[3391] <= 32'b00000000010000010000000100010011;
ROM[3392] <= 32'b00000000001100010010000000100011;
ROM[3393] <= 32'b00000000010000010000000100010011;
ROM[3394] <= 32'b00000000010000010010000000100011;
ROM[3395] <= 32'b00000000010000010000000100010011;
ROM[3396] <= 32'b00000000010100010010000000100011;
ROM[3397] <= 32'b00000000010000010000000100010011;
ROM[3398] <= 32'b00000000011000010010000000100011;
ROM[3399] <= 32'b00000000010000010000000100010011;
ROM[3400] <= 32'b00000001010000000000001110010011;
ROM[3401] <= 32'b00000000100000111000001110010011;
ROM[3402] <= 32'b01000000011100010000001110110011;
ROM[3403] <= 32'b00000000011100000000001000110011;
ROM[3404] <= 32'b00000000001000000000000110110011;
ROM[3405] <= 32'b01100111100000100110000011101111;
ROM[3406] <= 32'b00000010100100000000001110010011;
ROM[3407] <= 32'b00000000011100010010000000100011;
ROM[3408] <= 32'b00000000010000010000000100010011;
ROM[3409] <= 32'b00000000000000000011001110110111;
ROM[3410] <= 32'b01011001000000111000001110010011;
ROM[3411] <= 32'b00000000111000111000001110110011;
ROM[3412] <= 32'b00000000011100010010000000100011;
ROM[3413] <= 32'b00000000010000010000000100010011;
ROM[3414] <= 32'b00000000001100010010000000100011;
ROM[3415] <= 32'b00000000010000010000000100010011;
ROM[3416] <= 32'b00000000010000010010000000100011;
ROM[3417] <= 32'b00000000010000010000000100010011;
ROM[3418] <= 32'b00000000010100010010000000100011;
ROM[3419] <= 32'b00000000010000010000000100010011;
ROM[3420] <= 32'b00000000011000010010000000100011;
ROM[3421] <= 32'b00000000010000010000000100010011;
ROM[3422] <= 32'b00000001010000000000001110010011;
ROM[3423] <= 32'b00000000100000111000001110010011;
ROM[3424] <= 32'b01000000011100010000001110110011;
ROM[3425] <= 32'b00000000011100000000001000110011;
ROM[3426] <= 32'b00000000001000000000000110110011;
ROM[3427] <= 32'b01100010000000100110000011101111;
ROM[3428] <= 32'b00000011101000000000001110010011;
ROM[3429] <= 32'b00000000011100010010000000100011;
ROM[3430] <= 32'b00000000010000010000000100010011;
ROM[3431] <= 32'b00000000000000000011001110110111;
ROM[3432] <= 32'b01011110100000111000001110010011;
ROM[3433] <= 32'b00000000111000111000001110110011;
ROM[3434] <= 32'b00000000011100010010000000100011;
ROM[3435] <= 32'b00000000010000010000000100010011;
ROM[3436] <= 32'b00000000001100010010000000100011;
ROM[3437] <= 32'b00000000010000010000000100010011;
ROM[3438] <= 32'b00000000010000010010000000100011;
ROM[3439] <= 32'b00000000010000010000000100010011;
ROM[3440] <= 32'b00000000010100010010000000100011;
ROM[3441] <= 32'b00000000010000010000000100010011;
ROM[3442] <= 32'b00000000011000010010000000100011;
ROM[3443] <= 32'b00000000010000010000000100010011;
ROM[3444] <= 32'b00000001010000000000001110010011;
ROM[3445] <= 32'b00000000100000111000001110010011;
ROM[3446] <= 32'b01000000011100010000001110110011;
ROM[3447] <= 32'b00000000011100000000001000110011;
ROM[3448] <= 32'b00000000001000000000000110110011;
ROM[3449] <= 32'b01011100100000100110000011101111;
ROM[3450] <= 32'b00000010000000000000001110010011;
ROM[3451] <= 32'b00000000011100010010000000100011;
ROM[3452] <= 32'b00000000010000010000000100010011;
ROM[3453] <= 32'b00000000000000000011001110110111;
ROM[3454] <= 32'b01100100000000111000001110010011;
ROM[3455] <= 32'b00000000111000111000001110110011;
ROM[3456] <= 32'b00000000011100010010000000100011;
ROM[3457] <= 32'b00000000010000010000000100010011;
ROM[3458] <= 32'b00000000001100010010000000100011;
ROM[3459] <= 32'b00000000010000010000000100010011;
ROM[3460] <= 32'b00000000010000010010000000100011;
ROM[3461] <= 32'b00000000010000010000000100010011;
ROM[3462] <= 32'b00000000010100010010000000100011;
ROM[3463] <= 32'b00000000010000010000000100010011;
ROM[3464] <= 32'b00000000011000010010000000100011;
ROM[3465] <= 32'b00000000010000010000000100010011;
ROM[3466] <= 32'b00000001010000000000001110010011;
ROM[3467] <= 32'b00000000100000111000001110010011;
ROM[3468] <= 32'b01000000011100010000001110110011;
ROM[3469] <= 32'b00000000011100000000001000110011;
ROM[3470] <= 32'b00000000001000000000000110110011;
ROM[3471] <= 32'b01010111000000100110000011101111;
ROM[3472] <= 32'b00000000000000000011001110110111;
ROM[3473] <= 32'b01101000110000111000001110010011;
ROM[3474] <= 32'b00000000111000111000001110110011;
ROM[3475] <= 32'b00000000011100010010000000100011;
ROM[3476] <= 32'b00000000010000010000000100010011;
ROM[3477] <= 32'b00000000001100010010000000100011;
ROM[3478] <= 32'b00000000010000010000000100010011;
ROM[3479] <= 32'b00000000010000010010000000100011;
ROM[3480] <= 32'b00000000010000010000000100010011;
ROM[3481] <= 32'b00000000010100010010000000100011;
ROM[3482] <= 32'b00000000010000010000000100010011;
ROM[3483] <= 32'b00000000011000010010000000100011;
ROM[3484] <= 32'b00000000010000010000000100010011;
ROM[3485] <= 32'b00000001010000000000001110010011;
ROM[3486] <= 32'b00000000010000111000001110010011;
ROM[3487] <= 32'b01000000011100010000001110110011;
ROM[3488] <= 32'b00000000011100000000001000110011;
ROM[3489] <= 32'b00000000001000000000000110110011;
ROM[3490] <= 32'b00100100000100001010000011101111;
ROM[3491] <= 32'b11111111110000010000000100010011;
ROM[3492] <= 32'b00000000000000010010001110000011;
ROM[3493] <= 32'b00000000011100011010001000100011;
ROM[3494] <= 32'b00000000010000011010001110000011;
ROM[3495] <= 32'b00000000011100010010000000100011;
ROM[3496] <= 32'b00000000010000010000000100010011;
ROM[3497] <= 32'b00000000000100000000001110010011;
ROM[3498] <= 32'b00000000011100010010000000100011;
ROM[3499] <= 32'b00000000010000010000000100010011;
ROM[3500] <= 32'b11111111110000010000000100010011;
ROM[3501] <= 32'b00000000000000010010001110000011;
ROM[3502] <= 32'b11111111110000010000000100010011;
ROM[3503] <= 32'b00000000000000010010010000000011;
ROM[3504] <= 32'b00000000011101000010010010110011;
ROM[3505] <= 32'b00000000100000111010010100110011;
ROM[3506] <= 32'b00000000101001001000001110110011;
ROM[3507] <= 32'b00000000000100111000001110010011;
ROM[3508] <= 32'b00000000000100111111001110010011;
ROM[3509] <= 32'b00000000011100010010000000100011;
ROM[3510] <= 32'b00000000010000010000000100010011;
ROM[3511] <= 32'b11111111110000010000000100010011;
ROM[3512] <= 32'b00000000000000010010001110000011;
ROM[3513] <= 32'b00000000000000111000101001100011;
ROM[3514] <= 32'b00000000000000000100001110110111;
ROM[3515] <= 32'b11001001010000111000001110010011;
ROM[3516] <= 32'b00000000111000111000001110110011;
ROM[3517] <= 32'b00000000000000111000000011100111;
ROM[3518] <= 32'b00000000000000000000001110010011;
ROM[3519] <= 32'b00000000011100010010000000100011;
ROM[3520] <= 32'b00000000010000010000000100010011;
ROM[3521] <= 32'b11111111110000010000000100010011;
ROM[3522] <= 32'b00000000000000010010001110000011;
ROM[3523] <= 32'b00000000011100011010000000100011;
ROM[3524] <= 32'b00000000111000000000001110010011;
ROM[3525] <= 32'b00000000011100010010000000100011;
ROM[3526] <= 32'b00000000010000010000000100010011;
ROM[3527] <= 32'b00000000000000000011001110110111;
ROM[3528] <= 32'b01110110100000111000001110010011;
ROM[3529] <= 32'b00000000111000111000001110110011;
ROM[3530] <= 32'b00000000011100010010000000100011;
ROM[3531] <= 32'b00000000010000010000000100010011;
ROM[3532] <= 32'b00000000001100010010000000100011;
ROM[3533] <= 32'b00000000010000010000000100010011;
ROM[3534] <= 32'b00000000010000010010000000100011;
ROM[3535] <= 32'b00000000010000010000000100010011;
ROM[3536] <= 32'b00000000010100010010000000100011;
ROM[3537] <= 32'b00000000010000010000000100010011;
ROM[3538] <= 32'b00000000011000010010000000100011;
ROM[3539] <= 32'b00000000010000010000000100010011;
ROM[3540] <= 32'b00000001010000000000001110010011;
ROM[3541] <= 32'b00000000010000111000001110010011;
ROM[3542] <= 32'b01000000011100010000001110110011;
ROM[3543] <= 32'b00000000011100000000001000110011;
ROM[3544] <= 32'b00000000001000000000000110110011;
ROM[3545] <= 32'b01111101100100100101000011101111;
ROM[3546] <= 32'b00000101000000000000001110010011;
ROM[3547] <= 32'b00000000011100010010000000100011;
ROM[3548] <= 32'b00000000010000010000000100010011;
ROM[3549] <= 32'b00000000000000000011001110110111;
ROM[3550] <= 32'b01111100000000111000001110010011;
ROM[3551] <= 32'b00000000111000111000001110110011;
ROM[3552] <= 32'b00000000011100010010000000100011;
ROM[3553] <= 32'b00000000010000010000000100010011;
ROM[3554] <= 32'b00000000001100010010000000100011;
ROM[3555] <= 32'b00000000010000010000000100010011;
ROM[3556] <= 32'b00000000010000010010000000100011;
ROM[3557] <= 32'b00000000010000010000000100010011;
ROM[3558] <= 32'b00000000010100010010000000100011;
ROM[3559] <= 32'b00000000010000010000000100010011;
ROM[3560] <= 32'b00000000011000010010000000100011;
ROM[3561] <= 32'b00000000010000010000000100010011;
ROM[3562] <= 32'b00000001010000000000001110010011;
ROM[3563] <= 32'b00000000100000111000001110010011;
ROM[3564] <= 32'b01000000011100010000001110110011;
ROM[3565] <= 32'b00000000011100000000001000110011;
ROM[3566] <= 32'b00000000001000000000000110110011;
ROM[3567] <= 32'b00111111000000100110000011101111;
ROM[3568] <= 32'b00000111001000000000001110010011;
ROM[3569] <= 32'b00000000011100010010000000100011;
ROM[3570] <= 32'b00000000010000010000000100010011;
ROM[3571] <= 32'b00000000000000000100001110110111;
ROM[3572] <= 32'b10000001100000111000001110010011;
ROM[3573] <= 32'b00000000111000111000001110110011;
ROM[3574] <= 32'b00000000011100010010000000100011;
ROM[3575] <= 32'b00000000010000010000000100010011;
ROM[3576] <= 32'b00000000001100010010000000100011;
ROM[3577] <= 32'b00000000010000010000000100010011;
ROM[3578] <= 32'b00000000010000010010000000100011;
ROM[3579] <= 32'b00000000010000010000000100010011;
ROM[3580] <= 32'b00000000010100010010000000100011;
ROM[3581] <= 32'b00000000010000010000000100010011;
ROM[3582] <= 32'b00000000011000010010000000100011;
ROM[3583] <= 32'b00000000010000010000000100010011;
ROM[3584] <= 32'b00000001010000000000001110010011;
ROM[3585] <= 32'b00000000100000111000001110010011;
ROM[3586] <= 32'b01000000011100010000001110110011;
ROM[3587] <= 32'b00000000011100000000001000110011;
ROM[3588] <= 32'b00000000001000000000000110110011;
ROM[3589] <= 32'b00111001100000100110000011101111;
ROM[3590] <= 32'b00000110111100000000001110010011;
ROM[3591] <= 32'b00000000011100010010000000100011;
ROM[3592] <= 32'b00000000010000010000000100010011;
ROM[3593] <= 32'b00000000000000000100001110110111;
ROM[3594] <= 32'b10000111000000111000001110010011;
ROM[3595] <= 32'b00000000111000111000001110110011;
ROM[3596] <= 32'b00000000011100010010000000100011;
ROM[3597] <= 32'b00000000010000010000000100010011;
ROM[3598] <= 32'b00000000001100010010000000100011;
ROM[3599] <= 32'b00000000010000010000000100010011;
ROM[3600] <= 32'b00000000010000010010000000100011;
ROM[3601] <= 32'b00000000010000010000000100010011;
ROM[3602] <= 32'b00000000010100010010000000100011;
ROM[3603] <= 32'b00000000010000010000000100010011;
ROM[3604] <= 32'b00000000011000010010000000100011;
ROM[3605] <= 32'b00000000010000010000000100010011;
ROM[3606] <= 32'b00000001010000000000001110010011;
ROM[3607] <= 32'b00000000100000111000001110010011;
ROM[3608] <= 32'b01000000011100010000001110110011;
ROM[3609] <= 32'b00000000011100000000001000110011;
ROM[3610] <= 32'b00000000001000000000000110110011;
ROM[3611] <= 32'b00110100000000100110000011101111;
ROM[3612] <= 32'b00000110011100000000001110010011;
ROM[3613] <= 32'b00000000011100010010000000100011;
ROM[3614] <= 32'b00000000010000010000000100010011;
ROM[3615] <= 32'b00000000000000000100001110110111;
ROM[3616] <= 32'b10001100100000111000001110010011;
ROM[3617] <= 32'b00000000111000111000001110110011;
ROM[3618] <= 32'b00000000011100010010000000100011;
ROM[3619] <= 32'b00000000010000010000000100010011;
ROM[3620] <= 32'b00000000001100010010000000100011;
ROM[3621] <= 32'b00000000010000010000000100010011;
ROM[3622] <= 32'b00000000010000010010000000100011;
ROM[3623] <= 32'b00000000010000010000000100010011;
ROM[3624] <= 32'b00000000010100010010000000100011;
ROM[3625] <= 32'b00000000010000010000000100010011;
ROM[3626] <= 32'b00000000011000010010000000100011;
ROM[3627] <= 32'b00000000010000010000000100010011;
ROM[3628] <= 32'b00000001010000000000001110010011;
ROM[3629] <= 32'b00000000100000111000001110010011;
ROM[3630] <= 32'b01000000011100010000001110110011;
ROM[3631] <= 32'b00000000011100000000001000110011;
ROM[3632] <= 32'b00000000001000000000000110110011;
ROM[3633] <= 32'b00101110100000100110000011101111;
ROM[3634] <= 32'b00000111001000000000001110010011;
ROM[3635] <= 32'b00000000011100010010000000100011;
ROM[3636] <= 32'b00000000010000010000000100010011;
ROM[3637] <= 32'b00000000000000000100001110110111;
ROM[3638] <= 32'b10010010000000111000001110010011;
ROM[3639] <= 32'b00000000111000111000001110110011;
ROM[3640] <= 32'b00000000011100010010000000100011;
ROM[3641] <= 32'b00000000010000010000000100010011;
ROM[3642] <= 32'b00000000001100010010000000100011;
ROM[3643] <= 32'b00000000010000010000000100010011;
ROM[3644] <= 32'b00000000010000010010000000100011;
ROM[3645] <= 32'b00000000010000010000000100010011;
ROM[3646] <= 32'b00000000010100010010000000100011;
ROM[3647] <= 32'b00000000010000010000000100010011;
ROM[3648] <= 32'b00000000011000010010000000100011;
ROM[3649] <= 32'b00000000010000010000000100010011;
ROM[3650] <= 32'b00000001010000000000001110010011;
ROM[3651] <= 32'b00000000100000111000001110010011;
ROM[3652] <= 32'b01000000011100010000001110110011;
ROM[3653] <= 32'b00000000011100000000001000110011;
ROM[3654] <= 32'b00000000001000000000000110110011;
ROM[3655] <= 32'b00101001000000100110000011101111;
ROM[3656] <= 32'b00000110000100000000001110010011;
ROM[3657] <= 32'b00000000011100010010000000100011;
ROM[3658] <= 32'b00000000010000010000000100010011;
ROM[3659] <= 32'b00000000000000000100001110110111;
ROM[3660] <= 32'b10010111100000111000001110010011;
ROM[3661] <= 32'b00000000111000111000001110110011;
ROM[3662] <= 32'b00000000011100010010000000100011;
ROM[3663] <= 32'b00000000010000010000000100010011;
ROM[3664] <= 32'b00000000001100010010000000100011;
ROM[3665] <= 32'b00000000010000010000000100010011;
ROM[3666] <= 32'b00000000010000010010000000100011;
ROM[3667] <= 32'b00000000010000010000000100010011;
ROM[3668] <= 32'b00000000010100010010000000100011;
ROM[3669] <= 32'b00000000010000010000000100010011;
ROM[3670] <= 32'b00000000011000010010000000100011;
ROM[3671] <= 32'b00000000010000010000000100010011;
ROM[3672] <= 32'b00000001010000000000001110010011;
ROM[3673] <= 32'b00000000100000111000001110010011;
ROM[3674] <= 32'b01000000011100010000001110110011;
ROM[3675] <= 32'b00000000011100000000001000110011;
ROM[3676] <= 32'b00000000001000000000000110110011;
ROM[3677] <= 32'b00100011100000100110000011101111;
ROM[3678] <= 32'b00000110110100000000001110010011;
ROM[3679] <= 32'b00000000011100010010000000100011;
ROM[3680] <= 32'b00000000010000010000000100010011;
ROM[3681] <= 32'b00000000000000000100001110110111;
ROM[3682] <= 32'b10011101000000111000001110010011;
ROM[3683] <= 32'b00000000111000111000001110110011;
ROM[3684] <= 32'b00000000011100010010000000100011;
ROM[3685] <= 32'b00000000010000010000000100010011;
ROM[3686] <= 32'b00000000001100010010000000100011;
ROM[3687] <= 32'b00000000010000010000000100010011;
ROM[3688] <= 32'b00000000010000010010000000100011;
ROM[3689] <= 32'b00000000010000010000000100010011;
ROM[3690] <= 32'b00000000010100010010000000100011;
ROM[3691] <= 32'b00000000010000010000000100010011;
ROM[3692] <= 32'b00000000011000010010000000100011;
ROM[3693] <= 32'b00000000010000010000000100010011;
ROM[3694] <= 32'b00000001010000000000001110010011;
ROM[3695] <= 32'b00000000100000111000001110010011;
ROM[3696] <= 32'b01000000011100010000001110110011;
ROM[3697] <= 32'b00000000011100000000001000110011;
ROM[3698] <= 32'b00000000001000000000000110110011;
ROM[3699] <= 32'b00011110000000100110000011101111;
ROM[3700] <= 32'b00000010000000000000001110010011;
ROM[3701] <= 32'b00000000011100010010000000100011;
ROM[3702] <= 32'b00000000010000010000000100010011;
ROM[3703] <= 32'b00000000000000000100001110110111;
ROM[3704] <= 32'b10100010100000111000001110010011;
ROM[3705] <= 32'b00000000111000111000001110110011;
ROM[3706] <= 32'b00000000011100010010000000100011;
ROM[3707] <= 32'b00000000010000010000000100010011;
ROM[3708] <= 32'b00000000001100010010000000100011;
ROM[3709] <= 32'b00000000010000010000000100010011;
ROM[3710] <= 32'b00000000010000010010000000100011;
ROM[3711] <= 32'b00000000010000010000000100010011;
ROM[3712] <= 32'b00000000010100010010000000100011;
ROM[3713] <= 32'b00000000010000010000000100010011;
ROM[3714] <= 32'b00000000011000010010000000100011;
ROM[3715] <= 32'b00000000010000010000000100010011;
ROM[3716] <= 32'b00000001010000000000001110010011;
ROM[3717] <= 32'b00000000100000111000001110010011;
ROM[3718] <= 32'b01000000011100010000001110110011;
ROM[3719] <= 32'b00000000011100000000001000110011;
ROM[3720] <= 32'b00000000001000000000000110110011;
ROM[3721] <= 32'b00011000100000100110000011101111;
ROM[3722] <= 32'b00000110010100000000001110010011;
ROM[3723] <= 32'b00000000011100010010000000100011;
ROM[3724] <= 32'b00000000010000010000000100010011;
ROM[3725] <= 32'b00000000000000000100001110110111;
ROM[3726] <= 32'b10101000000000111000001110010011;
ROM[3727] <= 32'b00000000111000111000001110110011;
ROM[3728] <= 32'b00000000011100010010000000100011;
ROM[3729] <= 32'b00000000010000010000000100010011;
ROM[3730] <= 32'b00000000001100010010000000100011;
ROM[3731] <= 32'b00000000010000010000000100010011;
ROM[3732] <= 32'b00000000010000010010000000100011;
ROM[3733] <= 32'b00000000010000010000000100010011;
ROM[3734] <= 32'b00000000010100010010000000100011;
ROM[3735] <= 32'b00000000010000010000000100010011;
ROM[3736] <= 32'b00000000011000010010000000100011;
ROM[3737] <= 32'b00000000010000010000000100010011;
ROM[3738] <= 32'b00000001010000000000001110010011;
ROM[3739] <= 32'b00000000100000111000001110010011;
ROM[3740] <= 32'b01000000011100010000001110110011;
ROM[3741] <= 32'b00000000011100000000001000110011;
ROM[3742] <= 32'b00000000001000000000000110110011;
ROM[3743] <= 32'b00010011000000100110000011101111;
ROM[3744] <= 32'b00000110111000000000001110010011;
ROM[3745] <= 32'b00000000011100010010000000100011;
ROM[3746] <= 32'b00000000010000010000000100010011;
ROM[3747] <= 32'b00000000000000000100001110110111;
ROM[3748] <= 32'b10101101100000111000001110010011;
ROM[3749] <= 32'b00000000111000111000001110110011;
ROM[3750] <= 32'b00000000011100010010000000100011;
ROM[3751] <= 32'b00000000010000010000000100010011;
ROM[3752] <= 32'b00000000001100010010000000100011;
ROM[3753] <= 32'b00000000010000010000000100010011;
ROM[3754] <= 32'b00000000010000010010000000100011;
ROM[3755] <= 32'b00000000010000010000000100010011;
ROM[3756] <= 32'b00000000010100010010000000100011;
ROM[3757] <= 32'b00000000010000010000000100010011;
ROM[3758] <= 32'b00000000011000010010000000100011;
ROM[3759] <= 32'b00000000010000010000000100010011;
ROM[3760] <= 32'b00000001010000000000001110010011;
ROM[3761] <= 32'b00000000100000111000001110010011;
ROM[3762] <= 32'b01000000011100010000001110110011;
ROM[3763] <= 32'b00000000011100000000001000110011;
ROM[3764] <= 32'b00000000001000000000000110110011;
ROM[3765] <= 32'b00001101100000100110000011101111;
ROM[3766] <= 32'b00000110010000000000001110010011;
ROM[3767] <= 32'b00000000011100010010000000100011;
ROM[3768] <= 32'b00000000010000010000000100010011;
ROM[3769] <= 32'b00000000000000000100001110110111;
ROM[3770] <= 32'b10110011000000111000001110010011;
ROM[3771] <= 32'b00000000111000111000001110110011;
ROM[3772] <= 32'b00000000011100010010000000100011;
ROM[3773] <= 32'b00000000010000010000000100010011;
ROM[3774] <= 32'b00000000001100010010000000100011;
ROM[3775] <= 32'b00000000010000010000000100010011;
ROM[3776] <= 32'b00000000010000010010000000100011;
ROM[3777] <= 32'b00000000010000010000000100010011;
ROM[3778] <= 32'b00000000010100010010000000100011;
ROM[3779] <= 32'b00000000010000010000000100010011;
ROM[3780] <= 32'b00000000011000010010000000100011;
ROM[3781] <= 32'b00000000010000010000000100010011;
ROM[3782] <= 32'b00000001010000000000001110010011;
ROM[3783] <= 32'b00000000100000111000001110010011;
ROM[3784] <= 32'b01000000011100010000001110110011;
ROM[3785] <= 32'b00000000011100000000001000110011;
ROM[3786] <= 32'b00000000001000000000000110110011;
ROM[3787] <= 32'b00001000000000100110000011101111;
ROM[3788] <= 32'b00000110010100000000001110010011;
ROM[3789] <= 32'b00000000011100010010000000100011;
ROM[3790] <= 32'b00000000010000010000000100010011;
ROM[3791] <= 32'b00000000000000000100001110110111;
ROM[3792] <= 32'b10111000100000111000001110010011;
ROM[3793] <= 32'b00000000111000111000001110110011;
ROM[3794] <= 32'b00000000011100010010000000100011;
ROM[3795] <= 32'b00000000010000010000000100010011;
ROM[3796] <= 32'b00000000001100010010000000100011;
ROM[3797] <= 32'b00000000010000010000000100010011;
ROM[3798] <= 32'b00000000010000010010000000100011;
ROM[3799] <= 32'b00000000010000010000000100010011;
ROM[3800] <= 32'b00000000010100010010000000100011;
ROM[3801] <= 32'b00000000010000010000000100010011;
ROM[3802] <= 32'b00000000011000010010000000100011;
ROM[3803] <= 32'b00000000010000010000000100010011;
ROM[3804] <= 32'b00000001010000000000001110010011;
ROM[3805] <= 32'b00000000100000111000001110010011;
ROM[3806] <= 32'b01000000011100010000001110110011;
ROM[3807] <= 32'b00000000011100000000001000110011;
ROM[3808] <= 32'b00000000001000000000000110110011;
ROM[3809] <= 32'b00000010100000100110000011101111;
ROM[3810] <= 32'b00000110010000000000001110010011;
ROM[3811] <= 32'b00000000011100010010000000100011;
ROM[3812] <= 32'b00000000010000010000000100010011;
ROM[3813] <= 32'b00000000000000000100001110110111;
ROM[3814] <= 32'b10111110000000111000001110010011;
ROM[3815] <= 32'b00000000111000111000001110110011;
ROM[3816] <= 32'b00000000011100010010000000100011;
ROM[3817] <= 32'b00000000010000010000000100010011;
ROM[3818] <= 32'b00000000001100010010000000100011;
ROM[3819] <= 32'b00000000010000010000000100010011;
ROM[3820] <= 32'b00000000010000010010000000100011;
ROM[3821] <= 32'b00000000010000010000000100010011;
ROM[3822] <= 32'b00000000010100010010000000100011;
ROM[3823] <= 32'b00000000010000010000000100010011;
ROM[3824] <= 32'b00000000011000010010000000100011;
ROM[3825] <= 32'b00000000010000010000000100010011;
ROM[3826] <= 32'b00000001010000000000001110010011;
ROM[3827] <= 32'b00000000100000111000001110010011;
ROM[3828] <= 32'b01000000011100010000001110110011;
ROM[3829] <= 32'b00000000011100000000001000110011;
ROM[3830] <= 32'b00000000001000000000000110110011;
ROM[3831] <= 32'b01111101000100100101000011101111;
ROM[3832] <= 32'b00000010111000000000001110010011;
ROM[3833] <= 32'b00000000011100010010000000100011;
ROM[3834] <= 32'b00000000010000010000000100010011;
ROM[3835] <= 32'b00000000000000000100001110110111;
ROM[3836] <= 32'b11000011100000111000001110010011;
ROM[3837] <= 32'b00000000111000111000001110110011;
ROM[3838] <= 32'b00000000011100010010000000100011;
ROM[3839] <= 32'b00000000010000010000000100010011;
ROM[3840] <= 32'b00000000001100010010000000100011;
ROM[3841] <= 32'b00000000010000010000000100010011;
ROM[3842] <= 32'b00000000010000010010000000100011;
ROM[3843] <= 32'b00000000010000010000000100010011;
ROM[3844] <= 32'b00000000010100010010000000100011;
ROM[3845] <= 32'b00000000010000010000000100010011;
ROM[3846] <= 32'b00000000011000010010000000100011;
ROM[3847] <= 32'b00000000010000010000000100010011;
ROM[3848] <= 32'b00000001010000000000001110010011;
ROM[3849] <= 32'b00000000100000111000001110010011;
ROM[3850] <= 32'b01000000011100010000001110110011;
ROM[3851] <= 32'b00000000011100000000001000110011;
ROM[3852] <= 32'b00000000001000000000000110110011;
ROM[3853] <= 32'b01110111100100100101000011101111;
ROM[3854] <= 32'b00000000000000000100001110110111;
ROM[3855] <= 32'b11001000010000111000001110010011;
ROM[3856] <= 32'b00000000111000111000001110110011;
ROM[3857] <= 32'b00000000011100010010000000100011;
ROM[3858] <= 32'b00000000010000010000000100010011;
ROM[3859] <= 32'b00000000001100010010000000100011;
ROM[3860] <= 32'b00000000010000010000000100010011;
ROM[3861] <= 32'b00000000010000010010000000100011;
ROM[3862] <= 32'b00000000010000010000000100010011;
ROM[3863] <= 32'b00000000010100010010000000100011;
ROM[3864] <= 32'b00000000010000010000000100010011;
ROM[3865] <= 32'b00000000011000010010000000100011;
ROM[3866] <= 32'b00000000010000010000000100010011;
ROM[3867] <= 32'b00000001010000000000001110010011;
ROM[3868] <= 32'b00000000010000111000001110010011;
ROM[3869] <= 32'b01000000011100010000001110110011;
ROM[3870] <= 32'b00000000011100000000001000110011;
ROM[3871] <= 32'b00000000001000000000000110110011;
ROM[3872] <= 32'b00101110100000010011000011101111;
ROM[3873] <= 32'b11111111110000010000000100010011;
ROM[3874] <= 32'b00000000000000010010001110000011;
ROM[3875] <= 32'b00000000011101100010000000100011;
ROM[3876] <= 32'b00000101110000000000000011101111;
ROM[3877] <= 32'b00000000000000000100001110110111;
ROM[3878] <= 32'b11001110000000111000001110010011;
ROM[3879] <= 32'b00000000111000111000001110110011;
ROM[3880] <= 32'b00000000011100010010000000100011;
ROM[3881] <= 32'b00000000010000010000000100010011;
ROM[3882] <= 32'b00000000001100010010000000100011;
ROM[3883] <= 32'b00000000010000010000000100010011;
ROM[3884] <= 32'b00000000010000010010000000100011;
ROM[3885] <= 32'b00000000010000010000000100010011;
ROM[3886] <= 32'b00000000010100010010000000100011;
ROM[3887] <= 32'b00000000010000010000000100010011;
ROM[3888] <= 32'b00000000011000010010000000100011;
ROM[3889] <= 32'b00000000010000010000000100010011;
ROM[3890] <= 32'b00000001010000000000001110010011;
ROM[3891] <= 32'b00000000000000111000001110010011;
ROM[3892] <= 32'b01000000011100010000001110110011;
ROM[3893] <= 32'b00000000011100000000001000110011;
ROM[3894] <= 32'b00000000001000000000000110110011;
ROM[3895] <= 32'b11001111000011111100000011101111;
ROM[3896] <= 32'b11111111110000010000000100010011;
ROM[3897] <= 32'b00000000000000010010001110000011;
ROM[3898] <= 32'b00000000011101100010000000100011;
ROM[3899] <= 32'b10100001010111111110000011101111;
ROM[3900] <= 32'b00000000000000000000001110010011;
ROM[3901] <= 32'b00000000011100010010000000100011;
ROM[3902] <= 32'b00000000010000010000000100010011;
ROM[3903] <= 32'b00000001010000000000001110010011;
ROM[3904] <= 32'b01000000011100011000001110110011;
ROM[3905] <= 32'b00000000000000111010000010000011;
ROM[3906] <= 32'b11111111110000010000000100010011;
ROM[3907] <= 32'b00000000000000010010001110000011;
ROM[3908] <= 32'b00000000011100100010000000100011;
ROM[3909] <= 32'b00000000010000100000000100010011;
ROM[3910] <= 32'b00000001010000000000001110010011;
ROM[3911] <= 32'b01000000011100011000001110110011;
ROM[3912] <= 32'b00000000010000111010000110000011;
ROM[3913] <= 32'b00000000100000111010001000000011;
ROM[3914] <= 32'b00000000110000111010001010000011;
ROM[3915] <= 32'b00000001000000111010001100000011;
ROM[3916] <= 32'b00000000000000001000000011100111;
ROM[3917] <= 32'b00000000000000100010001110000011;
ROM[3918] <= 32'b00000000011100010010000000100011;
ROM[3919] <= 32'b00000000010000010000000100010011;
ROM[3920] <= 32'b00000100000100000000001110010011;
ROM[3921] <= 32'b00000000011100010010000000100011;
ROM[3922] <= 32'b00000000010000010000000100010011;
ROM[3923] <= 32'b11111111110000010000000100010011;
ROM[3924] <= 32'b00000000000000010010001110000011;
ROM[3925] <= 32'b11111111110000010000000100010011;
ROM[3926] <= 32'b00000000000000010010010000000011;
ROM[3927] <= 32'b00000000011101000010010010110011;
ROM[3928] <= 32'b00000000100000111010010100110011;
ROM[3929] <= 32'b00000000101001001000001110110011;
ROM[3930] <= 32'b00000000000100111000001110010011;
ROM[3931] <= 32'b00000000000100111111001110010011;
ROM[3932] <= 32'b00000000011100010010000000100011;
ROM[3933] <= 32'b00000000010000010000000100010011;
ROM[3934] <= 32'b11111111110000010000000100010011;
ROM[3935] <= 32'b00000000000000010010001110000011;
ROM[3936] <= 32'b00000000000000111000101001100011;
ROM[3937] <= 32'b00000000000000000101001110110111;
ROM[3938] <= 32'b11100101100000111000001110010011;
ROM[3939] <= 32'b00000000111000111000001110110011;
ROM[3940] <= 32'b00000000000000111000000011100111;
ROM[3941] <= 32'b00000000000000100010001110000011;
ROM[3942] <= 32'b00000000011100010010000000100011;
ROM[3943] <= 32'b00000000010000010000000100010011;
ROM[3944] <= 32'b00000100001000000000001110010011;
ROM[3945] <= 32'b00000000011100010010000000100011;
ROM[3946] <= 32'b00000000010000010000000100010011;
ROM[3947] <= 32'b11111111110000010000000100010011;
ROM[3948] <= 32'b00000000000000010010001110000011;
ROM[3949] <= 32'b11111111110000010000000100010011;
ROM[3950] <= 32'b00000000000000010010010000000011;
ROM[3951] <= 32'b00000000011101000010010010110011;
ROM[3952] <= 32'b00000000100000111010010100110011;
ROM[3953] <= 32'b00000000101001001000001110110011;
ROM[3954] <= 32'b00000000000100111000001110010011;
ROM[3955] <= 32'b00000000000100111111001110010011;
ROM[3956] <= 32'b00000000011100010010000000100011;
ROM[3957] <= 32'b00000000010000010000000100010011;
ROM[3958] <= 32'b11111111110000010000000100010011;
ROM[3959] <= 32'b00000000000000010010001110000011;
ROM[3960] <= 32'b00000000000000111000101001100011;
ROM[3961] <= 32'b00000000000000000101001110110111;
ROM[3962] <= 32'b11100001000000111000001110010011;
ROM[3963] <= 32'b00000000111000111000001110110011;
ROM[3964] <= 32'b00000000000000111000000011100111;
ROM[3965] <= 32'b00000000000000100010001110000011;
ROM[3966] <= 32'b00000000011100010010000000100011;
ROM[3967] <= 32'b00000000010000010000000100010011;
ROM[3968] <= 32'b00000100001100000000001110010011;
ROM[3969] <= 32'b00000000011100010010000000100011;
ROM[3970] <= 32'b00000000010000010000000100010011;
ROM[3971] <= 32'b11111111110000010000000100010011;
ROM[3972] <= 32'b00000000000000010010001110000011;
ROM[3973] <= 32'b11111111110000010000000100010011;
ROM[3974] <= 32'b00000000000000010010010000000011;
ROM[3975] <= 32'b00000000011101000010010010110011;
ROM[3976] <= 32'b00000000100000111010010100110011;
ROM[3977] <= 32'b00000000101001001000001110110011;
ROM[3978] <= 32'b00000000000100111000001110010011;
ROM[3979] <= 32'b00000000000100111111001110010011;
ROM[3980] <= 32'b00000000011100010010000000100011;
ROM[3981] <= 32'b00000000010000010000000100010011;
ROM[3982] <= 32'b11111111110000010000000100010011;
ROM[3983] <= 32'b00000000000000010010001110000011;
ROM[3984] <= 32'b00000000000000111000101001100011;
ROM[3985] <= 32'b00000000000000000101001110110111;
ROM[3986] <= 32'b11011100100000111000001110010011;
ROM[3987] <= 32'b00000000111000111000001110110011;
ROM[3988] <= 32'b00000000000000111000000011100111;
ROM[3989] <= 32'b00000000000000100010001110000011;
ROM[3990] <= 32'b00000000011100010010000000100011;
ROM[3991] <= 32'b00000000010000010000000100010011;
ROM[3992] <= 32'b00000100010000000000001110010011;
ROM[3993] <= 32'b00000000011100010010000000100011;
ROM[3994] <= 32'b00000000010000010000000100010011;
ROM[3995] <= 32'b11111111110000010000000100010011;
ROM[3996] <= 32'b00000000000000010010001110000011;
ROM[3997] <= 32'b11111111110000010000000100010011;
ROM[3998] <= 32'b00000000000000010010010000000011;
ROM[3999] <= 32'b00000000011101000010010010110011;
ROM[4000] <= 32'b00000000100000111010010100110011;
ROM[4001] <= 32'b00000000101001001000001110110011;
ROM[4002] <= 32'b00000000000100111000001110010011;
ROM[4003] <= 32'b00000000000100111111001110010011;
ROM[4004] <= 32'b00000000011100010010000000100011;
ROM[4005] <= 32'b00000000010000010000000100010011;
ROM[4006] <= 32'b11111111110000010000000100010011;
ROM[4007] <= 32'b00000000000000010010001110000011;
ROM[4008] <= 32'b00000000000000111000101001100011;
ROM[4009] <= 32'b00000000000000000101001110110111;
ROM[4010] <= 32'b11011000000000111000001110010011;
ROM[4011] <= 32'b00000000111000111000001110110011;
ROM[4012] <= 32'b00000000000000111000000011100111;
ROM[4013] <= 32'b00000000000000100010001110000011;
ROM[4014] <= 32'b00000000011100010010000000100011;
ROM[4015] <= 32'b00000000010000010000000100010011;
ROM[4016] <= 32'b00000100010100000000001110010011;
ROM[4017] <= 32'b00000000011100010010000000100011;
ROM[4018] <= 32'b00000000010000010000000100010011;
ROM[4019] <= 32'b11111111110000010000000100010011;
ROM[4020] <= 32'b00000000000000010010001110000011;
ROM[4021] <= 32'b11111111110000010000000100010011;
ROM[4022] <= 32'b00000000000000010010010000000011;
ROM[4023] <= 32'b00000000011101000010010010110011;
ROM[4024] <= 32'b00000000100000111010010100110011;
ROM[4025] <= 32'b00000000101001001000001110110011;
ROM[4026] <= 32'b00000000000100111000001110010011;
ROM[4027] <= 32'b00000000000100111111001110010011;
ROM[4028] <= 32'b00000000011100010010000000100011;
ROM[4029] <= 32'b00000000010000010000000100010011;
ROM[4030] <= 32'b11111111110000010000000100010011;
ROM[4031] <= 32'b00000000000000010010001110000011;
ROM[4032] <= 32'b00000000000000111000101001100011;
ROM[4033] <= 32'b00000000000000000101001110110111;
ROM[4034] <= 32'b11010011100000111000001110010011;
ROM[4035] <= 32'b00000000111000111000001110110011;
ROM[4036] <= 32'b00000000000000111000000011100111;
ROM[4037] <= 32'b00000000000000100010001110000011;
ROM[4038] <= 32'b00000000011100010010000000100011;
ROM[4039] <= 32'b00000000010000010000000100010011;
ROM[4040] <= 32'b00000100011000000000001110010011;
ROM[4041] <= 32'b00000000011100010010000000100011;
ROM[4042] <= 32'b00000000010000010000000100010011;
ROM[4043] <= 32'b11111111110000010000000100010011;
ROM[4044] <= 32'b00000000000000010010001110000011;
ROM[4045] <= 32'b11111111110000010000000100010011;
ROM[4046] <= 32'b00000000000000010010010000000011;
ROM[4047] <= 32'b00000000011101000010010010110011;
ROM[4048] <= 32'b00000000100000111010010100110011;
ROM[4049] <= 32'b00000000101001001000001110110011;
ROM[4050] <= 32'b00000000000100111000001110010011;
ROM[4051] <= 32'b00000000000100111111001110010011;
ROM[4052] <= 32'b00000000011100010010000000100011;
ROM[4053] <= 32'b00000000010000010000000100010011;
ROM[4054] <= 32'b11111111110000010000000100010011;
ROM[4055] <= 32'b00000000000000010010001110000011;
ROM[4056] <= 32'b00000000000000111000101001100011;
ROM[4057] <= 32'b00000000000000000101001110110111;
ROM[4058] <= 32'b11001111000000111000001110010011;
ROM[4059] <= 32'b00000000111000111000001110110011;
ROM[4060] <= 32'b00000000000000111000000011100111;
ROM[4061] <= 32'b00000000000000100010001110000011;
ROM[4062] <= 32'b00000000011100010010000000100011;
ROM[4063] <= 32'b00000000010000010000000100010011;
ROM[4064] <= 32'b00000100011100000000001110010011;
ROM[4065] <= 32'b00000000011100010010000000100011;
ROM[4066] <= 32'b00000000010000010000000100010011;
ROM[4067] <= 32'b11111111110000010000000100010011;
ROM[4068] <= 32'b00000000000000010010001110000011;
ROM[4069] <= 32'b11111111110000010000000100010011;
ROM[4070] <= 32'b00000000000000010010010000000011;
ROM[4071] <= 32'b00000000011101000010010010110011;
ROM[4072] <= 32'b00000000100000111010010100110011;
ROM[4073] <= 32'b00000000101001001000001110110011;
ROM[4074] <= 32'b00000000000100111000001110010011;
ROM[4075] <= 32'b00000000000100111111001110010011;
ROM[4076] <= 32'b00000000011100010010000000100011;
ROM[4077] <= 32'b00000000010000010000000100010011;
ROM[4078] <= 32'b11111111110000010000000100010011;
ROM[4079] <= 32'b00000000000000010010001110000011;
ROM[4080] <= 32'b00000000000000111000101001100011;
ROM[4081] <= 32'b00000000000000000101001110110111;
ROM[4082] <= 32'b11001010100000111000001110010011;
ROM[4083] <= 32'b00000000111000111000001110110011;
ROM[4084] <= 32'b00000000000000111000000011100111;
ROM[4085] <= 32'b00000000000000100010001110000011;
ROM[4086] <= 32'b00000000011100010010000000100011;
ROM[4087] <= 32'b00000000010000010000000100010011;
ROM[4088] <= 32'b00000100100000000000001110010011;
ROM[4089] <= 32'b00000000011100010010000000100011;
ROM[4090] <= 32'b00000000010000010000000100010011;
ROM[4091] <= 32'b11111111110000010000000100010011;
ROM[4092] <= 32'b00000000000000010010001110000011;
ROM[4093] <= 32'b11111111110000010000000100010011;
ROM[4094] <= 32'b00000000000000010010010000000011;
ROM[4095] <= 32'b00000000011101000010010010110011;
ROM[4096] <= 32'b00000000100000111010010100110011;
ROM[4097] <= 32'b00000000101001001000001110110011;
ROM[4098] <= 32'b00000000000100111000001110010011;
ROM[4099] <= 32'b00000000000100111111001110010011;
ROM[4100] <= 32'b00000000011100010010000000100011;
ROM[4101] <= 32'b00000000010000010000000100010011;
ROM[4102] <= 32'b11111111110000010000000100010011;
ROM[4103] <= 32'b00000000000000010010001110000011;
ROM[4104] <= 32'b00000000000000111000101001100011;
ROM[4105] <= 32'b00000000000000000101001110110111;
ROM[4106] <= 32'b11000110000000111000001110010011;
ROM[4107] <= 32'b00000000111000111000001110110011;
ROM[4108] <= 32'b00000000000000111000000011100111;
ROM[4109] <= 32'b00000000000000100010001110000011;
ROM[4110] <= 32'b00000000011100010010000000100011;
ROM[4111] <= 32'b00000000010000010000000100010011;
ROM[4112] <= 32'b00000100100100000000001110010011;
ROM[4113] <= 32'b00000000011100010010000000100011;
ROM[4114] <= 32'b00000000010000010000000100010011;
ROM[4115] <= 32'b11111111110000010000000100010011;
ROM[4116] <= 32'b00000000000000010010001110000011;
ROM[4117] <= 32'b11111111110000010000000100010011;
ROM[4118] <= 32'b00000000000000010010010000000011;
ROM[4119] <= 32'b00000000011101000010010010110011;
ROM[4120] <= 32'b00000000100000111010010100110011;
ROM[4121] <= 32'b00000000101001001000001110110011;
ROM[4122] <= 32'b00000000000100111000001110010011;
ROM[4123] <= 32'b00000000000100111111001110010011;
ROM[4124] <= 32'b00000000011100010010000000100011;
ROM[4125] <= 32'b00000000010000010000000100010011;
ROM[4126] <= 32'b11111111110000010000000100010011;
ROM[4127] <= 32'b00000000000000010010001110000011;
ROM[4128] <= 32'b00000000000000111000101001100011;
ROM[4129] <= 32'b00000000000000000101001110110111;
ROM[4130] <= 32'b11000001100000111000001110010011;
ROM[4131] <= 32'b00000000111000111000001110110011;
ROM[4132] <= 32'b00000000000000111000000011100111;
ROM[4133] <= 32'b00000000000000100010001110000011;
ROM[4134] <= 32'b00000000011100010010000000100011;
ROM[4135] <= 32'b00000000010000010000000100010011;
ROM[4136] <= 32'b00000100101000000000001110010011;
ROM[4137] <= 32'b00000000011100010010000000100011;
ROM[4138] <= 32'b00000000010000010000000100010011;
ROM[4139] <= 32'b11111111110000010000000100010011;
ROM[4140] <= 32'b00000000000000010010001110000011;
ROM[4141] <= 32'b11111111110000010000000100010011;
ROM[4142] <= 32'b00000000000000010010010000000011;
ROM[4143] <= 32'b00000000011101000010010010110011;
ROM[4144] <= 32'b00000000100000111010010100110011;
ROM[4145] <= 32'b00000000101001001000001110110011;
ROM[4146] <= 32'b00000000000100111000001110010011;
ROM[4147] <= 32'b00000000000100111111001110010011;
ROM[4148] <= 32'b00000000011100010010000000100011;
ROM[4149] <= 32'b00000000010000010000000100010011;
ROM[4150] <= 32'b11111111110000010000000100010011;
ROM[4151] <= 32'b00000000000000010010001110000011;
ROM[4152] <= 32'b00000000000000111000101001100011;
ROM[4153] <= 32'b00000000000000000101001110110111;
ROM[4154] <= 32'b10111101000000111000001110010011;
ROM[4155] <= 32'b00000000111000111000001110110011;
ROM[4156] <= 32'b00000000000000111000000011100111;
ROM[4157] <= 32'b00000000000000100010001110000011;
ROM[4158] <= 32'b00000000011100010010000000100011;
ROM[4159] <= 32'b00000000010000010000000100010011;
ROM[4160] <= 32'b00000100101100000000001110010011;
ROM[4161] <= 32'b00000000011100010010000000100011;
ROM[4162] <= 32'b00000000010000010000000100010011;
ROM[4163] <= 32'b11111111110000010000000100010011;
ROM[4164] <= 32'b00000000000000010010001110000011;
ROM[4165] <= 32'b11111111110000010000000100010011;
ROM[4166] <= 32'b00000000000000010010010000000011;
ROM[4167] <= 32'b00000000011101000010010010110011;
ROM[4168] <= 32'b00000000100000111010010100110011;
ROM[4169] <= 32'b00000000101001001000001110110011;
ROM[4170] <= 32'b00000000000100111000001110010011;
ROM[4171] <= 32'b00000000000100111111001110010011;
ROM[4172] <= 32'b00000000011100010010000000100011;
ROM[4173] <= 32'b00000000010000010000000100010011;
ROM[4174] <= 32'b11111111110000010000000100010011;
ROM[4175] <= 32'b00000000000000010010001110000011;
ROM[4176] <= 32'b00000000000000111000101001100011;
ROM[4177] <= 32'b00000000000000000101001110110111;
ROM[4178] <= 32'b10111000100000111000001110010011;
ROM[4179] <= 32'b00000000111000111000001110110011;
ROM[4180] <= 32'b00000000000000111000000011100111;
ROM[4181] <= 32'b00000000000000100010001110000011;
ROM[4182] <= 32'b00000000011100010010000000100011;
ROM[4183] <= 32'b00000000010000010000000100010011;
ROM[4184] <= 32'b00000100110000000000001110010011;
ROM[4185] <= 32'b00000000011100010010000000100011;
ROM[4186] <= 32'b00000000010000010000000100010011;
ROM[4187] <= 32'b11111111110000010000000100010011;
ROM[4188] <= 32'b00000000000000010010001110000011;
ROM[4189] <= 32'b11111111110000010000000100010011;
ROM[4190] <= 32'b00000000000000010010010000000011;
ROM[4191] <= 32'b00000000011101000010010010110011;
ROM[4192] <= 32'b00000000100000111010010100110011;
ROM[4193] <= 32'b00000000101001001000001110110011;
ROM[4194] <= 32'b00000000000100111000001110010011;
ROM[4195] <= 32'b00000000000100111111001110010011;
ROM[4196] <= 32'b00000000011100010010000000100011;
ROM[4197] <= 32'b00000000010000010000000100010011;
ROM[4198] <= 32'b11111111110000010000000100010011;
ROM[4199] <= 32'b00000000000000010010001110000011;
ROM[4200] <= 32'b00000000000000111000101001100011;
ROM[4201] <= 32'b00000000000000000101001110110111;
ROM[4202] <= 32'b10110100000000111000001110010011;
ROM[4203] <= 32'b00000000111000111000001110110011;
ROM[4204] <= 32'b00000000000000111000000011100111;
ROM[4205] <= 32'b00000000000000100010001110000011;
ROM[4206] <= 32'b00000000011100010010000000100011;
ROM[4207] <= 32'b00000000010000010000000100010011;
ROM[4208] <= 32'b00000100110100000000001110010011;
ROM[4209] <= 32'b00000000011100010010000000100011;
ROM[4210] <= 32'b00000000010000010000000100010011;
ROM[4211] <= 32'b11111111110000010000000100010011;
ROM[4212] <= 32'b00000000000000010010001110000011;
ROM[4213] <= 32'b11111111110000010000000100010011;
ROM[4214] <= 32'b00000000000000010010010000000011;
ROM[4215] <= 32'b00000000011101000010010010110011;
ROM[4216] <= 32'b00000000100000111010010100110011;
ROM[4217] <= 32'b00000000101001001000001110110011;
ROM[4218] <= 32'b00000000000100111000001110010011;
ROM[4219] <= 32'b00000000000100111111001110010011;
ROM[4220] <= 32'b00000000011100010010000000100011;
ROM[4221] <= 32'b00000000010000010000000100010011;
ROM[4222] <= 32'b11111111110000010000000100010011;
ROM[4223] <= 32'b00000000000000010010001110000011;
ROM[4224] <= 32'b00000000000000111000101001100011;
ROM[4225] <= 32'b00000000000000000101001110110111;
ROM[4226] <= 32'b10101111100000111000001110010011;
ROM[4227] <= 32'b00000000111000111000001110110011;
ROM[4228] <= 32'b00000000000000111000000011100111;
ROM[4229] <= 32'b00000000000000100010001110000011;
ROM[4230] <= 32'b00000000011100010010000000100011;
ROM[4231] <= 32'b00000000010000010000000100010011;
ROM[4232] <= 32'b00000100111000000000001110010011;
ROM[4233] <= 32'b00000000011100010010000000100011;
ROM[4234] <= 32'b00000000010000010000000100010011;
ROM[4235] <= 32'b11111111110000010000000100010011;
ROM[4236] <= 32'b00000000000000010010001110000011;
ROM[4237] <= 32'b11111111110000010000000100010011;
ROM[4238] <= 32'b00000000000000010010010000000011;
ROM[4239] <= 32'b00000000011101000010010010110011;
ROM[4240] <= 32'b00000000100000111010010100110011;
ROM[4241] <= 32'b00000000101001001000001110110011;
ROM[4242] <= 32'b00000000000100111000001110010011;
ROM[4243] <= 32'b00000000000100111111001110010011;
ROM[4244] <= 32'b00000000011100010010000000100011;
ROM[4245] <= 32'b00000000010000010000000100010011;
ROM[4246] <= 32'b11111111110000010000000100010011;
ROM[4247] <= 32'b00000000000000010010001110000011;
ROM[4248] <= 32'b00000000000000111000101001100011;
ROM[4249] <= 32'b00000000000000000101001110110111;
ROM[4250] <= 32'b10101011000000111000001110010011;
ROM[4251] <= 32'b00000000111000111000001110110011;
ROM[4252] <= 32'b00000000000000111000000011100111;
ROM[4253] <= 32'b00000000000000100010001110000011;
ROM[4254] <= 32'b00000000011100010010000000100011;
ROM[4255] <= 32'b00000000010000010000000100010011;
ROM[4256] <= 32'b00000100111100000000001110010011;
ROM[4257] <= 32'b00000000011100010010000000100011;
ROM[4258] <= 32'b00000000010000010000000100010011;
ROM[4259] <= 32'b11111111110000010000000100010011;
ROM[4260] <= 32'b00000000000000010010001110000011;
ROM[4261] <= 32'b11111111110000010000000100010011;
ROM[4262] <= 32'b00000000000000010010010000000011;
ROM[4263] <= 32'b00000000011101000010010010110011;
ROM[4264] <= 32'b00000000100000111010010100110011;
ROM[4265] <= 32'b00000000101001001000001110110011;
ROM[4266] <= 32'b00000000000100111000001110010011;
ROM[4267] <= 32'b00000000000100111111001110010011;
ROM[4268] <= 32'b00000000011100010010000000100011;
ROM[4269] <= 32'b00000000010000010000000100010011;
ROM[4270] <= 32'b11111111110000010000000100010011;
ROM[4271] <= 32'b00000000000000010010001110000011;
ROM[4272] <= 32'b00000000000000111000101001100011;
ROM[4273] <= 32'b00000000000000000101001110110111;
ROM[4274] <= 32'b10100110100000111000001110010011;
ROM[4275] <= 32'b00000000111000111000001110110011;
ROM[4276] <= 32'b00000000000000111000000011100111;
ROM[4277] <= 32'b00000000000000100010001110000011;
ROM[4278] <= 32'b00000000011100010010000000100011;
ROM[4279] <= 32'b00000000010000010000000100010011;
ROM[4280] <= 32'b00000101000000000000001110010011;
ROM[4281] <= 32'b00000000011100010010000000100011;
ROM[4282] <= 32'b00000000010000010000000100010011;
ROM[4283] <= 32'b11111111110000010000000100010011;
ROM[4284] <= 32'b00000000000000010010001110000011;
ROM[4285] <= 32'b11111111110000010000000100010011;
ROM[4286] <= 32'b00000000000000010010010000000011;
ROM[4287] <= 32'b00000000011101000010010010110011;
ROM[4288] <= 32'b00000000100000111010010100110011;
ROM[4289] <= 32'b00000000101001001000001110110011;
ROM[4290] <= 32'b00000000000100111000001110010011;
ROM[4291] <= 32'b00000000000100111111001110010011;
ROM[4292] <= 32'b00000000011100010010000000100011;
ROM[4293] <= 32'b00000000010000010000000100010011;
ROM[4294] <= 32'b11111111110000010000000100010011;
ROM[4295] <= 32'b00000000000000010010001110000011;
ROM[4296] <= 32'b00000000000000111000101001100011;
ROM[4297] <= 32'b00000000000000000101001110110111;
ROM[4298] <= 32'b10100010000000111000001110010011;
ROM[4299] <= 32'b00000000111000111000001110110011;
ROM[4300] <= 32'b00000000000000111000000011100111;
ROM[4301] <= 32'b00000000000000100010001110000011;
ROM[4302] <= 32'b00000000011100010010000000100011;
ROM[4303] <= 32'b00000000010000010000000100010011;
ROM[4304] <= 32'b00000101000100000000001110010011;
ROM[4305] <= 32'b00000000011100010010000000100011;
ROM[4306] <= 32'b00000000010000010000000100010011;
ROM[4307] <= 32'b11111111110000010000000100010011;
ROM[4308] <= 32'b00000000000000010010001110000011;
ROM[4309] <= 32'b11111111110000010000000100010011;
ROM[4310] <= 32'b00000000000000010010010000000011;
ROM[4311] <= 32'b00000000011101000010010010110011;
ROM[4312] <= 32'b00000000100000111010010100110011;
ROM[4313] <= 32'b00000000101001001000001110110011;
ROM[4314] <= 32'b00000000000100111000001110010011;
ROM[4315] <= 32'b00000000000100111111001110010011;
ROM[4316] <= 32'b00000000011100010010000000100011;
ROM[4317] <= 32'b00000000010000010000000100010011;
ROM[4318] <= 32'b11111111110000010000000100010011;
ROM[4319] <= 32'b00000000000000010010001110000011;
ROM[4320] <= 32'b00000000000000111000101001100011;
ROM[4321] <= 32'b00000000000000000101001110110111;
ROM[4322] <= 32'b10011101100000111000001110010011;
ROM[4323] <= 32'b00000000111000111000001110110011;
ROM[4324] <= 32'b00000000000000111000000011100111;
ROM[4325] <= 32'b00000000000000100010001110000011;
ROM[4326] <= 32'b00000000011100010010000000100011;
ROM[4327] <= 32'b00000000010000010000000100010011;
ROM[4328] <= 32'b00000101001000000000001110010011;
ROM[4329] <= 32'b00000000011100010010000000100011;
ROM[4330] <= 32'b00000000010000010000000100010011;
ROM[4331] <= 32'b11111111110000010000000100010011;
ROM[4332] <= 32'b00000000000000010010001110000011;
ROM[4333] <= 32'b11111111110000010000000100010011;
ROM[4334] <= 32'b00000000000000010010010000000011;
ROM[4335] <= 32'b00000000011101000010010010110011;
ROM[4336] <= 32'b00000000100000111010010100110011;
ROM[4337] <= 32'b00000000101001001000001110110011;
ROM[4338] <= 32'b00000000000100111000001110010011;
ROM[4339] <= 32'b00000000000100111111001110010011;
ROM[4340] <= 32'b00000000011100010010000000100011;
ROM[4341] <= 32'b00000000010000010000000100010011;
ROM[4342] <= 32'b11111111110000010000000100010011;
ROM[4343] <= 32'b00000000000000010010001110000011;
ROM[4344] <= 32'b00000000000000111000101001100011;
ROM[4345] <= 32'b00000000000000000101001110110111;
ROM[4346] <= 32'b10011001000000111000001110010011;
ROM[4347] <= 32'b00000000111000111000001110110011;
ROM[4348] <= 32'b00000000000000111000000011100111;
ROM[4349] <= 32'b00000000000000100010001110000011;
ROM[4350] <= 32'b00000000011100010010000000100011;
ROM[4351] <= 32'b00000000010000010000000100010011;
ROM[4352] <= 32'b00000101001100000000001110010011;
ROM[4353] <= 32'b00000000011100010010000000100011;
ROM[4354] <= 32'b00000000010000010000000100010011;
ROM[4355] <= 32'b11111111110000010000000100010011;
ROM[4356] <= 32'b00000000000000010010001110000011;
ROM[4357] <= 32'b11111111110000010000000100010011;
ROM[4358] <= 32'b00000000000000010010010000000011;
ROM[4359] <= 32'b00000000011101000010010010110011;
ROM[4360] <= 32'b00000000100000111010010100110011;
ROM[4361] <= 32'b00000000101001001000001110110011;
ROM[4362] <= 32'b00000000000100111000001110010011;
ROM[4363] <= 32'b00000000000100111111001110010011;
ROM[4364] <= 32'b00000000011100010010000000100011;
ROM[4365] <= 32'b00000000010000010000000100010011;
ROM[4366] <= 32'b11111111110000010000000100010011;
ROM[4367] <= 32'b00000000000000010010001110000011;
ROM[4368] <= 32'b00000000000000111000101001100011;
ROM[4369] <= 32'b00000000000000000101001110110111;
ROM[4370] <= 32'b10010100100000111000001110010011;
ROM[4371] <= 32'b00000000111000111000001110110011;
ROM[4372] <= 32'b00000000000000111000000011100111;
ROM[4373] <= 32'b00000000000000100010001110000011;
ROM[4374] <= 32'b00000000011100010010000000100011;
ROM[4375] <= 32'b00000000010000010000000100010011;
ROM[4376] <= 32'b00000101010000000000001110010011;
ROM[4377] <= 32'b00000000011100010010000000100011;
ROM[4378] <= 32'b00000000010000010000000100010011;
ROM[4379] <= 32'b11111111110000010000000100010011;
ROM[4380] <= 32'b00000000000000010010001110000011;
ROM[4381] <= 32'b11111111110000010000000100010011;
ROM[4382] <= 32'b00000000000000010010010000000011;
ROM[4383] <= 32'b00000000011101000010010010110011;
ROM[4384] <= 32'b00000000100000111010010100110011;
ROM[4385] <= 32'b00000000101001001000001110110011;
ROM[4386] <= 32'b00000000000100111000001110010011;
ROM[4387] <= 32'b00000000000100111111001110010011;
ROM[4388] <= 32'b00000000011100010010000000100011;
ROM[4389] <= 32'b00000000010000010000000100010011;
ROM[4390] <= 32'b11111111110000010000000100010011;
ROM[4391] <= 32'b00000000000000010010001110000011;
ROM[4392] <= 32'b00000000000000111000101001100011;
ROM[4393] <= 32'b00000000000000000101001110110111;
ROM[4394] <= 32'b10010000000000111000001110010011;
ROM[4395] <= 32'b00000000111000111000001110110011;
ROM[4396] <= 32'b00000000000000111000000011100111;
ROM[4397] <= 32'b00000000000000100010001110000011;
ROM[4398] <= 32'b00000000011100010010000000100011;
ROM[4399] <= 32'b00000000010000010000000100010011;
ROM[4400] <= 32'b00000101010100000000001110010011;
ROM[4401] <= 32'b00000000011100010010000000100011;
ROM[4402] <= 32'b00000000010000010000000100010011;
ROM[4403] <= 32'b11111111110000010000000100010011;
ROM[4404] <= 32'b00000000000000010010001110000011;
ROM[4405] <= 32'b11111111110000010000000100010011;
ROM[4406] <= 32'b00000000000000010010010000000011;
ROM[4407] <= 32'b00000000011101000010010010110011;
ROM[4408] <= 32'b00000000100000111010010100110011;
ROM[4409] <= 32'b00000000101001001000001110110011;
ROM[4410] <= 32'b00000000000100111000001110010011;
ROM[4411] <= 32'b00000000000100111111001110010011;
ROM[4412] <= 32'b00000000011100010010000000100011;
ROM[4413] <= 32'b00000000010000010000000100010011;
ROM[4414] <= 32'b11111111110000010000000100010011;
ROM[4415] <= 32'b00000000000000010010001110000011;
ROM[4416] <= 32'b00000000000000111000101001100011;
ROM[4417] <= 32'b00000000000000000101001110110111;
ROM[4418] <= 32'b10001011100000111000001110010011;
ROM[4419] <= 32'b00000000111000111000001110110011;
ROM[4420] <= 32'b00000000000000111000000011100111;
ROM[4421] <= 32'b00000000000000100010001110000011;
ROM[4422] <= 32'b00000000011100010010000000100011;
ROM[4423] <= 32'b00000000010000010000000100010011;
ROM[4424] <= 32'b00000101011000000000001110010011;
ROM[4425] <= 32'b00000000011100010010000000100011;
ROM[4426] <= 32'b00000000010000010000000100010011;
ROM[4427] <= 32'b11111111110000010000000100010011;
ROM[4428] <= 32'b00000000000000010010001110000011;
ROM[4429] <= 32'b11111111110000010000000100010011;
ROM[4430] <= 32'b00000000000000010010010000000011;
ROM[4431] <= 32'b00000000011101000010010010110011;
ROM[4432] <= 32'b00000000100000111010010100110011;
ROM[4433] <= 32'b00000000101001001000001110110011;
ROM[4434] <= 32'b00000000000100111000001110010011;
ROM[4435] <= 32'b00000000000100111111001110010011;
ROM[4436] <= 32'b00000000011100010010000000100011;
ROM[4437] <= 32'b00000000010000010000000100010011;
ROM[4438] <= 32'b11111111110000010000000100010011;
ROM[4439] <= 32'b00000000000000010010001110000011;
ROM[4440] <= 32'b00000000000000111000101001100011;
ROM[4441] <= 32'b00000000000000000101001110110111;
ROM[4442] <= 32'b10000111000000111000001110010011;
ROM[4443] <= 32'b00000000111000111000001110110011;
ROM[4444] <= 32'b00000000000000111000000011100111;
ROM[4445] <= 32'b00000000000000100010001110000011;
ROM[4446] <= 32'b00000000011100010010000000100011;
ROM[4447] <= 32'b00000000010000010000000100010011;
ROM[4448] <= 32'b00000101011100000000001110010011;
ROM[4449] <= 32'b00000000011100010010000000100011;
ROM[4450] <= 32'b00000000010000010000000100010011;
ROM[4451] <= 32'b11111111110000010000000100010011;
ROM[4452] <= 32'b00000000000000010010001110000011;
ROM[4453] <= 32'b11111111110000010000000100010011;
ROM[4454] <= 32'b00000000000000010010010000000011;
ROM[4455] <= 32'b00000000011101000010010010110011;
ROM[4456] <= 32'b00000000100000111010010100110011;
ROM[4457] <= 32'b00000000101001001000001110110011;
ROM[4458] <= 32'b00000000000100111000001110010011;
ROM[4459] <= 32'b00000000000100111111001110010011;
ROM[4460] <= 32'b00000000011100010010000000100011;
ROM[4461] <= 32'b00000000010000010000000100010011;
ROM[4462] <= 32'b11111111110000010000000100010011;
ROM[4463] <= 32'b00000000000000010010001110000011;
ROM[4464] <= 32'b00000000000000111000101001100011;
ROM[4465] <= 32'b00000000000000000101001110110111;
ROM[4466] <= 32'b10000010100000111000001110010011;
ROM[4467] <= 32'b00000000111000111000001110110011;
ROM[4468] <= 32'b00000000000000111000000011100111;
ROM[4469] <= 32'b00000000000000100010001110000011;
ROM[4470] <= 32'b00000000011100010010000000100011;
ROM[4471] <= 32'b00000000010000010000000100010011;
ROM[4472] <= 32'b00000101100000000000001110010011;
ROM[4473] <= 32'b00000000011100010010000000100011;
ROM[4474] <= 32'b00000000010000010000000100010011;
ROM[4475] <= 32'b11111111110000010000000100010011;
ROM[4476] <= 32'b00000000000000010010001110000011;
ROM[4477] <= 32'b11111111110000010000000100010011;
ROM[4478] <= 32'b00000000000000010010010000000011;
ROM[4479] <= 32'b00000000011101000010010010110011;
ROM[4480] <= 32'b00000000100000111010010100110011;
ROM[4481] <= 32'b00000000101001001000001110110011;
ROM[4482] <= 32'b00000000000100111000001110010011;
ROM[4483] <= 32'b00000000000100111111001110010011;
ROM[4484] <= 32'b00000000011100010010000000100011;
ROM[4485] <= 32'b00000000010000010000000100010011;
ROM[4486] <= 32'b11111111110000010000000100010011;
ROM[4487] <= 32'b00000000000000010010001110000011;
ROM[4488] <= 32'b00000000000000111000101001100011;
ROM[4489] <= 32'b00000000000000000100001110110111;
ROM[4490] <= 32'b01111110000000111000001110010011;
ROM[4491] <= 32'b00000000111000111000001110110011;
ROM[4492] <= 32'b00000000000000111000000011100111;
ROM[4493] <= 32'b00000000000000100010001110000011;
ROM[4494] <= 32'b00000000011100010010000000100011;
ROM[4495] <= 32'b00000000010000010000000100010011;
ROM[4496] <= 32'b00000101100100000000001110010011;
ROM[4497] <= 32'b00000000011100010010000000100011;
ROM[4498] <= 32'b00000000010000010000000100010011;
ROM[4499] <= 32'b11111111110000010000000100010011;
ROM[4500] <= 32'b00000000000000010010001110000011;
ROM[4501] <= 32'b11111111110000010000000100010011;
ROM[4502] <= 32'b00000000000000010010010000000011;
ROM[4503] <= 32'b00000000011101000010010010110011;
ROM[4504] <= 32'b00000000100000111010010100110011;
ROM[4505] <= 32'b00000000101001001000001110110011;
ROM[4506] <= 32'b00000000000100111000001110010011;
ROM[4507] <= 32'b00000000000100111111001110010011;
ROM[4508] <= 32'b00000000011100010010000000100011;
ROM[4509] <= 32'b00000000010000010000000100010011;
ROM[4510] <= 32'b11111111110000010000000100010011;
ROM[4511] <= 32'b00000000000000010010001110000011;
ROM[4512] <= 32'b00000000000000111000101001100011;
ROM[4513] <= 32'b00000000000000000100001110110111;
ROM[4514] <= 32'b01111001100000111000001110010011;
ROM[4515] <= 32'b00000000111000111000001110110011;
ROM[4516] <= 32'b00000000000000111000000011100111;
ROM[4517] <= 32'b00000000000000100010001110000011;
ROM[4518] <= 32'b00000000011100010010000000100011;
ROM[4519] <= 32'b00000000010000010000000100010011;
ROM[4520] <= 32'b00000101101000000000001110010011;
ROM[4521] <= 32'b00000000011100010010000000100011;
ROM[4522] <= 32'b00000000010000010000000100010011;
ROM[4523] <= 32'b11111111110000010000000100010011;
ROM[4524] <= 32'b00000000000000010010001110000011;
ROM[4525] <= 32'b11111111110000010000000100010011;
ROM[4526] <= 32'b00000000000000010010010000000011;
ROM[4527] <= 32'b00000000011101000010010010110011;
ROM[4528] <= 32'b00000000100000111010010100110011;
ROM[4529] <= 32'b00000000101001001000001110110011;
ROM[4530] <= 32'b00000000000100111000001110010011;
ROM[4531] <= 32'b00000000000100111111001110010011;
ROM[4532] <= 32'b00000000011100010010000000100011;
ROM[4533] <= 32'b00000000010000010000000100010011;
ROM[4534] <= 32'b11111111110000010000000100010011;
ROM[4535] <= 32'b00000000000000010010001110000011;
ROM[4536] <= 32'b00000000000000111000101001100011;
ROM[4537] <= 32'b00000000000000000100001110110111;
ROM[4538] <= 32'b01110101000000111000001110010011;
ROM[4539] <= 32'b00000000111000111000001110110011;
ROM[4540] <= 32'b00000000000000111000000011100111;
ROM[4541] <= 32'b00000000000100000000001110010011;
ROM[4542] <= 32'b00000000011100010010000000100011;
ROM[4543] <= 32'b00000000010000010000000100010011;
ROM[4544] <= 32'b11111111110000010000000100010011;
ROM[4545] <= 32'b00000000000000010010001110000011;
ROM[4546] <= 32'b01000000011100000000001110110011;
ROM[4547] <= 32'b00000000011100010010000000100011;
ROM[4548] <= 32'b00000000010000010000000100010011;
ROM[4549] <= 32'b00000001010000000000001110010011;
ROM[4550] <= 32'b01000000011100011000001110110011;
ROM[4551] <= 32'b00000000000000111010000010000011;
ROM[4552] <= 32'b11111111110000010000000100010011;
ROM[4553] <= 32'b00000000000000010010001110000011;
ROM[4554] <= 32'b00000000011100100010000000100011;
ROM[4555] <= 32'b00000000010000100000000100010011;
ROM[4556] <= 32'b00000001010000000000001110010011;
ROM[4557] <= 32'b01000000011100011000001110110011;
ROM[4558] <= 32'b00000000010000111010000110000011;
ROM[4559] <= 32'b00000000100000111010001000000011;
ROM[4560] <= 32'b00000000110000111010001010000011;
ROM[4561] <= 32'b00000001000000111010001100000011;
ROM[4562] <= 32'b00000000000000001000000011100111;
ROM[4563] <= 32'b00000100100000000000000011101111;
ROM[4564] <= 32'b00000101101000000000001110010011;
ROM[4565] <= 32'b00000000011100010010000000100011;
ROM[4566] <= 32'b00000000010000010000000100010011;
ROM[4567] <= 32'b00000001010000000000001110010011;
ROM[4568] <= 32'b01000000011100011000001110110011;
ROM[4569] <= 32'b00000000000000111010000010000011;
ROM[4570] <= 32'b11111111110000010000000100010011;
ROM[4571] <= 32'b00000000000000010010001110000011;
ROM[4572] <= 32'b00000000011100100010000000100011;
ROM[4573] <= 32'b00000000010000100000000100010011;
ROM[4574] <= 32'b00000001010000000000001110010011;
ROM[4575] <= 32'b01000000011100011000001110110011;
ROM[4576] <= 32'b00000000010000111010000110000011;
ROM[4577] <= 32'b00000000100000111010001000000011;
ROM[4578] <= 32'b00000000110000111010001010000011;
ROM[4579] <= 32'b00000001000000111010001100000011;
ROM[4580] <= 32'b00000000000000001000000011100111;
ROM[4581] <= 32'b00000100100000000000000011101111;
ROM[4582] <= 32'b00000101100100000000001110010011;
ROM[4583] <= 32'b00000000011100010010000000100011;
ROM[4584] <= 32'b00000000010000010000000100010011;
ROM[4585] <= 32'b00000001010000000000001110010011;
ROM[4586] <= 32'b01000000011100011000001110110011;
ROM[4587] <= 32'b00000000000000111010000010000011;
ROM[4588] <= 32'b11111111110000010000000100010011;
ROM[4589] <= 32'b00000000000000010010001110000011;
ROM[4590] <= 32'b00000000011100100010000000100011;
ROM[4591] <= 32'b00000000010000100000000100010011;
ROM[4592] <= 32'b00000001010000000000001110010011;
ROM[4593] <= 32'b01000000011100011000001110110011;
ROM[4594] <= 32'b00000000010000111010000110000011;
ROM[4595] <= 32'b00000000100000111010001000000011;
ROM[4596] <= 32'b00000000110000111010001010000011;
ROM[4597] <= 32'b00000001000000111010001100000011;
ROM[4598] <= 32'b00000000000000001000000011100111;
ROM[4599] <= 32'b00000100100000000000000011101111;
ROM[4600] <= 32'b00000101100000000000001110010011;
ROM[4601] <= 32'b00000000011100010010000000100011;
ROM[4602] <= 32'b00000000010000010000000100010011;
ROM[4603] <= 32'b00000001010000000000001110010011;
ROM[4604] <= 32'b01000000011100011000001110110011;
ROM[4605] <= 32'b00000000000000111010000010000011;
ROM[4606] <= 32'b11111111110000010000000100010011;
ROM[4607] <= 32'b00000000000000010010001110000011;
ROM[4608] <= 32'b00000000011100100010000000100011;
ROM[4609] <= 32'b00000000010000100000000100010011;
ROM[4610] <= 32'b00000001010000000000001110010011;
ROM[4611] <= 32'b01000000011100011000001110110011;
ROM[4612] <= 32'b00000000010000111010000110000011;
ROM[4613] <= 32'b00000000100000111010001000000011;
ROM[4614] <= 32'b00000000110000111010001010000011;
ROM[4615] <= 32'b00000001000000111010001100000011;
ROM[4616] <= 32'b00000000000000001000000011100111;
ROM[4617] <= 32'b00000100100000000000000011101111;
ROM[4618] <= 32'b00000101011100000000001110010011;
ROM[4619] <= 32'b00000000011100010010000000100011;
ROM[4620] <= 32'b00000000010000010000000100010011;
ROM[4621] <= 32'b00000001010000000000001110010011;
ROM[4622] <= 32'b01000000011100011000001110110011;
ROM[4623] <= 32'b00000000000000111010000010000011;
ROM[4624] <= 32'b11111111110000010000000100010011;
ROM[4625] <= 32'b00000000000000010010001110000011;
ROM[4626] <= 32'b00000000011100100010000000100011;
ROM[4627] <= 32'b00000000010000100000000100010011;
ROM[4628] <= 32'b00000001010000000000001110010011;
ROM[4629] <= 32'b01000000011100011000001110110011;
ROM[4630] <= 32'b00000000010000111010000110000011;
ROM[4631] <= 32'b00000000100000111010001000000011;
ROM[4632] <= 32'b00000000110000111010001010000011;
ROM[4633] <= 32'b00000001000000111010001100000011;
ROM[4634] <= 32'b00000000000000001000000011100111;
ROM[4635] <= 32'b00000100100000000000000011101111;
ROM[4636] <= 32'b00000101011000000000001110010011;
ROM[4637] <= 32'b00000000011100010010000000100011;
ROM[4638] <= 32'b00000000010000010000000100010011;
ROM[4639] <= 32'b00000001010000000000001110010011;
ROM[4640] <= 32'b01000000011100011000001110110011;
ROM[4641] <= 32'b00000000000000111010000010000011;
ROM[4642] <= 32'b11111111110000010000000100010011;
ROM[4643] <= 32'b00000000000000010010001110000011;
ROM[4644] <= 32'b00000000011100100010000000100011;
ROM[4645] <= 32'b00000000010000100000000100010011;
ROM[4646] <= 32'b00000001010000000000001110010011;
ROM[4647] <= 32'b01000000011100011000001110110011;
ROM[4648] <= 32'b00000000010000111010000110000011;
ROM[4649] <= 32'b00000000100000111010001000000011;
ROM[4650] <= 32'b00000000110000111010001010000011;
ROM[4651] <= 32'b00000001000000111010001100000011;
ROM[4652] <= 32'b00000000000000001000000011100111;
ROM[4653] <= 32'b00000100100000000000000011101111;
ROM[4654] <= 32'b00000101010100000000001110010011;
ROM[4655] <= 32'b00000000011100010010000000100011;
ROM[4656] <= 32'b00000000010000010000000100010011;
ROM[4657] <= 32'b00000001010000000000001110010011;
ROM[4658] <= 32'b01000000011100011000001110110011;
ROM[4659] <= 32'b00000000000000111010000010000011;
ROM[4660] <= 32'b11111111110000010000000100010011;
ROM[4661] <= 32'b00000000000000010010001110000011;
ROM[4662] <= 32'b00000000011100100010000000100011;
ROM[4663] <= 32'b00000000010000100000000100010011;
ROM[4664] <= 32'b00000001010000000000001110010011;
ROM[4665] <= 32'b01000000011100011000001110110011;
ROM[4666] <= 32'b00000000010000111010000110000011;
ROM[4667] <= 32'b00000000100000111010001000000011;
ROM[4668] <= 32'b00000000110000111010001010000011;
ROM[4669] <= 32'b00000001000000111010001100000011;
ROM[4670] <= 32'b00000000000000001000000011100111;
ROM[4671] <= 32'b00000100100000000000000011101111;
ROM[4672] <= 32'b00000101010000000000001110010011;
ROM[4673] <= 32'b00000000011100010010000000100011;
ROM[4674] <= 32'b00000000010000010000000100010011;
ROM[4675] <= 32'b00000001010000000000001110010011;
ROM[4676] <= 32'b01000000011100011000001110110011;
ROM[4677] <= 32'b00000000000000111010000010000011;
ROM[4678] <= 32'b11111111110000010000000100010011;
ROM[4679] <= 32'b00000000000000010010001110000011;
ROM[4680] <= 32'b00000000011100100010000000100011;
ROM[4681] <= 32'b00000000010000100000000100010011;
ROM[4682] <= 32'b00000001010000000000001110010011;
ROM[4683] <= 32'b01000000011100011000001110110011;
ROM[4684] <= 32'b00000000010000111010000110000011;
ROM[4685] <= 32'b00000000100000111010001000000011;
ROM[4686] <= 32'b00000000110000111010001010000011;
ROM[4687] <= 32'b00000001000000111010001100000011;
ROM[4688] <= 32'b00000000000000001000000011100111;
ROM[4689] <= 32'b00000100100000000000000011101111;
ROM[4690] <= 32'b00000101001100000000001110010011;
ROM[4691] <= 32'b00000000011100010010000000100011;
ROM[4692] <= 32'b00000000010000010000000100010011;
ROM[4693] <= 32'b00000001010000000000001110010011;
ROM[4694] <= 32'b01000000011100011000001110110011;
ROM[4695] <= 32'b00000000000000111010000010000011;
ROM[4696] <= 32'b11111111110000010000000100010011;
ROM[4697] <= 32'b00000000000000010010001110000011;
ROM[4698] <= 32'b00000000011100100010000000100011;
ROM[4699] <= 32'b00000000010000100000000100010011;
ROM[4700] <= 32'b00000001010000000000001110010011;
ROM[4701] <= 32'b01000000011100011000001110110011;
ROM[4702] <= 32'b00000000010000111010000110000011;
ROM[4703] <= 32'b00000000100000111010001000000011;
ROM[4704] <= 32'b00000000110000111010001010000011;
ROM[4705] <= 32'b00000001000000111010001100000011;
ROM[4706] <= 32'b00000000000000001000000011100111;
ROM[4707] <= 32'b00000100100000000000000011101111;
ROM[4708] <= 32'b00000101001000000000001110010011;
ROM[4709] <= 32'b00000000011100010010000000100011;
ROM[4710] <= 32'b00000000010000010000000100010011;
ROM[4711] <= 32'b00000001010000000000001110010011;
ROM[4712] <= 32'b01000000011100011000001110110011;
ROM[4713] <= 32'b00000000000000111010000010000011;
ROM[4714] <= 32'b11111111110000010000000100010011;
ROM[4715] <= 32'b00000000000000010010001110000011;
ROM[4716] <= 32'b00000000011100100010000000100011;
ROM[4717] <= 32'b00000000010000100000000100010011;
ROM[4718] <= 32'b00000001010000000000001110010011;
ROM[4719] <= 32'b01000000011100011000001110110011;
ROM[4720] <= 32'b00000000010000111010000110000011;
ROM[4721] <= 32'b00000000100000111010001000000011;
ROM[4722] <= 32'b00000000110000111010001010000011;
ROM[4723] <= 32'b00000001000000111010001100000011;
ROM[4724] <= 32'b00000000000000001000000011100111;
ROM[4725] <= 32'b00000100100000000000000011101111;
ROM[4726] <= 32'b00000101000100000000001110010011;
ROM[4727] <= 32'b00000000011100010010000000100011;
ROM[4728] <= 32'b00000000010000010000000100010011;
ROM[4729] <= 32'b00000001010000000000001110010011;
ROM[4730] <= 32'b01000000011100011000001110110011;
ROM[4731] <= 32'b00000000000000111010000010000011;
ROM[4732] <= 32'b11111111110000010000000100010011;
ROM[4733] <= 32'b00000000000000010010001110000011;
ROM[4734] <= 32'b00000000011100100010000000100011;
ROM[4735] <= 32'b00000000010000100000000100010011;
ROM[4736] <= 32'b00000001010000000000001110010011;
ROM[4737] <= 32'b01000000011100011000001110110011;
ROM[4738] <= 32'b00000000010000111010000110000011;
ROM[4739] <= 32'b00000000100000111010001000000011;
ROM[4740] <= 32'b00000000110000111010001010000011;
ROM[4741] <= 32'b00000001000000111010001100000011;
ROM[4742] <= 32'b00000000000000001000000011100111;
ROM[4743] <= 32'b00000100100000000000000011101111;
ROM[4744] <= 32'b00000101000000000000001110010011;
ROM[4745] <= 32'b00000000011100010010000000100011;
ROM[4746] <= 32'b00000000010000010000000100010011;
ROM[4747] <= 32'b00000001010000000000001110010011;
ROM[4748] <= 32'b01000000011100011000001110110011;
ROM[4749] <= 32'b00000000000000111010000010000011;
ROM[4750] <= 32'b11111111110000010000000100010011;
ROM[4751] <= 32'b00000000000000010010001110000011;
ROM[4752] <= 32'b00000000011100100010000000100011;
ROM[4753] <= 32'b00000000010000100000000100010011;
ROM[4754] <= 32'b00000001010000000000001110010011;
ROM[4755] <= 32'b01000000011100011000001110110011;
ROM[4756] <= 32'b00000000010000111010000110000011;
ROM[4757] <= 32'b00000000100000111010001000000011;
ROM[4758] <= 32'b00000000110000111010001010000011;
ROM[4759] <= 32'b00000001000000111010001100000011;
ROM[4760] <= 32'b00000000000000001000000011100111;
ROM[4761] <= 32'b00000100100000000000000011101111;
ROM[4762] <= 32'b00000100111100000000001110010011;
ROM[4763] <= 32'b00000000011100010010000000100011;
ROM[4764] <= 32'b00000000010000010000000100010011;
ROM[4765] <= 32'b00000001010000000000001110010011;
ROM[4766] <= 32'b01000000011100011000001110110011;
ROM[4767] <= 32'b00000000000000111010000010000011;
ROM[4768] <= 32'b11111111110000010000000100010011;
ROM[4769] <= 32'b00000000000000010010001110000011;
ROM[4770] <= 32'b00000000011100100010000000100011;
ROM[4771] <= 32'b00000000010000100000000100010011;
ROM[4772] <= 32'b00000001010000000000001110010011;
ROM[4773] <= 32'b01000000011100011000001110110011;
ROM[4774] <= 32'b00000000010000111010000110000011;
ROM[4775] <= 32'b00000000100000111010001000000011;
ROM[4776] <= 32'b00000000110000111010001010000011;
ROM[4777] <= 32'b00000001000000111010001100000011;
ROM[4778] <= 32'b00000000000000001000000011100111;
ROM[4779] <= 32'b00000100100000000000000011101111;
ROM[4780] <= 32'b00000100111000000000001110010011;
ROM[4781] <= 32'b00000000011100010010000000100011;
ROM[4782] <= 32'b00000000010000010000000100010011;
ROM[4783] <= 32'b00000001010000000000001110010011;
ROM[4784] <= 32'b01000000011100011000001110110011;
ROM[4785] <= 32'b00000000000000111010000010000011;
ROM[4786] <= 32'b11111111110000010000000100010011;
ROM[4787] <= 32'b00000000000000010010001110000011;
ROM[4788] <= 32'b00000000011100100010000000100011;
ROM[4789] <= 32'b00000000010000100000000100010011;
ROM[4790] <= 32'b00000001010000000000001110010011;
ROM[4791] <= 32'b01000000011100011000001110110011;
ROM[4792] <= 32'b00000000010000111010000110000011;
ROM[4793] <= 32'b00000000100000111010001000000011;
ROM[4794] <= 32'b00000000110000111010001010000011;
ROM[4795] <= 32'b00000001000000111010001100000011;
ROM[4796] <= 32'b00000000000000001000000011100111;
ROM[4797] <= 32'b00000100100000000000000011101111;
ROM[4798] <= 32'b00000100110100000000001110010011;
ROM[4799] <= 32'b00000000011100010010000000100011;
ROM[4800] <= 32'b00000000010000010000000100010011;
ROM[4801] <= 32'b00000001010000000000001110010011;
ROM[4802] <= 32'b01000000011100011000001110110011;
ROM[4803] <= 32'b00000000000000111010000010000011;
ROM[4804] <= 32'b11111111110000010000000100010011;
ROM[4805] <= 32'b00000000000000010010001110000011;
ROM[4806] <= 32'b00000000011100100010000000100011;
ROM[4807] <= 32'b00000000010000100000000100010011;
ROM[4808] <= 32'b00000001010000000000001110010011;
ROM[4809] <= 32'b01000000011100011000001110110011;
ROM[4810] <= 32'b00000000010000111010000110000011;
ROM[4811] <= 32'b00000000100000111010001000000011;
ROM[4812] <= 32'b00000000110000111010001010000011;
ROM[4813] <= 32'b00000001000000111010001100000011;
ROM[4814] <= 32'b00000000000000001000000011100111;
ROM[4815] <= 32'b00000100100000000000000011101111;
ROM[4816] <= 32'b00000100110000000000001110010011;
ROM[4817] <= 32'b00000000011100010010000000100011;
ROM[4818] <= 32'b00000000010000010000000100010011;
ROM[4819] <= 32'b00000001010000000000001110010011;
ROM[4820] <= 32'b01000000011100011000001110110011;
ROM[4821] <= 32'b00000000000000111010000010000011;
ROM[4822] <= 32'b11111111110000010000000100010011;
ROM[4823] <= 32'b00000000000000010010001110000011;
ROM[4824] <= 32'b00000000011100100010000000100011;
ROM[4825] <= 32'b00000000010000100000000100010011;
ROM[4826] <= 32'b00000001010000000000001110010011;
ROM[4827] <= 32'b01000000011100011000001110110011;
ROM[4828] <= 32'b00000000010000111010000110000011;
ROM[4829] <= 32'b00000000100000111010001000000011;
ROM[4830] <= 32'b00000000110000111010001010000011;
ROM[4831] <= 32'b00000001000000111010001100000011;
ROM[4832] <= 32'b00000000000000001000000011100111;
ROM[4833] <= 32'b00000100100000000000000011101111;
ROM[4834] <= 32'b00000100101100000000001110010011;
ROM[4835] <= 32'b00000000011100010010000000100011;
ROM[4836] <= 32'b00000000010000010000000100010011;
ROM[4837] <= 32'b00000001010000000000001110010011;
ROM[4838] <= 32'b01000000011100011000001110110011;
ROM[4839] <= 32'b00000000000000111010000010000011;
ROM[4840] <= 32'b11111111110000010000000100010011;
ROM[4841] <= 32'b00000000000000010010001110000011;
ROM[4842] <= 32'b00000000011100100010000000100011;
ROM[4843] <= 32'b00000000010000100000000100010011;
ROM[4844] <= 32'b00000001010000000000001110010011;
ROM[4845] <= 32'b01000000011100011000001110110011;
ROM[4846] <= 32'b00000000010000111010000110000011;
ROM[4847] <= 32'b00000000100000111010001000000011;
ROM[4848] <= 32'b00000000110000111010001010000011;
ROM[4849] <= 32'b00000001000000111010001100000011;
ROM[4850] <= 32'b00000000000000001000000011100111;
ROM[4851] <= 32'b00000100100000000000000011101111;
ROM[4852] <= 32'b00000100101000000000001110010011;
ROM[4853] <= 32'b00000000011100010010000000100011;
ROM[4854] <= 32'b00000000010000010000000100010011;
ROM[4855] <= 32'b00000001010000000000001110010011;
ROM[4856] <= 32'b01000000011100011000001110110011;
ROM[4857] <= 32'b00000000000000111010000010000011;
ROM[4858] <= 32'b11111111110000010000000100010011;
ROM[4859] <= 32'b00000000000000010010001110000011;
ROM[4860] <= 32'b00000000011100100010000000100011;
ROM[4861] <= 32'b00000000010000100000000100010011;
ROM[4862] <= 32'b00000001010000000000001110010011;
ROM[4863] <= 32'b01000000011100011000001110110011;
ROM[4864] <= 32'b00000000010000111010000110000011;
ROM[4865] <= 32'b00000000100000111010001000000011;
ROM[4866] <= 32'b00000000110000111010001010000011;
ROM[4867] <= 32'b00000001000000111010001100000011;
ROM[4868] <= 32'b00000000000000001000000011100111;
ROM[4869] <= 32'b00000100100000000000000011101111;
ROM[4870] <= 32'b00000100100100000000001110010011;
ROM[4871] <= 32'b00000000011100010010000000100011;
ROM[4872] <= 32'b00000000010000010000000100010011;
ROM[4873] <= 32'b00000001010000000000001110010011;
ROM[4874] <= 32'b01000000011100011000001110110011;
ROM[4875] <= 32'b00000000000000111010000010000011;
ROM[4876] <= 32'b11111111110000010000000100010011;
ROM[4877] <= 32'b00000000000000010010001110000011;
ROM[4878] <= 32'b00000000011100100010000000100011;
ROM[4879] <= 32'b00000000010000100000000100010011;
ROM[4880] <= 32'b00000001010000000000001110010011;
ROM[4881] <= 32'b01000000011100011000001110110011;
ROM[4882] <= 32'b00000000010000111010000110000011;
ROM[4883] <= 32'b00000000100000111010001000000011;
ROM[4884] <= 32'b00000000110000111010001010000011;
ROM[4885] <= 32'b00000001000000111010001100000011;
ROM[4886] <= 32'b00000000000000001000000011100111;
ROM[4887] <= 32'b00000100100000000000000011101111;
ROM[4888] <= 32'b00000100100000000000001110010011;
ROM[4889] <= 32'b00000000011100010010000000100011;
ROM[4890] <= 32'b00000000010000010000000100010011;
ROM[4891] <= 32'b00000001010000000000001110010011;
ROM[4892] <= 32'b01000000011100011000001110110011;
ROM[4893] <= 32'b00000000000000111010000010000011;
ROM[4894] <= 32'b11111111110000010000000100010011;
ROM[4895] <= 32'b00000000000000010010001110000011;
ROM[4896] <= 32'b00000000011100100010000000100011;
ROM[4897] <= 32'b00000000010000100000000100010011;
ROM[4898] <= 32'b00000001010000000000001110010011;
ROM[4899] <= 32'b01000000011100011000001110110011;
ROM[4900] <= 32'b00000000010000111010000110000011;
ROM[4901] <= 32'b00000000100000111010001000000011;
ROM[4902] <= 32'b00000000110000111010001010000011;
ROM[4903] <= 32'b00000001000000111010001100000011;
ROM[4904] <= 32'b00000000000000001000000011100111;
ROM[4905] <= 32'b00000100100000000000000011101111;
ROM[4906] <= 32'b00000100011100000000001110010011;
ROM[4907] <= 32'b00000000011100010010000000100011;
ROM[4908] <= 32'b00000000010000010000000100010011;
ROM[4909] <= 32'b00000001010000000000001110010011;
ROM[4910] <= 32'b01000000011100011000001110110011;
ROM[4911] <= 32'b00000000000000111010000010000011;
ROM[4912] <= 32'b11111111110000010000000100010011;
ROM[4913] <= 32'b00000000000000010010001110000011;
ROM[4914] <= 32'b00000000011100100010000000100011;
ROM[4915] <= 32'b00000000010000100000000100010011;
ROM[4916] <= 32'b00000001010000000000001110010011;
ROM[4917] <= 32'b01000000011100011000001110110011;
ROM[4918] <= 32'b00000000010000111010000110000011;
ROM[4919] <= 32'b00000000100000111010001000000011;
ROM[4920] <= 32'b00000000110000111010001010000011;
ROM[4921] <= 32'b00000001000000111010001100000011;
ROM[4922] <= 32'b00000000000000001000000011100111;
ROM[4923] <= 32'b00000100100000000000000011101111;
ROM[4924] <= 32'b00000100011000000000001110010011;
ROM[4925] <= 32'b00000000011100010010000000100011;
ROM[4926] <= 32'b00000000010000010000000100010011;
ROM[4927] <= 32'b00000001010000000000001110010011;
ROM[4928] <= 32'b01000000011100011000001110110011;
ROM[4929] <= 32'b00000000000000111010000010000011;
ROM[4930] <= 32'b11111111110000010000000100010011;
ROM[4931] <= 32'b00000000000000010010001110000011;
ROM[4932] <= 32'b00000000011100100010000000100011;
ROM[4933] <= 32'b00000000010000100000000100010011;
ROM[4934] <= 32'b00000001010000000000001110010011;
ROM[4935] <= 32'b01000000011100011000001110110011;
ROM[4936] <= 32'b00000000010000111010000110000011;
ROM[4937] <= 32'b00000000100000111010001000000011;
ROM[4938] <= 32'b00000000110000111010001010000011;
ROM[4939] <= 32'b00000001000000111010001100000011;
ROM[4940] <= 32'b00000000000000001000000011100111;
ROM[4941] <= 32'b00000100100000000000000011101111;
ROM[4942] <= 32'b00000100010100000000001110010011;
ROM[4943] <= 32'b00000000011100010010000000100011;
ROM[4944] <= 32'b00000000010000010000000100010011;
ROM[4945] <= 32'b00000001010000000000001110010011;
ROM[4946] <= 32'b01000000011100011000001110110011;
ROM[4947] <= 32'b00000000000000111010000010000011;
ROM[4948] <= 32'b11111111110000010000000100010011;
ROM[4949] <= 32'b00000000000000010010001110000011;
ROM[4950] <= 32'b00000000011100100010000000100011;
ROM[4951] <= 32'b00000000010000100000000100010011;
ROM[4952] <= 32'b00000001010000000000001110010011;
ROM[4953] <= 32'b01000000011100011000001110110011;
ROM[4954] <= 32'b00000000010000111010000110000011;
ROM[4955] <= 32'b00000000100000111010001000000011;
ROM[4956] <= 32'b00000000110000111010001010000011;
ROM[4957] <= 32'b00000001000000111010001100000011;
ROM[4958] <= 32'b00000000000000001000000011100111;
ROM[4959] <= 32'b00000100100000000000000011101111;
ROM[4960] <= 32'b00000100010000000000001110010011;
ROM[4961] <= 32'b00000000011100010010000000100011;
ROM[4962] <= 32'b00000000010000010000000100010011;
ROM[4963] <= 32'b00000001010000000000001110010011;
ROM[4964] <= 32'b01000000011100011000001110110011;
ROM[4965] <= 32'b00000000000000111010000010000011;
ROM[4966] <= 32'b11111111110000010000000100010011;
ROM[4967] <= 32'b00000000000000010010001110000011;
ROM[4968] <= 32'b00000000011100100010000000100011;
ROM[4969] <= 32'b00000000010000100000000100010011;
ROM[4970] <= 32'b00000001010000000000001110010011;
ROM[4971] <= 32'b01000000011100011000001110110011;
ROM[4972] <= 32'b00000000010000111010000110000011;
ROM[4973] <= 32'b00000000100000111010001000000011;
ROM[4974] <= 32'b00000000110000111010001010000011;
ROM[4975] <= 32'b00000001000000111010001100000011;
ROM[4976] <= 32'b00000000000000001000000011100111;
ROM[4977] <= 32'b00000100100000000000000011101111;
ROM[4978] <= 32'b00000100001100000000001110010011;
ROM[4979] <= 32'b00000000011100010010000000100011;
ROM[4980] <= 32'b00000000010000010000000100010011;
ROM[4981] <= 32'b00000001010000000000001110010011;
ROM[4982] <= 32'b01000000011100011000001110110011;
ROM[4983] <= 32'b00000000000000111010000010000011;
ROM[4984] <= 32'b11111111110000010000000100010011;
ROM[4985] <= 32'b00000000000000010010001110000011;
ROM[4986] <= 32'b00000000011100100010000000100011;
ROM[4987] <= 32'b00000000010000100000000100010011;
ROM[4988] <= 32'b00000001010000000000001110010011;
ROM[4989] <= 32'b01000000011100011000001110110011;
ROM[4990] <= 32'b00000000010000111010000110000011;
ROM[4991] <= 32'b00000000100000111010001000000011;
ROM[4992] <= 32'b00000000110000111010001010000011;
ROM[4993] <= 32'b00000001000000111010001100000011;
ROM[4994] <= 32'b00000000000000001000000011100111;
ROM[4995] <= 32'b00000100100000000000000011101111;
ROM[4996] <= 32'b00000100001000000000001110010011;
ROM[4997] <= 32'b00000000011100010010000000100011;
ROM[4998] <= 32'b00000000010000010000000100010011;
ROM[4999] <= 32'b00000001010000000000001110010011;
ROM[5000] <= 32'b01000000011100011000001110110011;
ROM[5001] <= 32'b00000000000000111010000010000011;
ROM[5002] <= 32'b11111111110000010000000100010011;
ROM[5003] <= 32'b00000000000000010010001110000011;
ROM[5004] <= 32'b00000000011100100010000000100011;
ROM[5005] <= 32'b00000000010000100000000100010011;
ROM[5006] <= 32'b00000001010000000000001110010011;
ROM[5007] <= 32'b01000000011100011000001110110011;
ROM[5008] <= 32'b00000000010000111010000110000011;
ROM[5009] <= 32'b00000000100000111010001000000011;
ROM[5010] <= 32'b00000000110000111010001010000011;
ROM[5011] <= 32'b00000001000000111010001100000011;
ROM[5012] <= 32'b00000000000000001000000011100111;
ROM[5013] <= 32'b00000100100000000000000011101111;
ROM[5014] <= 32'b00000100000100000000001110010011;
ROM[5015] <= 32'b00000000011100010010000000100011;
ROM[5016] <= 32'b00000000010000010000000100010011;
ROM[5017] <= 32'b00000001010000000000001110010011;
ROM[5018] <= 32'b01000000011100011000001110110011;
ROM[5019] <= 32'b00000000000000111010000010000011;
ROM[5020] <= 32'b11111111110000010000000100010011;
ROM[5021] <= 32'b00000000000000010010001110000011;
ROM[5022] <= 32'b00000000011100100010000000100011;
ROM[5023] <= 32'b00000000010000100000000100010011;
ROM[5024] <= 32'b00000001010000000000001110010011;
ROM[5025] <= 32'b01000000011100011000001110110011;
ROM[5026] <= 32'b00000000010000111010000110000011;
ROM[5027] <= 32'b00000000100000111010001000000011;
ROM[5028] <= 32'b00000000110000111010001010000011;
ROM[5029] <= 32'b00000001000000111010001100000011;
ROM[5030] <= 32'b00000000000000001000000011100111;
ROM[5031] <= 32'b00000000000000010010000000100011;
ROM[5032] <= 32'b00000000010000010000000100010011;
ROM[5033] <= 32'b00000000000000010010000000100011;
ROM[5034] <= 32'b00000000010000010000000100010011;
ROM[5035] <= 32'b00000000000000010010000000100011;
ROM[5036] <= 32'b00000000010000010000000100010011;
ROM[5037] <= 32'b00000000000000010010000000100011;
ROM[5038] <= 32'b00000000010000010000000100010011;
ROM[5039] <= 32'b00000000000000010010000000100011;
ROM[5040] <= 32'b00000000010000010000000100010011;
ROM[5041] <= 32'b00000000000000010010000000100011;
ROM[5042] <= 32'b00000000010000010000000100010011;
ROM[5043] <= 32'b00000000000000010010000000100011;
ROM[5044] <= 32'b00000000010000010000000100010011;
ROM[5045] <= 32'b00000000000000010010000000100011;
ROM[5046] <= 32'b00000000010000010000000100010011;
ROM[5047] <= 32'b00000000000000010010000000100011;
ROM[5048] <= 32'b00000000010000010000000100010011;
ROM[5049] <= 32'b00000000000000010010000000100011;
ROM[5050] <= 32'b00000000010000010000000100010011;
ROM[5051] <= 32'b00000000000000010010000000100011;
ROM[5052] <= 32'b00000000010000010000000100010011;
ROM[5053] <= 32'b00000000000000010010000000100011;
ROM[5054] <= 32'b00000000010000010000000100010011;
ROM[5055] <= 32'b00000000000000010010000000100011;
ROM[5056] <= 32'b00000000010000010000000100010011;
ROM[5057] <= 32'b00000000000000010010000000100011;
ROM[5058] <= 32'b00000000010000010000000100010011;
ROM[5059] <= 32'b00000000000000010010000000100011;
ROM[5060] <= 32'b00000000010000010000000100010011;
ROM[5061] <= 32'b00000000000000010010000000100011;
ROM[5062] <= 32'b00000000010000010000000100010011;
ROM[5063] <= 32'b00000000010100000000001110010011;
ROM[5064] <= 32'b00000000011100010010000000100011;
ROM[5065] <= 32'b00000000010000010000000100010011;
ROM[5066] <= 32'b00000000000000000101001110110111;
ROM[5067] <= 32'b11110111010000111000001110010011;
ROM[5068] <= 32'b00000000111000111000001110110011;
ROM[5069] <= 32'b00000000011100010010000000100011;
ROM[5070] <= 32'b00000000010000010000000100010011;
ROM[5071] <= 32'b00000000001100010010000000100011;
ROM[5072] <= 32'b00000000010000010000000100010011;
ROM[5073] <= 32'b00000000010000010010000000100011;
ROM[5074] <= 32'b00000000010000010000000100010011;
ROM[5075] <= 32'b00000000010100010010000000100011;
ROM[5076] <= 32'b00000000010000010000000100010011;
ROM[5077] <= 32'b00000000011000010010000000100011;
ROM[5078] <= 32'b00000000010000010000000100010011;
ROM[5079] <= 32'b00000001010000000000001110010011;
ROM[5080] <= 32'b00000000010000111000001110010011;
ROM[5081] <= 32'b01000000011100010000001110110011;
ROM[5082] <= 32'b00000000011100000000001000110011;
ROM[5083] <= 32'b00000000001000000000000110110011;
ROM[5084] <= 32'b10010001000011111011000011101111;
ROM[5085] <= 32'b11111111110000010000000100010011;
ROM[5086] <= 32'b00000000000000010010001110000011;
ROM[5087] <= 32'b00000000011100011010000000100011;
ROM[5088] <= 32'b00000000010000000000001110010011;
ROM[5089] <= 32'b00000000011100010010000000100011;
ROM[5090] <= 32'b00000000010000010000000100010011;
ROM[5091] <= 32'b00000000000000000101001110110111;
ROM[5092] <= 32'b11111101100000111000001110010011;
ROM[5093] <= 32'b00000000111000111000001110110011;
ROM[5094] <= 32'b00000000011100010010000000100011;
ROM[5095] <= 32'b00000000010000010000000100010011;
ROM[5096] <= 32'b00000000001100010010000000100011;
ROM[5097] <= 32'b00000000010000010000000100010011;
ROM[5098] <= 32'b00000000010000010010000000100011;
ROM[5099] <= 32'b00000000010000010000000100010011;
ROM[5100] <= 32'b00000000010100010010000000100011;
ROM[5101] <= 32'b00000000010000010000000100010011;
ROM[5102] <= 32'b00000000011000010010000000100011;
ROM[5103] <= 32'b00000000010000010000000100010011;
ROM[5104] <= 32'b00000001010000000000001110010011;
ROM[5105] <= 32'b00000000010000111000001110010011;
ROM[5106] <= 32'b01000000011100010000001110110011;
ROM[5107] <= 32'b00000000011100000000001000110011;
ROM[5108] <= 32'b00000000001000000000000110110011;
ROM[5109] <= 32'b01110110100000100100000011101111;
ROM[5110] <= 32'b00000100101000000000001110010011;
ROM[5111] <= 32'b00000000011100010010000000100011;
ROM[5112] <= 32'b00000000010000010000000100010011;
ROM[5113] <= 32'b00000000000000000101001110110111;
ROM[5114] <= 32'b00000011000000111000001110010011;
ROM[5115] <= 32'b00000000111000111000001110110011;
ROM[5116] <= 32'b00000000011100010010000000100011;
ROM[5117] <= 32'b00000000010000010000000100010011;
ROM[5118] <= 32'b00000000001100010010000000100011;
ROM[5119] <= 32'b00000000010000010000000100010011;
ROM[5120] <= 32'b00000000010000010010000000100011;
ROM[5121] <= 32'b00000000010000010000000100010011;
ROM[5122] <= 32'b00000000010100010010000000100011;
ROM[5123] <= 32'b00000000010000010000000100010011;
ROM[5124] <= 32'b00000000011000010010000000100011;
ROM[5125] <= 32'b00000000010000010000000100010011;
ROM[5126] <= 32'b00000001010000000000001110010011;
ROM[5127] <= 32'b00000000100000111000001110010011;
ROM[5128] <= 32'b01000000011100010000001110110011;
ROM[5129] <= 32'b00000000011100000000001000110011;
ROM[5130] <= 32'b00000000001000000000000110110011;
ROM[5131] <= 32'b00111000000100100100000011101111;
ROM[5132] <= 32'b00000100000100000000001110010011;
ROM[5133] <= 32'b00000000011100010010000000100011;
ROM[5134] <= 32'b00000000010000010000000100010011;
ROM[5135] <= 32'b00000000000000000101001110110111;
ROM[5136] <= 32'b00001000100000111000001110010011;
ROM[5137] <= 32'b00000000111000111000001110110011;
ROM[5138] <= 32'b00000000011100010010000000100011;
ROM[5139] <= 32'b00000000010000010000000100010011;
ROM[5140] <= 32'b00000000001100010010000000100011;
ROM[5141] <= 32'b00000000010000010000000100010011;
ROM[5142] <= 32'b00000000010000010010000000100011;
ROM[5143] <= 32'b00000000010000010000000100010011;
ROM[5144] <= 32'b00000000010100010010000000100011;
ROM[5145] <= 32'b00000000010000010000000100010011;
ROM[5146] <= 32'b00000000011000010010000000100011;
ROM[5147] <= 32'b00000000010000010000000100010011;
ROM[5148] <= 32'b00000001010000000000001110010011;
ROM[5149] <= 32'b00000000100000111000001110010011;
ROM[5150] <= 32'b01000000011100010000001110110011;
ROM[5151] <= 32'b00000000011100000000001000110011;
ROM[5152] <= 32'b00000000001000000000000110110011;
ROM[5153] <= 32'b00110010100100100100000011101111;
ROM[5154] <= 32'b00000100001100000000001110010011;
ROM[5155] <= 32'b00000000011100010010000000100011;
ROM[5156] <= 32'b00000000010000010000000100010011;
ROM[5157] <= 32'b00000000000000000101001110110111;
ROM[5158] <= 32'b00001110000000111000001110010011;
ROM[5159] <= 32'b00000000111000111000001110110011;
ROM[5160] <= 32'b00000000011100010010000000100011;
ROM[5161] <= 32'b00000000010000010000000100010011;
ROM[5162] <= 32'b00000000001100010010000000100011;
ROM[5163] <= 32'b00000000010000010000000100010011;
ROM[5164] <= 32'b00000000010000010010000000100011;
ROM[5165] <= 32'b00000000010000010000000100010011;
ROM[5166] <= 32'b00000000010100010010000000100011;
ROM[5167] <= 32'b00000000010000010000000100010011;
ROM[5168] <= 32'b00000000011000010010000000100011;
ROM[5169] <= 32'b00000000010000010000000100010011;
ROM[5170] <= 32'b00000001010000000000001110010011;
ROM[5171] <= 32'b00000000100000111000001110010011;
ROM[5172] <= 32'b01000000011100010000001110110011;
ROM[5173] <= 32'b00000000011100000000001000110011;
ROM[5174] <= 32'b00000000001000000000000110110011;
ROM[5175] <= 32'b00101101000100100100000011101111;
ROM[5176] <= 32'b00000100101100000000001110010011;
ROM[5177] <= 32'b00000000011100010010000000100011;
ROM[5178] <= 32'b00000000010000010000000100010011;
ROM[5179] <= 32'b00000000000000000101001110110111;
ROM[5180] <= 32'b00010011100000111000001110010011;
ROM[5181] <= 32'b00000000111000111000001110110011;
ROM[5182] <= 32'b00000000011100010010000000100011;
ROM[5183] <= 32'b00000000010000010000000100010011;
ROM[5184] <= 32'b00000000001100010010000000100011;
ROM[5185] <= 32'b00000000010000010000000100010011;
ROM[5186] <= 32'b00000000010000010010000000100011;
ROM[5187] <= 32'b00000000010000010000000100010011;
ROM[5188] <= 32'b00000000010100010010000000100011;
ROM[5189] <= 32'b00000000010000010000000100010011;
ROM[5190] <= 32'b00000000011000010010000000100011;
ROM[5191] <= 32'b00000000010000010000000100010011;
ROM[5192] <= 32'b00000001010000000000001110010011;
ROM[5193] <= 32'b00000000100000111000001110010011;
ROM[5194] <= 32'b01000000011100010000001110110011;
ROM[5195] <= 32'b00000000011100000000001000110011;
ROM[5196] <= 32'b00000000001000000000000110110011;
ROM[5197] <= 32'b00100111100100100100000011101111;
ROM[5198] <= 32'b00000000000000011010001110000011;
ROM[5199] <= 32'b00000000011100010010000000100011;
ROM[5200] <= 32'b00000000010000010000000100010011;
ROM[5201] <= 32'b00000000000000000000001110010011;
ROM[5202] <= 32'b00000000011100010010000000100011;
ROM[5203] <= 32'b00000000010000010000000100010011;
ROM[5204] <= 32'b00000000010000000000001110010011;
ROM[5205] <= 32'b00000000011100010010000000100011;
ROM[5206] <= 32'b00000000010000010000000100010011;
ROM[5207] <= 32'b00000000000000000101001110110111;
ROM[5208] <= 32'b00011010100000111000001110010011;
ROM[5209] <= 32'b00000000111000111000001110110011;
ROM[5210] <= 32'b00000000011100010010000000100011;
ROM[5211] <= 32'b00000000010000010000000100010011;
ROM[5212] <= 32'b00000000001100010010000000100011;
ROM[5213] <= 32'b00000000010000010000000100010011;
ROM[5214] <= 32'b00000000010000010010000000100011;
ROM[5215] <= 32'b00000000010000010000000100010011;
ROM[5216] <= 32'b00000000010100010010000000100011;
ROM[5217] <= 32'b00000000010000010000000100010011;
ROM[5218] <= 32'b00000000011000010010000000100011;
ROM[5219] <= 32'b00000000010000010000000100010011;
ROM[5220] <= 32'b00000001010000000000001110010011;
ROM[5221] <= 32'b00000000100000111000001110010011;
ROM[5222] <= 32'b01000000011100010000001110110011;
ROM[5223] <= 32'b00000000011100000000001000110011;
ROM[5224] <= 32'b00000000001000000000000110110011;
ROM[5225] <= 32'b01101000100000001100000011101111;
ROM[5226] <= 32'b11111111110000010000000100010011;
ROM[5227] <= 32'b00000000000000010010001110000011;
ROM[5228] <= 32'b11111111110000010000000100010011;
ROM[5229] <= 32'b00000000000000010010010000000011;
ROM[5230] <= 32'b00000000011101000000001110110011;
ROM[5231] <= 32'b00000000011100010010000000100011;
ROM[5232] <= 32'b00000000010000010000000100010011;
ROM[5233] <= 32'b11111111110000010000000100010011;
ROM[5234] <= 32'b00000000000000010010001110000011;
ROM[5235] <= 32'b00000000000000111000001100010011;
ROM[5236] <= 32'b11111111110000010000000100010011;
ROM[5237] <= 32'b00000000000000010010001110000011;
ROM[5238] <= 32'b00000000110100110000010000110011;
ROM[5239] <= 32'b00000000011101000010000000100011;
ROM[5240] <= 32'b00000000101100000000001110010011;
ROM[5241] <= 32'b00000000011100010010000000100011;
ROM[5242] <= 32'b00000000010000010000000100010011;
ROM[5243] <= 32'b00000000000000000101001110110111;
ROM[5244] <= 32'b00100011100000111000001110010011;
ROM[5245] <= 32'b00000000111000111000001110110011;
ROM[5246] <= 32'b00000000011100010010000000100011;
ROM[5247] <= 32'b00000000010000010000000100010011;
ROM[5248] <= 32'b00000000001100010010000000100011;
ROM[5249] <= 32'b00000000010000010000000100010011;
ROM[5250] <= 32'b00000000010000010010000000100011;
ROM[5251] <= 32'b00000000010000010000000100010011;
ROM[5252] <= 32'b00000000010100010010000000100011;
ROM[5253] <= 32'b00000000010000010000000100010011;
ROM[5254] <= 32'b00000000011000010010000000100011;
ROM[5255] <= 32'b00000000010000010000000100010011;
ROM[5256] <= 32'b00000001010000000000001110010011;
ROM[5257] <= 32'b00000000010000111000001110010011;
ROM[5258] <= 32'b01000000011100010000001110110011;
ROM[5259] <= 32'b00000000011100000000001000110011;
ROM[5260] <= 32'b00000000001000000000000110110011;
ROM[5261] <= 32'b01010000100000100100000011101111;
ROM[5262] <= 32'b00000101000000000000001110010011;
ROM[5263] <= 32'b00000000011100010010000000100011;
ROM[5264] <= 32'b00000000010000010000000100010011;
ROM[5265] <= 32'b00000000000000000101001110110111;
ROM[5266] <= 32'b00101001000000111000001110010011;
ROM[5267] <= 32'b00000000111000111000001110110011;
ROM[5268] <= 32'b00000000011100010010000000100011;
ROM[5269] <= 32'b00000000010000010000000100010011;
ROM[5270] <= 32'b00000000001100010010000000100011;
ROM[5271] <= 32'b00000000010000010000000100010011;
ROM[5272] <= 32'b00000000010000010010000000100011;
ROM[5273] <= 32'b00000000010000010000000100010011;
ROM[5274] <= 32'b00000000010100010010000000100011;
ROM[5275] <= 32'b00000000010000010000000100010011;
ROM[5276] <= 32'b00000000011000010010000000100011;
ROM[5277] <= 32'b00000000010000010000000100010011;
ROM[5278] <= 32'b00000001010000000000001110010011;
ROM[5279] <= 32'b00000000100000111000001110010011;
ROM[5280] <= 32'b01000000011100010000001110110011;
ROM[5281] <= 32'b00000000011100000000001000110011;
ROM[5282] <= 32'b00000000001000000000000110110011;
ROM[5283] <= 32'b00010010000100100100000011101111;
ROM[5284] <= 32'b00000101001000000000001110010011;
ROM[5285] <= 32'b00000000011100010010000000100011;
ROM[5286] <= 32'b00000000010000010000000100010011;
ROM[5287] <= 32'b00000000000000000101001110110111;
ROM[5288] <= 32'b00101110100000111000001110010011;
ROM[5289] <= 32'b00000000111000111000001110110011;
ROM[5290] <= 32'b00000000011100010010000000100011;
ROM[5291] <= 32'b00000000010000010000000100010011;
ROM[5292] <= 32'b00000000001100010010000000100011;
ROM[5293] <= 32'b00000000010000010000000100010011;
ROM[5294] <= 32'b00000000010000010010000000100011;
ROM[5295] <= 32'b00000000010000010000000100010011;
ROM[5296] <= 32'b00000000010100010010000000100011;
ROM[5297] <= 32'b00000000010000010000000100010011;
ROM[5298] <= 32'b00000000011000010010000000100011;
ROM[5299] <= 32'b00000000010000010000000100010011;
ROM[5300] <= 32'b00000001010000000000001110010011;
ROM[5301] <= 32'b00000000100000111000001110010011;
ROM[5302] <= 32'b01000000011100010000001110110011;
ROM[5303] <= 32'b00000000011100000000001000110011;
ROM[5304] <= 32'b00000000001000000000000110110011;
ROM[5305] <= 32'b00001100100100100100000011101111;
ROM[5306] <= 32'b00000100111100000000001110010011;
ROM[5307] <= 32'b00000000011100010010000000100011;
ROM[5308] <= 32'b00000000010000010000000100010011;
ROM[5309] <= 32'b00000000000000000101001110110111;
ROM[5310] <= 32'b00110100000000111000001110010011;
ROM[5311] <= 32'b00000000111000111000001110110011;
ROM[5312] <= 32'b00000000011100010010000000100011;
ROM[5313] <= 32'b00000000010000010000000100010011;
ROM[5314] <= 32'b00000000001100010010000000100011;
ROM[5315] <= 32'b00000000010000010000000100010011;
ROM[5316] <= 32'b00000000010000010010000000100011;
ROM[5317] <= 32'b00000000010000010000000100010011;
ROM[5318] <= 32'b00000000010100010010000000100011;
ROM[5319] <= 32'b00000000010000010000000100010011;
ROM[5320] <= 32'b00000000011000010010000000100011;
ROM[5321] <= 32'b00000000010000010000000100010011;
ROM[5322] <= 32'b00000001010000000000001110010011;
ROM[5323] <= 32'b00000000100000111000001110010011;
ROM[5324] <= 32'b01000000011100010000001110110011;
ROM[5325] <= 32'b00000000011100000000001000110011;
ROM[5326] <= 32'b00000000001000000000000110110011;
ROM[5327] <= 32'b00000111000100100100000011101111;
ROM[5328] <= 32'b00000100011100000000001110010011;
ROM[5329] <= 32'b00000000011100010010000000100011;
ROM[5330] <= 32'b00000000010000010000000100010011;
ROM[5331] <= 32'b00000000000000000101001110110111;
ROM[5332] <= 32'b00111001100000111000001110010011;
ROM[5333] <= 32'b00000000111000111000001110110011;
ROM[5334] <= 32'b00000000011100010010000000100011;
ROM[5335] <= 32'b00000000010000010000000100010011;
ROM[5336] <= 32'b00000000001100010010000000100011;
ROM[5337] <= 32'b00000000010000010000000100010011;
ROM[5338] <= 32'b00000000010000010010000000100011;
ROM[5339] <= 32'b00000000010000010000000100010011;
ROM[5340] <= 32'b00000000010100010010000000100011;
ROM[5341] <= 32'b00000000010000010000000100010011;
ROM[5342] <= 32'b00000000011000010010000000100011;
ROM[5343] <= 32'b00000000010000010000000100010011;
ROM[5344] <= 32'b00000001010000000000001110010011;
ROM[5345] <= 32'b00000000100000111000001110010011;
ROM[5346] <= 32'b01000000011100010000001110110011;
ROM[5347] <= 32'b00000000011100000000001000110011;
ROM[5348] <= 32'b00000000001000000000000110110011;
ROM[5349] <= 32'b00000001100100100100000011101111;
ROM[5350] <= 32'b00000101001000000000001110010011;
ROM[5351] <= 32'b00000000011100010010000000100011;
ROM[5352] <= 32'b00000000010000010000000100010011;
ROM[5353] <= 32'b00000000000000000101001110110111;
ROM[5354] <= 32'b00111111000000111000001110010011;
ROM[5355] <= 32'b00000000111000111000001110110011;
ROM[5356] <= 32'b00000000011100010010000000100011;
ROM[5357] <= 32'b00000000010000010000000100010011;
ROM[5358] <= 32'b00000000001100010010000000100011;
ROM[5359] <= 32'b00000000010000010000000100010011;
ROM[5360] <= 32'b00000000010000010010000000100011;
ROM[5361] <= 32'b00000000010000010000000100010011;
ROM[5362] <= 32'b00000000010100010010000000100011;
ROM[5363] <= 32'b00000000010000010000000100010011;
ROM[5364] <= 32'b00000000011000010010000000100011;
ROM[5365] <= 32'b00000000010000010000000100010011;
ROM[5366] <= 32'b00000001010000000000001110010011;
ROM[5367] <= 32'b00000000100000111000001110010011;
ROM[5368] <= 32'b01000000011100010000001110110011;
ROM[5369] <= 32'b00000000011100000000001000110011;
ROM[5370] <= 32'b00000000001000000000000110110011;
ROM[5371] <= 32'b01111100000000100100000011101111;
ROM[5372] <= 32'b00000100000100000000001110010011;
ROM[5373] <= 32'b00000000011100010010000000100011;
ROM[5374] <= 32'b00000000010000010000000100010011;
ROM[5375] <= 32'b00000000000000000101001110110111;
ROM[5376] <= 32'b01000100100000111000001110010011;
ROM[5377] <= 32'b00000000111000111000001110110011;
ROM[5378] <= 32'b00000000011100010010000000100011;
ROM[5379] <= 32'b00000000010000010000000100010011;
ROM[5380] <= 32'b00000000001100010010000000100011;
ROM[5381] <= 32'b00000000010000010000000100010011;
ROM[5382] <= 32'b00000000010000010010000000100011;
ROM[5383] <= 32'b00000000010000010000000100010011;
ROM[5384] <= 32'b00000000010100010010000000100011;
ROM[5385] <= 32'b00000000010000010000000100010011;
ROM[5386] <= 32'b00000000011000010010000000100011;
ROM[5387] <= 32'b00000000010000010000000100010011;
ROM[5388] <= 32'b00000001010000000000001110010011;
ROM[5389] <= 32'b00000000100000111000001110010011;
ROM[5390] <= 32'b01000000011100010000001110110011;
ROM[5391] <= 32'b00000000011100000000001000110011;
ROM[5392] <= 32'b00000000001000000000000110110011;
ROM[5393] <= 32'b01110110100000100100000011101111;
ROM[5394] <= 32'b00000100110100000000001110010011;
ROM[5395] <= 32'b00000000011100010010000000100011;
ROM[5396] <= 32'b00000000010000010000000100010011;
ROM[5397] <= 32'b00000000000000000101001110110111;
ROM[5398] <= 32'b01001010000000111000001110010011;
ROM[5399] <= 32'b00000000111000111000001110110011;
ROM[5400] <= 32'b00000000011100010010000000100011;
ROM[5401] <= 32'b00000000010000010000000100010011;
ROM[5402] <= 32'b00000000001100010010000000100011;
ROM[5403] <= 32'b00000000010000010000000100010011;
ROM[5404] <= 32'b00000000010000010010000000100011;
ROM[5405] <= 32'b00000000010000010000000100010011;
ROM[5406] <= 32'b00000000010100010010000000100011;
ROM[5407] <= 32'b00000000010000010000000100010011;
ROM[5408] <= 32'b00000000011000010010000000100011;
ROM[5409] <= 32'b00000000010000010000000100010011;
ROM[5410] <= 32'b00000001010000000000001110010011;
ROM[5411] <= 32'b00000000100000111000001110010011;
ROM[5412] <= 32'b01000000011100010000001110110011;
ROM[5413] <= 32'b00000000011100000000001000110011;
ROM[5414] <= 32'b00000000001000000000000110110011;
ROM[5415] <= 32'b01110001000000100100000011101111;
ROM[5416] <= 32'b00000100110100000000001110010011;
ROM[5417] <= 32'b00000000011100010010000000100011;
ROM[5418] <= 32'b00000000010000010000000100010011;
ROM[5419] <= 32'b00000000000000000101001110110111;
ROM[5420] <= 32'b01001111100000111000001110010011;
ROM[5421] <= 32'b00000000111000111000001110110011;
ROM[5422] <= 32'b00000000011100010010000000100011;
ROM[5423] <= 32'b00000000010000010000000100010011;
ROM[5424] <= 32'b00000000001100010010000000100011;
ROM[5425] <= 32'b00000000010000010000000100010011;
ROM[5426] <= 32'b00000000010000010010000000100011;
ROM[5427] <= 32'b00000000010000010000000100010011;
ROM[5428] <= 32'b00000000010100010010000000100011;
ROM[5429] <= 32'b00000000010000010000000100010011;
ROM[5430] <= 32'b00000000011000010010000000100011;
ROM[5431] <= 32'b00000000010000010000000100010011;
ROM[5432] <= 32'b00000001010000000000001110010011;
ROM[5433] <= 32'b00000000100000111000001110010011;
ROM[5434] <= 32'b01000000011100010000001110110011;
ROM[5435] <= 32'b00000000011100000000001000110011;
ROM[5436] <= 32'b00000000001000000000000110110011;
ROM[5437] <= 32'b01101011100000100100000011101111;
ROM[5438] <= 32'b00000100100100000000001110010011;
ROM[5439] <= 32'b00000000011100010010000000100011;
ROM[5440] <= 32'b00000000010000010000000100010011;
ROM[5441] <= 32'b00000000000000000101001110110111;
ROM[5442] <= 32'b01010101000000111000001110010011;
ROM[5443] <= 32'b00000000111000111000001110110011;
ROM[5444] <= 32'b00000000011100010010000000100011;
ROM[5445] <= 32'b00000000010000010000000100010011;
ROM[5446] <= 32'b00000000001100010010000000100011;
ROM[5447] <= 32'b00000000010000010000000100010011;
ROM[5448] <= 32'b00000000010000010010000000100011;
ROM[5449] <= 32'b00000000010000010000000100010011;
ROM[5450] <= 32'b00000000010100010010000000100011;
ROM[5451] <= 32'b00000000010000010000000100010011;
ROM[5452] <= 32'b00000000011000010010000000100011;
ROM[5453] <= 32'b00000000010000010000000100010011;
ROM[5454] <= 32'b00000001010000000000001110010011;
ROM[5455] <= 32'b00000000100000111000001110010011;
ROM[5456] <= 32'b01000000011100010000001110110011;
ROM[5457] <= 32'b00000000011100000000001000110011;
ROM[5458] <= 32'b00000000001000000000000110110011;
ROM[5459] <= 32'b01100110000000100100000011101111;
ROM[5460] <= 32'b00000100111000000000001110010011;
ROM[5461] <= 32'b00000000011100010010000000100011;
ROM[5462] <= 32'b00000000010000010000000100010011;
ROM[5463] <= 32'b00000000000000000101001110110111;
ROM[5464] <= 32'b01011010100000111000001110010011;
ROM[5465] <= 32'b00000000111000111000001110110011;
ROM[5466] <= 32'b00000000011100010010000000100011;
ROM[5467] <= 32'b00000000010000010000000100010011;
ROM[5468] <= 32'b00000000001100010010000000100011;
ROM[5469] <= 32'b00000000010000010000000100010011;
ROM[5470] <= 32'b00000000010000010010000000100011;
ROM[5471] <= 32'b00000000010000010000000100010011;
ROM[5472] <= 32'b00000000010100010010000000100011;
ROM[5473] <= 32'b00000000010000010000000100010011;
ROM[5474] <= 32'b00000000011000010010000000100011;
ROM[5475] <= 32'b00000000010000010000000100010011;
ROM[5476] <= 32'b00000001010000000000001110010011;
ROM[5477] <= 32'b00000000100000111000001110010011;
ROM[5478] <= 32'b01000000011100010000001110110011;
ROM[5479] <= 32'b00000000011100000000001000110011;
ROM[5480] <= 32'b00000000001000000000000110110011;
ROM[5481] <= 32'b01100000100000100100000011101111;
ROM[5482] <= 32'b00000100011100000000001110010011;
ROM[5483] <= 32'b00000000011100010010000000100011;
ROM[5484] <= 32'b00000000010000010000000100010011;
ROM[5485] <= 32'b00000000000000000101001110110111;
ROM[5486] <= 32'b01100000000000111000001110010011;
ROM[5487] <= 32'b00000000111000111000001110110011;
ROM[5488] <= 32'b00000000011100010010000000100011;
ROM[5489] <= 32'b00000000010000010000000100010011;
ROM[5490] <= 32'b00000000001100010010000000100011;
ROM[5491] <= 32'b00000000010000010000000100010011;
ROM[5492] <= 32'b00000000010000010010000000100011;
ROM[5493] <= 32'b00000000010000010000000100010011;
ROM[5494] <= 32'b00000000010100010010000000100011;
ROM[5495] <= 32'b00000000010000010000000100010011;
ROM[5496] <= 32'b00000000011000010010000000100011;
ROM[5497] <= 32'b00000000010000010000000100010011;
ROM[5498] <= 32'b00000001010000000000001110010011;
ROM[5499] <= 32'b00000000100000111000001110010011;
ROM[5500] <= 32'b01000000011100010000001110110011;
ROM[5501] <= 32'b00000000011100000000001000110011;
ROM[5502] <= 32'b00000000001000000000000110110011;
ROM[5503] <= 32'b01011011000000100100000011101111;
ROM[5504] <= 32'b00000000000000011010001110000011;
ROM[5505] <= 32'b00000000011100010010000000100011;
ROM[5506] <= 32'b00000000010000010000000100010011;
ROM[5507] <= 32'b00000000000100000000001110010011;
ROM[5508] <= 32'b00000000011100010010000000100011;
ROM[5509] <= 32'b00000000010000010000000100010011;
ROM[5510] <= 32'b00000000010000000000001110010011;
ROM[5511] <= 32'b00000000011100010010000000100011;
ROM[5512] <= 32'b00000000010000010000000100010011;
ROM[5513] <= 32'b00000000000000000101001110110111;
ROM[5514] <= 32'b01100111000000111000001110010011;
ROM[5515] <= 32'b00000000111000111000001110110011;
ROM[5516] <= 32'b00000000011100010010000000100011;
ROM[5517] <= 32'b00000000010000010000000100010011;
ROM[5518] <= 32'b00000000001100010010000000100011;
ROM[5519] <= 32'b00000000010000010000000100010011;
ROM[5520] <= 32'b00000000010000010010000000100011;
ROM[5521] <= 32'b00000000010000010000000100010011;
ROM[5522] <= 32'b00000000010100010010000000100011;
ROM[5523] <= 32'b00000000010000010000000100010011;
ROM[5524] <= 32'b00000000011000010010000000100011;
ROM[5525] <= 32'b00000000010000010000000100010011;
ROM[5526] <= 32'b00000001010000000000001110010011;
ROM[5527] <= 32'b00000000100000111000001110010011;
ROM[5528] <= 32'b01000000011100010000001110110011;
ROM[5529] <= 32'b00000000011100000000001000110011;
ROM[5530] <= 32'b00000000001000000000000110110011;
ROM[5531] <= 32'b00011100000000001100000011101111;
ROM[5532] <= 32'b11111111110000010000000100010011;
ROM[5533] <= 32'b00000000000000010010001110000011;
ROM[5534] <= 32'b11111111110000010000000100010011;
ROM[5535] <= 32'b00000000000000010010010000000011;
ROM[5536] <= 32'b00000000011101000000001110110011;
ROM[5537] <= 32'b00000000011100010010000000100011;
ROM[5538] <= 32'b00000000010000010000000100010011;
ROM[5539] <= 32'b11111111110000010000000100010011;
ROM[5540] <= 32'b00000000000000010010001110000011;
ROM[5541] <= 32'b00000000000000111000001100010011;
ROM[5542] <= 32'b11111111110000010000000100010011;
ROM[5543] <= 32'b00000000000000010010001110000011;
ROM[5544] <= 32'b00000000110100110000010000110011;
ROM[5545] <= 32'b00000000011101000010000000100011;
ROM[5546] <= 32'b00000000100000000000001110010011;
ROM[5547] <= 32'b00000000011100010010000000100011;
ROM[5548] <= 32'b00000000010000010000000100010011;
ROM[5549] <= 32'b00000000000000000101001110110111;
ROM[5550] <= 32'b01110000000000111000001110010011;
ROM[5551] <= 32'b00000000111000111000001110110011;
ROM[5552] <= 32'b00000000011100010010000000100011;
ROM[5553] <= 32'b00000000010000010000000100010011;
ROM[5554] <= 32'b00000000001100010010000000100011;
ROM[5555] <= 32'b00000000010000010000000100010011;
ROM[5556] <= 32'b00000000010000010010000000100011;
ROM[5557] <= 32'b00000000010000010000000100010011;
ROM[5558] <= 32'b00000000010100010010000000100011;
ROM[5559] <= 32'b00000000010000010000000100010011;
ROM[5560] <= 32'b00000000011000010010000000100011;
ROM[5561] <= 32'b00000000010000010000000100010011;
ROM[5562] <= 32'b00000001010000000000001110010011;
ROM[5563] <= 32'b00000000010000111000001110010011;
ROM[5564] <= 32'b01000000011100010000001110110011;
ROM[5565] <= 32'b00000000011100000000001000110011;
ROM[5566] <= 32'b00000000001000000000000110110011;
ROM[5567] <= 32'b00000100000000100100000011101111;
ROM[5568] <= 32'b00000100110000000000001110010011;
ROM[5569] <= 32'b00000000011100010010000000100011;
ROM[5570] <= 32'b00000000010000010000000100010011;
ROM[5571] <= 32'b00000000000000000101001110110111;
ROM[5572] <= 32'b01110101100000111000001110010011;
ROM[5573] <= 32'b00000000111000111000001110110011;
ROM[5574] <= 32'b00000000011100010010000000100011;
ROM[5575] <= 32'b00000000010000010000000100010011;
ROM[5576] <= 32'b00000000001100010010000000100011;
ROM[5577] <= 32'b00000000010000010000000100010011;
ROM[5578] <= 32'b00000000010000010010000000100011;
ROM[5579] <= 32'b00000000010000010000000100010011;
ROM[5580] <= 32'b00000000010100010010000000100011;
ROM[5581] <= 32'b00000000010000010000000100010011;
ROM[5582] <= 32'b00000000011000010010000000100011;
ROM[5583] <= 32'b00000000010000010000000100010011;
ROM[5584] <= 32'b00000001010000000000001110010011;
ROM[5585] <= 32'b00000000100000111000001110010011;
ROM[5586] <= 32'b01000000011100010000001110110011;
ROM[5587] <= 32'b00000000011100000000001000110011;
ROM[5588] <= 32'b00000000001000000000000110110011;
ROM[5589] <= 32'b01000101100000100100000011101111;
ROM[5590] <= 32'b00000100000100000000001110010011;
ROM[5591] <= 32'b00000000011100010010000000100011;
ROM[5592] <= 32'b00000000010000010000000100010011;
ROM[5593] <= 32'b00000000000000000101001110110111;
ROM[5594] <= 32'b01111011000000111000001110010011;
ROM[5595] <= 32'b00000000111000111000001110110011;
ROM[5596] <= 32'b00000000011100010010000000100011;
ROM[5597] <= 32'b00000000010000010000000100010011;
ROM[5598] <= 32'b00000000001100010010000000100011;
ROM[5599] <= 32'b00000000010000010000000100010011;
ROM[5600] <= 32'b00000000010000010010000000100011;
ROM[5601] <= 32'b00000000010000010000000100010011;
ROM[5602] <= 32'b00000000010100010010000000100011;
ROM[5603] <= 32'b00000000010000010000000100010011;
ROM[5604] <= 32'b00000000011000010010000000100011;
ROM[5605] <= 32'b00000000010000010000000100010011;
ROM[5606] <= 32'b00000001010000000000001110010011;
ROM[5607] <= 32'b00000000100000111000001110010011;
ROM[5608] <= 32'b01000000011100010000001110110011;
ROM[5609] <= 32'b00000000011100000000001000110011;
ROM[5610] <= 32'b00000000001000000000000110110011;
ROM[5611] <= 32'b01000000000000100100000011101111;
ROM[5612] <= 32'b00000100111000000000001110010011;
ROM[5613] <= 32'b00000000011100010010000000100011;
ROM[5614] <= 32'b00000000010000010000000100010011;
ROM[5615] <= 32'b00000000000000000110001110110111;
ROM[5616] <= 32'b10000000100000111000001110010011;
ROM[5617] <= 32'b00000000111000111000001110110011;
ROM[5618] <= 32'b00000000011100010010000000100011;
ROM[5619] <= 32'b00000000010000010000000100010011;
ROM[5620] <= 32'b00000000001100010010000000100011;
ROM[5621] <= 32'b00000000010000010000000100010011;
ROM[5622] <= 32'b00000000010000010010000000100011;
ROM[5623] <= 32'b00000000010000010000000100010011;
ROM[5624] <= 32'b00000000010100010010000000100011;
ROM[5625] <= 32'b00000000010000010000000100010011;
ROM[5626] <= 32'b00000000011000010010000000100011;
ROM[5627] <= 32'b00000000010000010000000100010011;
ROM[5628] <= 32'b00000001010000000000001110010011;
ROM[5629] <= 32'b00000000100000111000001110010011;
ROM[5630] <= 32'b01000000011100010000001110110011;
ROM[5631] <= 32'b00000000011100000000001000110011;
ROM[5632] <= 32'b00000000001000000000000110110011;
ROM[5633] <= 32'b00111010100000100100000011101111;
ROM[5634] <= 32'b00000100011100000000001110010011;
ROM[5635] <= 32'b00000000011100010010000000100011;
ROM[5636] <= 32'b00000000010000010000000100010011;
ROM[5637] <= 32'b00000000000000000110001110110111;
ROM[5638] <= 32'b10000110000000111000001110010011;
ROM[5639] <= 32'b00000000111000111000001110110011;
ROM[5640] <= 32'b00000000011100010010000000100011;
ROM[5641] <= 32'b00000000010000010000000100010011;
ROM[5642] <= 32'b00000000001100010010000000100011;
ROM[5643] <= 32'b00000000010000010000000100010011;
ROM[5644] <= 32'b00000000010000010010000000100011;
ROM[5645] <= 32'b00000000010000010000000100010011;
ROM[5646] <= 32'b00000000010100010010000000100011;
ROM[5647] <= 32'b00000000010000010000000100010011;
ROM[5648] <= 32'b00000000011000010010000000100011;
ROM[5649] <= 32'b00000000010000010000000100010011;
ROM[5650] <= 32'b00000001010000000000001110010011;
ROM[5651] <= 32'b00000000100000111000001110010011;
ROM[5652] <= 32'b01000000011100010000001110110011;
ROM[5653] <= 32'b00000000011100000000001000110011;
ROM[5654] <= 32'b00000000001000000000000110110011;
ROM[5655] <= 32'b00110101000000100100000011101111;
ROM[5656] <= 32'b00000101010100000000001110010011;
ROM[5657] <= 32'b00000000011100010010000000100011;
ROM[5658] <= 32'b00000000010000010000000100010011;
ROM[5659] <= 32'b00000000000000000110001110110111;
ROM[5660] <= 32'b10001011100000111000001110010011;
ROM[5661] <= 32'b00000000111000111000001110110011;
ROM[5662] <= 32'b00000000011100010010000000100011;
ROM[5663] <= 32'b00000000010000010000000100010011;
ROM[5664] <= 32'b00000000001100010010000000100011;
ROM[5665] <= 32'b00000000010000010000000100010011;
ROM[5666] <= 32'b00000000010000010010000000100011;
ROM[5667] <= 32'b00000000010000010000000100010011;
ROM[5668] <= 32'b00000000010100010010000000100011;
ROM[5669] <= 32'b00000000010000010000000100010011;
ROM[5670] <= 32'b00000000011000010010000000100011;
ROM[5671] <= 32'b00000000010000010000000100010011;
ROM[5672] <= 32'b00000001010000000000001110010011;
ROM[5673] <= 32'b00000000100000111000001110010011;
ROM[5674] <= 32'b01000000011100010000001110110011;
ROM[5675] <= 32'b00000000011100000000001000110011;
ROM[5676] <= 32'b00000000001000000000000110110011;
ROM[5677] <= 32'b00101111100000100100000011101111;
ROM[5678] <= 32'b00000100000100000000001110010011;
ROM[5679] <= 32'b00000000011100010010000000100011;
ROM[5680] <= 32'b00000000010000010000000100010011;
ROM[5681] <= 32'b00000000000000000110001110110111;
ROM[5682] <= 32'b10010001000000111000001110010011;
ROM[5683] <= 32'b00000000111000111000001110110011;
ROM[5684] <= 32'b00000000011100010010000000100011;
ROM[5685] <= 32'b00000000010000010000000100010011;
ROM[5686] <= 32'b00000000001100010010000000100011;
ROM[5687] <= 32'b00000000010000010000000100010011;
ROM[5688] <= 32'b00000000010000010010000000100011;
ROM[5689] <= 32'b00000000010000010000000100010011;
ROM[5690] <= 32'b00000000010100010010000000100011;
ROM[5691] <= 32'b00000000010000010000000100010011;
ROM[5692] <= 32'b00000000011000010010000000100011;
ROM[5693] <= 32'b00000000010000010000000100010011;
ROM[5694] <= 32'b00000001010000000000001110010011;
ROM[5695] <= 32'b00000000100000111000001110010011;
ROM[5696] <= 32'b01000000011100010000001110110011;
ROM[5697] <= 32'b00000000011100000000001000110011;
ROM[5698] <= 32'b00000000001000000000000110110011;
ROM[5699] <= 32'b00101010000000100100000011101111;
ROM[5700] <= 32'b00000100011100000000001110010011;
ROM[5701] <= 32'b00000000011100010010000000100011;
ROM[5702] <= 32'b00000000010000010000000100010011;
ROM[5703] <= 32'b00000000000000000110001110110111;
ROM[5704] <= 32'b10010110100000111000001110010011;
ROM[5705] <= 32'b00000000111000111000001110110011;
ROM[5706] <= 32'b00000000011100010010000000100011;
ROM[5707] <= 32'b00000000010000010000000100010011;
ROM[5708] <= 32'b00000000001100010010000000100011;
ROM[5709] <= 32'b00000000010000010000000100010011;
ROM[5710] <= 32'b00000000010000010010000000100011;
ROM[5711] <= 32'b00000000010000010000000100010011;
ROM[5712] <= 32'b00000000010100010010000000100011;
ROM[5713] <= 32'b00000000010000010000000100010011;
ROM[5714] <= 32'b00000000011000010010000000100011;
ROM[5715] <= 32'b00000000010000010000000100010011;
ROM[5716] <= 32'b00000001010000000000001110010011;
ROM[5717] <= 32'b00000000100000111000001110010011;
ROM[5718] <= 32'b01000000011100010000001110110011;
ROM[5719] <= 32'b00000000011100000000001000110011;
ROM[5720] <= 32'b00000000001000000000000110110011;
ROM[5721] <= 32'b00100100100000100100000011101111;
ROM[5722] <= 32'b00000100010100000000001110010011;
ROM[5723] <= 32'b00000000011100010010000000100011;
ROM[5724] <= 32'b00000000010000010000000100010011;
ROM[5725] <= 32'b00000000000000000110001110110111;
ROM[5726] <= 32'b10011100000000111000001110010011;
ROM[5727] <= 32'b00000000111000111000001110110011;
ROM[5728] <= 32'b00000000011100010010000000100011;
ROM[5729] <= 32'b00000000010000010000000100010011;
ROM[5730] <= 32'b00000000001100010010000000100011;
ROM[5731] <= 32'b00000000010000010000000100010011;
ROM[5732] <= 32'b00000000010000010010000000100011;
ROM[5733] <= 32'b00000000010000010000000100010011;
ROM[5734] <= 32'b00000000010100010010000000100011;
ROM[5735] <= 32'b00000000010000010000000100010011;
ROM[5736] <= 32'b00000000011000010010000000100011;
ROM[5737] <= 32'b00000000010000010000000100010011;
ROM[5738] <= 32'b00000001010000000000001110010011;
ROM[5739] <= 32'b00000000100000111000001110010011;
ROM[5740] <= 32'b01000000011100010000001110110011;
ROM[5741] <= 32'b00000000011100000000001000110011;
ROM[5742] <= 32'b00000000001000000000000110110011;
ROM[5743] <= 32'b00011111000000100100000011101111;
ROM[5744] <= 32'b00000000000000011010001110000011;
ROM[5745] <= 32'b00000000011100010010000000100011;
ROM[5746] <= 32'b00000000010000010000000100010011;
ROM[5747] <= 32'b00000000001000000000001110010011;
ROM[5748] <= 32'b00000000011100010010000000100011;
ROM[5749] <= 32'b00000000010000010000000100010011;
ROM[5750] <= 32'b00000000010000000000001110010011;
ROM[5751] <= 32'b00000000011100010010000000100011;
ROM[5752] <= 32'b00000000010000010000000100010011;
ROM[5753] <= 32'b00000000000000000110001110110111;
ROM[5754] <= 32'b10100011000000111000001110010011;
ROM[5755] <= 32'b00000000111000111000001110110011;
ROM[5756] <= 32'b00000000011100010010000000100011;
ROM[5757] <= 32'b00000000010000010000000100010011;
ROM[5758] <= 32'b00000000001100010010000000100011;
ROM[5759] <= 32'b00000000010000010000000100010011;
ROM[5760] <= 32'b00000000010000010010000000100011;
ROM[5761] <= 32'b00000000010000010000000100010011;
ROM[5762] <= 32'b00000000010100010010000000100011;
ROM[5763] <= 32'b00000000010000010000000100010011;
ROM[5764] <= 32'b00000000011000010010000000100011;
ROM[5765] <= 32'b00000000010000010000000100010011;
ROM[5766] <= 32'b00000001010000000000001110010011;
ROM[5767] <= 32'b00000000100000111000001110010011;
ROM[5768] <= 32'b01000000011100010000001110110011;
ROM[5769] <= 32'b00000000011100000000001000110011;
ROM[5770] <= 32'b00000000001000000000000110110011;
ROM[5771] <= 32'b01100000000100001011000011101111;
ROM[5772] <= 32'b11111111110000010000000100010011;
ROM[5773] <= 32'b00000000000000010010001110000011;
ROM[5774] <= 32'b11111111110000010000000100010011;
ROM[5775] <= 32'b00000000000000010010010000000011;
ROM[5776] <= 32'b00000000011101000000001110110011;
ROM[5777] <= 32'b00000000011100010010000000100011;
ROM[5778] <= 32'b00000000010000010000000100010011;
ROM[5779] <= 32'b11111111110000010000000100010011;
ROM[5780] <= 32'b00000000000000010010001110000011;
ROM[5781] <= 32'b00000000000000111000001100010011;
ROM[5782] <= 32'b11111111110000010000000100010011;
ROM[5783] <= 32'b00000000000000010010001110000011;
ROM[5784] <= 32'b00000000110100110000010000110011;
ROM[5785] <= 32'b00000000011101000010000000100011;
ROM[5786] <= 32'b00000000100000000000001110010011;
ROM[5787] <= 32'b00000000011100010010000000100011;
ROM[5788] <= 32'b00000000010000010000000100010011;
ROM[5789] <= 32'b00000000000000000110001110110111;
ROM[5790] <= 32'b10101100000000111000001110010011;
ROM[5791] <= 32'b00000000111000111000001110110011;
ROM[5792] <= 32'b00000000011100010010000000100011;
ROM[5793] <= 32'b00000000010000010000000100010011;
ROM[5794] <= 32'b00000000001100010010000000100011;
ROM[5795] <= 32'b00000000010000010000000100010011;
ROM[5796] <= 32'b00000000010000010010000000100011;
ROM[5797] <= 32'b00000000010000010000000100010011;
ROM[5798] <= 32'b00000000010100010010000000100011;
ROM[5799] <= 32'b00000000010000010000000100010011;
ROM[5800] <= 32'b00000000011000010010000000100011;
ROM[5801] <= 32'b00000000010000010000000100010011;
ROM[5802] <= 32'b00000001010000000000001110010011;
ROM[5803] <= 32'b00000000010000111000001110010011;
ROM[5804] <= 32'b01000000011100010000001110110011;
ROM[5805] <= 32'b00000000011100000000001000110011;
ROM[5806] <= 32'b00000000001000000000000110110011;
ROM[5807] <= 32'b01001000000100100011000011101111;
ROM[5808] <= 32'b00000100001100000000001110010011;
ROM[5809] <= 32'b00000000011100010010000000100011;
ROM[5810] <= 32'b00000000010000010000000100010011;
ROM[5811] <= 32'b00000000000000000110001110110111;
ROM[5812] <= 32'b10110001100000111000001110010011;
ROM[5813] <= 32'b00000000111000111000001110110011;
ROM[5814] <= 32'b00000000011100010010000000100011;
ROM[5815] <= 32'b00000000010000010000000100010011;
ROM[5816] <= 32'b00000000001100010010000000100011;
ROM[5817] <= 32'b00000000010000010000000100010011;
ROM[5818] <= 32'b00000000010000010010000000100011;
ROM[5819] <= 32'b00000000010000010000000100010011;
ROM[5820] <= 32'b00000000010100010010000000100011;
ROM[5821] <= 32'b00000000010000010000000100010011;
ROM[5822] <= 32'b00000000011000010010000000100011;
ROM[5823] <= 32'b00000000010000010000000100010011;
ROM[5824] <= 32'b00000001010000000000001110010011;
ROM[5825] <= 32'b00000000100000111000001110010011;
ROM[5826] <= 32'b01000000011100010000001110110011;
ROM[5827] <= 32'b00000000011100000000001000110011;
ROM[5828] <= 32'b00000000001000000000000110110011;
ROM[5829] <= 32'b00001001100000100100000011101111;
ROM[5830] <= 32'b00000100111100000000001110010011;
ROM[5831] <= 32'b00000000011100010010000000100011;
ROM[5832] <= 32'b00000000010000010000000100010011;
ROM[5833] <= 32'b00000000000000000110001110110111;
ROM[5834] <= 32'b10110111000000111000001110010011;
ROM[5835] <= 32'b00000000111000111000001110110011;
ROM[5836] <= 32'b00000000011100010010000000100011;
ROM[5837] <= 32'b00000000010000010000000100010011;
ROM[5838] <= 32'b00000000001100010010000000100011;
ROM[5839] <= 32'b00000000010000010000000100010011;
ROM[5840] <= 32'b00000000010000010010000000100011;
ROM[5841] <= 32'b00000000010000010000000100010011;
ROM[5842] <= 32'b00000000010100010010000000100011;
ROM[5843] <= 32'b00000000010000010000000100010011;
ROM[5844] <= 32'b00000000011000010010000000100011;
ROM[5845] <= 32'b00000000010000010000000100010011;
ROM[5846] <= 32'b00000001010000000000001110010011;
ROM[5847] <= 32'b00000000100000111000001110010011;
ROM[5848] <= 32'b01000000011100010000001110110011;
ROM[5849] <= 32'b00000000011100000000001000110011;
ROM[5850] <= 32'b00000000001000000000000110110011;
ROM[5851] <= 32'b00000100000000100100000011101111;
ROM[5852] <= 32'b00000100110100000000001110010011;
ROM[5853] <= 32'b00000000011100010010000000100011;
ROM[5854] <= 32'b00000000010000010000000100010011;
ROM[5855] <= 32'b00000000000000000110001110110111;
ROM[5856] <= 32'b10111100100000111000001110010011;
ROM[5857] <= 32'b00000000111000111000001110110011;
ROM[5858] <= 32'b00000000011100010010000000100011;
ROM[5859] <= 32'b00000000010000010000000100010011;
ROM[5860] <= 32'b00000000001100010010000000100011;
ROM[5861] <= 32'b00000000010000010000000100010011;
ROM[5862] <= 32'b00000000010000010010000000100011;
ROM[5863] <= 32'b00000000010000010000000100010011;
ROM[5864] <= 32'b00000000010100010010000000100011;
ROM[5865] <= 32'b00000000010000010000000100010011;
ROM[5866] <= 32'b00000000011000010010000000100011;
ROM[5867] <= 32'b00000000010000010000000100010011;
ROM[5868] <= 32'b00000001010000000000001110010011;
ROM[5869] <= 32'b00000000100000111000001110010011;
ROM[5870] <= 32'b01000000011100010000001110110011;
ROM[5871] <= 32'b00000000011100000000001000110011;
ROM[5872] <= 32'b00000000001000000000000110110011;
ROM[5873] <= 32'b01111110100100100011000011101111;
ROM[5874] <= 32'b00000101000000000000001110010011;
ROM[5875] <= 32'b00000000011100010010000000100011;
ROM[5876] <= 32'b00000000010000010000000100010011;
ROM[5877] <= 32'b00000000000000000110001110110111;
ROM[5878] <= 32'b11000010000000111000001110010011;
ROM[5879] <= 32'b00000000111000111000001110110011;
ROM[5880] <= 32'b00000000011100010010000000100011;
ROM[5881] <= 32'b00000000010000010000000100010011;
ROM[5882] <= 32'b00000000001100010010000000100011;
ROM[5883] <= 32'b00000000010000010000000100010011;
ROM[5884] <= 32'b00000000010000010010000000100011;
ROM[5885] <= 32'b00000000010000010000000100010011;
ROM[5886] <= 32'b00000000010100010010000000100011;
ROM[5887] <= 32'b00000000010000010000000100010011;
ROM[5888] <= 32'b00000000011000010010000000100011;
ROM[5889] <= 32'b00000000010000010000000100010011;
ROM[5890] <= 32'b00000001010000000000001110010011;
ROM[5891] <= 32'b00000000100000111000001110010011;
ROM[5892] <= 32'b01000000011100010000001110110011;
ROM[5893] <= 32'b00000000011100000000001000110011;
ROM[5894] <= 32'b00000000001000000000000110110011;
ROM[5895] <= 32'b01111001000100100011000011101111;
ROM[5896] <= 32'b00000100100100000000001110010011;
ROM[5897] <= 32'b00000000011100010010000000100011;
ROM[5898] <= 32'b00000000010000010000000100010011;
ROM[5899] <= 32'b00000000000000000110001110110111;
ROM[5900] <= 32'b11000111100000111000001110010011;
ROM[5901] <= 32'b00000000111000111000001110110011;
ROM[5902] <= 32'b00000000011100010010000000100011;
ROM[5903] <= 32'b00000000010000010000000100010011;
ROM[5904] <= 32'b00000000001100010010000000100011;
ROM[5905] <= 32'b00000000010000010000000100010011;
ROM[5906] <= 32'b00000000010000010010000000100011;
ROM[5907] <= 32'b00000000010000010000000100010011;
ROM[5908] <= 32'b00000000010100010010000000100011;
ROM[5909] <= 32'b00000000010000010000000100010011;
ROM[5910] <= 32'b00000000011000010010000000100011;
ROM[5911] <= 32'b00000000010000010000000100010011;
ROM[5912] <= 32'b00000001010000000000001110010011;
ROM[5913] <= 32'b00000000100000111000001110010011;
ROM[5914] <= 32'b01000000011100010000001110110011;
ROM[5915] <= 32'b00000000011100000000001000110011;
ROM[5916] <= 32'b00000000001000000000000110110011;
ROM[5917] <= 32'b01110011100100100011000011101111;
ROM[5918] <= 32'b00000100110000000000001110010011;
ROM[5919] <= 32'b00000000011100010010000000100011;
ROM[5920] <= 32'b00000000010000010000000100010011;
ROM[5921] <= 32'b00000000000000000110001110110111;
ROM[5922] <= 32'b11001101000000111000001110010011;
ROM[5923] <= 32'b00000000111000111000001110110011;
ROM[5924] <= 32'b00000000011100010010000000100011;
ROM[5925] <= 32'b00000000010000010000000100010011;
ROM[5926] <= 32'b00000000001100010010000000100011;
ROM[5927] <= 32'b00000000010000010000000100010011;
ROM[5928] <= 32'b00000000010000010010000000100011;
ROM[5929] <= 32'b00000000010000010000000100010011;
ROM[5930] <= 32'b00000000010100010010000000100011;
ROM[5931] <= 32'b00000000010000010000000100010011;
ROM[5932] <= 32'b00000000011000010010000000100011;
ROM[5933] <= 32'b00000000010000010000000100010011;
ROM[5934] <= 32'b00000001010000000000001110010011;
ROM[5935] <= 32'b00000000100000111000001110010011;
ROM[5936] <= 32'b01000000011100010000001110110011;
ROM[5937] <= 32'b00000000011100000000001000110011;
ROM[5938] <= 32'b00000000001000000000000110110011;
ROM[5939] <= 32'b01101110000100100011000011101111;
ROM[5940] <= 32'b00000100010100000000001110010011;
ROM[5941] <= 32'b00000000011100010010000000100011;
ROM[5942] <= 32'b00000000010000010000000100010011;
ROM[5943] <= 32'b00000000000000000110001110110111;
ROM[5944] <= 32'b11010010100000111000001110010011;
ROM[5945] <= 32'b00000000111000111000001110110011;
ROM[5946] <= 32'b00000000011100010010000000100011;
ROM[5947] <= 32'b00000000010000010000000100010011;
ROM[5948] <= 32'b00000000001100010010000000100011;
ROM[5949] <= 32'b00000000010000010000000100010011;
ROM[5950] <= 32'b00000000010000010010000000100011;
ROM[5951] <= 32'b00000000010000010000000100010011;
ROM[5952] <= 32'b00000000010100010010000000100011;
ROM[5953] <= 32'b00000000010000010000000100010011;
ROM[5954] <= 32'b00000000011000010010000000100011;
ROM[5955] <= 32'b00000000010000010000000100010011;
ROM[5956] <= 32'b00000001010000000000001110010011;
ROM[5957] <= 32'b00000000100000111000001110010011;
ROM[5958] <= 32'b01000000011100010000001110110011;
ROM[5959] <= 32'b00000000011100000000001000110011;
ROM[5960] <= 32'b00000000001000000000000110110011;
ROM[5961] <= 32'b01101000100100100011000011101111;
ROM[5962] <= 32'b00000101001000000000001110010011;
ROM[5963] <= 32'b00000000011100010010000000100011;
ROM[5964] <= 32'b00000000010000010000000100010011;
ROM[5965] <= 32'b00000000000000000110001110110111;
ROM[5966] <= 32'b11011000000000111000001110010011;
ROM[5967] <= 32'b00000000111000111000001110110011;
ROM[5968] <= 32'b00000000011100010010000000100011;
ROM[5969] <= 32'b00000000010000010000000100010011;
ROM[5970] <= 32'b00000000001100010010000000100011;
ROM[5971] <= 32'b00000000010000010000000100010011;
ROM[5972] <= 32'b00000000010000010010000000100011;
ROM[5973] <= 32'b00000000010000010000000100010011;
ROM[5974] <= 32'b00000000010100010010000000100011;
ROM[5975] <= 32'b00000000010000010000000100010011;
ROM[5976] <= 32'b00000000011000010010000000100011;
ROM[5977] <= 32'b00000000010000010000000100010011;
ROM[5978] <= 32'b00000001010000000000001110010011;
ROM[5979] <= 32'b00000000100000111000001110010011;
ROM[5980] <= 32'b01000000011100010000001110110011;
ROM[5981] <= 32'b00000000011100000000001000110011;
ROM[5982] <= 32'b00000000001000000000000110110011;
ROM[5983] <= 32'b01100011000100100011000011101111;
ROM[5984] <= 32'b00000000000000011010001110000011;
ROM[5985] <= 32'b00000000011100010010000000100011;
ROM[5986] <= 32'b00000000010000010000000100010011;
ROM[5987] <= 32'b00000000001100000000001110010011;
ROM[5988] <= 32'b00000000011100010010000000100011;
ROM[5989] <= 32'b00000000010000010000000100010011;
ROM[5990] <= 32'b00000000010000000000001110010011;
ROM[5991] <= 32'b00000000011100010010000000100011;
ROM[5992] <= 32'b00000000010000010000000100010011;
ROM[5993] <= 32'b00000000000000000110001110110111;
ROM[5994] <= 32'b11011111000000111000001110010011;
ROM[5995] <= 32'b00000000111000111000001110110011;
ROM[5996] <= 32'b00000000011100010010000000100011;
ROM[5997] <= 32'b00000000010000010000000100010011;
ROM[5998] <= 32'b00000000001100010010000000100011;
ROM[5999] <= 32'b00000000010000010000000100010011;
ROM[6000] <= 32'b00000000010000010010000000100011;
ROM[6001] <= 32'b00000000010000010000000100010011;
ROM[6002] <= 32'b00000000010100010010000000100011;
ROM[6003] <= 32'b00000000010000010000000100010011;
ROM[6004] <= 32'b00000000011000010010000000100011;
ROM[6005] <= 32'b00000000010000010000000100010011;
ROM[6006] <= 32'b00000001010000000000001110010011;
ROM[6007] <= 32'b00000000100000111000001110010011;
ROM[6008] <= 32'b01000000011100010000001110110011;
ROM[6009] <= 32'b00000000011100000000001000110011;
ROM[6010] <= 32'b00000000001000000000000110110011;
ROM[6011] <= 32'b00100100000100001011000011101111;
ROM[6012] <= 32'b11111111110000010000000100010011;
ROM[6013] <= 32'b00000000000000010010001110000011;
ROM[6014] <= 32'b11111111110000010000000100010011;
ROM[6015] <= 32'b00000000000000010010010000000011;
ROM[6016] <= 32'b00000000011101000000001110110011;
ROM[6017] <= 32'b00000000011100010010000000100011;
ROM[6018] <= 32'b00000000010000010000000100010011;
ROM[6019] <= 32'b11111111110000010000000100010011;
ROM[6020] <= 32'b00000000000000010010001110000011;
ROM[6021] <= 32'b00000000000000111000001100010011;
ROM[6022] <= 32'b11111111110000010000000100010011;
ROM[6023] <= 32'b00000000000000010010001110000011;
ROM[6024] <= 32'b00000000110100110000010000110011;
ROM[6025] <= 32'b00000000011101000010000000100011;
ROM[6026] <= 32'b00000000011100000000001110010011;
ROM[6027] <= 32'b00000000011100010010000000100011;
ROM[6028] <= 32'b00000000010000010000000100010011;
ROM[6029] <= 32'b00000000000000000110001110110111;
ROM[6030] <= 32'b11101000000000111000001110010011;
ROM[6031] <= 32'b00000000111000111000001110110011;
ROM[6032] <= 32'b00000000011100010010000000100011;
ROM[6033] <= 32'b00000000010000010000000100010011;
ROM[6034] <= 32'b00000000001100010010000000100011;
ROM[6035] <= 32'b00000000010000010000000100010011;
ROM[6036] <= 32'b00000000010000010010000000100011;
ROM[6037] <= 32'b00000000010000010000000100010011;
ROM[6038] <= 32'b00000000010100010010000000100011;
ROM[6039] <= 32'b00000000010000010000000100010011;
ROM[6040] <= 32'b00000000011000010010000000100011;
ROM[6041] <= 32'b00000000010000010000000100010011;
ROM[6042] <= 32'b00000001010000000000001110010011;
ROM[6043] <= 32'b00000000010000111000001110010011;
ROM[6044] <= 32'b01000000011100010000001110110011;
ROM[6045] <= 32'b00000000011100000000001000110011;
ROM[6046] <= 32'b00000000001000000000000110110011;
ROM[6047] <= 32'b00001100000100100011000011101111;
ROM[6048] <= 32'b00000101011000000000001110010011;
ROM[6049] <= 32'b00000000011100010010000000100011;
ROM[6050] <= 32'b00000000010000010000000100010011;
ROM[6051] <= 32'b00000000000000000110001110110111;
ROM[6052] <= 32'b11101101100000111000001110010011;
ROM[6053] <= 32'b00000000111000111000001110110011;
ROM[6054] <= 32'b00000000011100010010000000100011;
ROM[6055] <= 32'b00000000010000010000000100010011;
ROM[6056] <= 32'b00000000001100010010000000100011;
ROM[6057] <= 32'b00000000010000010000000100010011;
ROM[6058] <= 32'b00000000010000010010000000100011;
ROM[6059] <= 32'b00000000010000010000000100010011;
ROM[6060] <= 32'b00000000010100010010000000100011;
ROM[6061] <= 32'b00000000010000010000000100010011;
ROM[6062] <= 32'b00000000011000010010000000100011;
ROM[6063] <= 32'b00000000010000010000000100010011;
ROM[6064] <= 32'b00000001010000000000001110010011;
ROM[6065] <= 32'b00000000100000111000001110010011;
ROM[6066] <= 32'b01000000011100010000001110110011;
ROM[6067] <= 32'b00000000011100000000001000110011;
ROM[6068] <= 32'b00000000001000000000000110110011;
ROM[6069] <= 32'b01001101100100100011000011101111;
ROM[6070] <= 32'b00000100100100000000001110010011;
ROM[6071] <= 32'b00000000011100010010000000100011;
ROM[6072] <= 32'b00000000010000010000000100010011;
ROM[6073] <= 32'b00000000000000000110001110110111;
ROM[6074] <= 32'b11110011000000111000001110010011;
ROM[6075] <= 32'b00000000111000111000001110110011;
ROM[6076] <= 32'b00000000011100010010000000100011;
ROM[6077] <= 32'b00000000010000010000000100010011;
ROM[6078] <= 32'b00000000001100010010000000100011;
ROM[6079] <= 32'b00000000010000010000000100010011;
ROM[6080] <= 32'b00000000010000010010000000100011;
ROM[6081] <= 32'b00000000010000010000000100010011;
ROM[6082] <= 32'b00000000010100010010000000100011;
ROM[6083] <= 32'b00000000010000010000000100010011;
ROM[6084] <= 32'b00000000011000010010000000100011;
ROM[6085] <= 32'b00000000010000010000000100010011;
ROM[6086] <= 32'b00000001010000000000001110010011;
ROM[6087] <= 32'b00000000100000111000001110010011;
ROM[6088] <= 32'b01000000011100010000001110110011;
ROM[6089] <= 32'b00000000011100000000001000110011;
ROM[6090] <= 32'b00000000001000000000000110110011;
ROM[6091] <= 32'b01001000000100100011000011101111;
ROM[6092] <= 32'b00000101001000000000001110010011;
ROM[6093] <= 32'b00000000011100010010000000100011;
ROM[6094] <= 32'b00000000010000010000000100010011;
ROM[6095] <= 32'b00000000000000000110001110110111;
ROM[6096] <= 32'b11111000100000111000001110010011;
ROM[6097] <= 32'b00000000111000111000001110110011;
ROM[6098] <= 32'b00000000011100010010000000100011;
ROM[6099] <= 32'b00000000010000010000000100010011;
ROM[6100] <= 32'b00000000001100010010000000100011;
ROM[6101] <= 32'b00000000010000010000000100010011;
ROM[6102] <= 32'b00000000010000010010000000100011;
ROM[6103] <= 32'b00000000010000010000000100010011;
ROM[6104] <= 32'b00000000010100010010000000100011;
ROM[6105] <= 32'b00000000010000010000000100010011;
ROM[6106] <= 32'b00000000011000010010000000100011;
ROM[6107] <= 32'b00000000010000010000000100010011;
ROM[6108] <= 32'b00000001010000000000001110010011;
ROM[6109] <= 32'b00000000100000111000001110010011;
ROM[6110] <= 32'b01000000011100010000001110110011;
ROM[6111] <= 32'b00000000011100000000001000110011;
ROM[6112] <= 32'b00000000001000000000000110110011;
ROM[6113] <= 32'b01000010100100100011000011101111;
ROM[6114] <= 32'b00000101010000000000001110010011;
ROM[6115] <= 32'b00000000011100010010000000100011;
ROM[6116] <= 32'b00000000010000010000000100010011;
ROM[6117] <= 32'b00000000000000000110001110110111;
ROM[6118] <= 32'b11111110000000111000001110010011;
ROM[6119] <= 32'b00000000111000111000001110110011;
ROM[6120] <= 32'b00000000011100010010000000100011;
ROM[6121] <= 32'b00000000010000010000000100010011;
ROM[6122] <= 32'b00000000001100010010000000100011;
ROM[6123] <= 32'b00000000010000010000000100010011;
ROM[6124] <= 32'b00000000010000010010000000100011;
ROM[6125] <= 32'b00000000010000010000000100010011;
ROM[6126] <= 32'b00000000010100010010000000100011;
ROM[6127] <= 32'b00000000010000010000000100010011;
ROM[6128] <= 32'b00000000011000010010000000100011;
ROM[6129] <= 32'b00000000010000010000000100010011;
ROM[6130] <= 32'b00000001010000000000001110010011;
ROM[6131] <= 32'b00000000100000111000001110010011;
ROM[6132] <= 32'b01000000011100010000001110110011;
ROM[6133] <= 32'b00000000011100000000001000110011;
ROM[6134] <= 32'b00000000001000000000000110110011;
ROM[6135] <= 32'b00111101000100100011000011101111;
ROM[6136] <= 32'b00000101010100000000001110010011;
ROM[6137] <= 32'b00000000011100010010000000100011;
ROM[6138] <= 32'b00000000010000010000000100010011;
ROM[6139] <= 32'b00000000000000000110001110110111;
ROM[6140] <= 32'b00000011100000111000001110010011;
ROM[6141] <= 32'b00000000111000111000001110110011;
ROM[6142] <= 32'b00000000011100010010000000100011;
ROM[6143] <= 32'b00000000010000010000000100010011;
ROM[6144] <= 32'b00000000001100010010000000100011;
ROM[6145] <= 32'b00000000010000010000000100010011;
ROM[6146] <= 32'b00000000010000010010000000100011;
ROM[6147] <= 32'b00000000010000010000000100010011;
ROM[6148] <= 32'b00000000010100010010000000100011;
ROM[6149] <= 32'b00000000010000010000000100010011;
ROM[6150] <= 32'b00000000011000010010000000100011;
ROM[6151] <= 32'b00000000010000010000000100010011;
ROM[6152] <= 32'b00000001010000000000001110010011;
ROM[6153] <= 32'b00000000100000111000001110010011;
ROM[6154] <= 32'b01000000011100010000001110110011;
ROM[6155] <= 32'b00000000011100000000001000110011;
ROM[6156] <= 32'b00000000001000000000000110110011;
ROM[6157] <= 32'b00110111100100100011000011101111;
ROM[6158] <= 32'b00000100000100000000001110010011;
ROM[6159] <= 32'b00000000011100010010000000100011;
ROM[6160] <= 32'b00000000010000010000000100010011;
ROM[6161] <= 32'b00000000000000000110001110110111;
ROM[6162] <= 32'b00001001000000111000001110010011;
ROM[6163] <= 32'b00000000111000111000001110110011;
ROM[6164] <= 32'b00000000011100010010000000100011;
ROM[6165] <= 32'b00000000010000010000000100010011;
ROM[6166] <= 32'b00000000001100010010000000100011;
ROM[6167] <= 32'b00000000010000010000000100010011;
ROM[6168] <= 32'b00000000010000010010000000100011;
ROM[6169] <= 32'b00000000010000010000000100010011;
ROM[6170] <= 32'b00000000010100010010000000100011;
ROM[6171] <= 32'b00000000010000010000000100010011;
ROM[6172] <= 32'b00000000011000010010000000100011;
ROM[6173] <= 32'b00000000010000010000000100010011;
ROM[6174] <= 32'b00000001010000000000001110010011;
ROM[6175] <= 32'b00000000100000111000001110010011;
ROM[6176] <= 32'b01000000011100010000001110110011;
ROM[6177] <= 32'b00000000011100000000001000110011;
ROM[6178] <= 32'b00000000001000000000000110110011;
ROM[6179] <= 32'b00110010000100100011000011101111;
ROM[6180] <= 32'b00000100110000000000001110010011;
ROM[6181] <= 32'b00000000011100010010000000100011;
ROM[6182] <= 32'b00000000010000010000000100010011;
ROM[6183] <= 32'b00000000000000000110001110110111;
ROM[6184] <= 32'b00001110100000111000001110010011;
ROM[6185] <= 32'b00000000111000111000001110110011;
ROM[6186] <= 32'b00000000011100010010000000100011;
ROM[6187] <= 32'b00000000010000010000000100010011;
ROM[6188] <= 32'b00000000001100010010000000100011;
ROM[6189] <= 32'b00000000010000010000000100010011;
ROM[6190] <= 32'b00000000010000010010000000100011;
ROM[6191] <= 32'b00000000010000010000000100010011;
ROM[6192] <= 32'b00000000010100010010000000100011;
ROM[6193] <= 32'b00000000010000010000000100010011;
ROM[6194] <= 32'b00000000011000010010000000100011;
ROM[6195] <= 32'b00000000010000010000000100010011;
ROM[6196] <= 32'b00000001010000000000001110010011;
ROM[6197] <= 32'b00000000100000111000001110010011;
ROM[6198] <= 32'b01000000011100010000001110110011;
ROM[6199] <= 32'b00000000011100000000001000110011;
ROM[6200] <= 32'b00000000001000000000000110110011;
ROM[6201] <= 32'b00101100100100100011000011101111;
ROM[6202] <= 32'b00000000000000011010001110000011;
ROM[6203] <= 32'b00000000011100010010000000100011;
ROM[6204] <= 32'b00000000010000010000000100010011;
ROM[6205] <= 32'b00000000010000000000001110010011;
ROM[6206] <= 32'b00000000011100010010000000100011;
ROM[6207] <= 32'b00000000010000010000000100010011;
ROM[6208] <= 32'b00000000010000000000001110010011;
ROM[6209] <= 32'b00000000011100010010000000100011;
ROM[6210] <= 32'b00000000010000010000000100010011;
ROM[6211] <= 32'b00000000000000000110001110110111;
ROM[6212] <= 32'b00010101100000111000001110010011;
ROM[6213] <= 32'b00000000111000111000001110110011;
ROM[6214] <= 32'b00000000011100010010000000100011;
ROM[6215] <= 32'b00000000010000010000000100010011;
ROM[6216] <= 32'b00000000001100010010000000100011;
ROM[6217] <= 32'b00000000010000010000000100010011;
ROM[6218] <= 32'b00000000010000010010000000100011;
ROM[6219] <= 32'b00000000010000010000000100010011;
ROM[6220] <= 32'b00000000010100010010000000100011;
ROM[6221] <= 32'b00000000010000010000000100010011;
ROM[6222] <= 32'b00000000011000010010000000100011;
ROM[6223] <= 32'b00000000010000010000000100010011;
ROM[6224] <= 32'b00000001010000000000001110010011;
ROM[6225] <= 32'b00000000100000111000001110010011;
ROM[6226] <= 32'b01000000011100010000001110110011;
ROM[6227] <= 32'b00000000011100000000001000110011;
ROM[6228] <= 32'b00000000001000000000000110110011;
ROM[6229] <= 32'b01101101100000001011000011101111;
ROM[6230] <= 32'b11111111110000010000000100010011;
ROM[6231] <= 32'b00000000000000010010001110000011;
ROM[6232] <= 32'b11111111110000010000000100010011;
ROM[6233] <= 32'b00000000000000010010010000000011;
ROM[6234] <= 32'b00000000011101000000001110110011;
ROM[6235] <= 32'b00000000011100010010000000100011;
ROM[6236] <= 32'b00000000010000010000000100010011;
ROM[6237] <= 32'b11111111110000010000000100010011;
ROM[6238] <= 32'b00000000000000010010001110000011;
ROM[6239] <= 32'b00000000000000111000001100010011;
ROM[6240] <= 32'b11111111110000010000000100010011;
ROM[6241] <= 32'b00000000000000010010001110000011;
ROM[6242] <= 32'b00000000110100110000010000110011;
ROM[6243] <= 32'b00000000011101000010000000100011;
ROM[6244] <= 32'b00000000010100000000001110010011;
ROM[6245] <= 32'b00000000011100010010000000100011;
ROM[6246] <= 32'b00000000010000010000000100010011;
ROM[6247] <= 32'b00000000000000000110001110110111;
ROM[6248] <= 32'b00011110100000111000001110010011;
ROM[6249] <= 32'b00000000111000111000001110110011;
ROM[6250] <= 32'b00000000011100010010000000100011;
ROM[6251] <= 32'b00000000010000010000000100010011;
ROM[6252] <= 32'b00000000001100010010000000100011;
ROM[6253] <= 32'b00000000010000010000000100010011;
ROM[6254] <= 32'b00000000010000010010000000100011;
ROM[6255] <= 32'b00000000010000010000000100010011;
ROM[6256] <= 32'b00000000010100010010000000100011;
ROM[6257] <= 32'b00000000010000010000000100010011;
ROM[6258] <= 32'b00000000011000010010000000100011;
ROM[6259] <= 32'b00000000010000010000000100010011;
ROM[6260] <= 32'b00000001010000000000001110010011;
ROM[6261] <= 32'b00000000010000111000001110010011;
ROM[6262] <= 32'b01000000011100010000001110110011;
ROM[6263] <= 32'b00000000011100000000001000110011;
ROM[6264] <= 32'b00000000001000000000000110110011;
ROM[6265] <= 32'b11101001110111111001000011101111;
ROM[6266] <= 32'b11111111110000010000000100010011;
ROM[6267] <= 32'b00000000000000010010001110000011;
ROM[6268] <= 32'b00000010011100011010111000100011;
ROM[6269] <= 32'b00000000010000000000001110010011;
ROM[6270] <= 32'b00000000011100010010000000100011;
ROM[6271] <= 32'b00000000010000010000000100010011;
ROM[6272] <= 32'b00000011110000011010001110000011;
ROM[6273] <= 32'b00000000011100010010000000100011;
ROM[6274] <= 32'b00000000010000010000000100010011;
ROM[6275] <= 32'b00000000000000000000001110010011;
ROM[6276] <= 32'b00000000011100010010000000100011;
ROM[6277] <= 32'b00000000010000010000000100010011;
ROM[6278] <= 32'b00000000010000000000001110010011;
ROM[6279] <= 32'b00000000011100010010000000100011;
ROM[6280] <= 32'b00000000010000010000000100010011;
ROM[6281] <= 32'b00000000000000000110001110110111;
ROM[6282] <= 32'b00100111000000111000001110010011;
ROM[6283] <= 32'b00000000111000111000001110110011;
ROM[6284] <= 32'b00000000011100010010000000100011;
ROM[6285] <= 32'b00000000010000010000000100010011;
ROM[6286] <= 32'b00000000001100010010000000100011;
ROM[6287] <= 32'b00000000010000010000000100010011;
ROM[6288] <= 32'b00000000010000010010000000100011;
ROM[6289] <= 32'b00000000010000010000000100010011;
ROM[6290] <= 32'b00000000010100010010000000100011;
ROM[6291] <= 32'b00000000010000010000000100010011;
ROM[6292] <= 32'b00000000011000010010000000100011;
ROM[6293] <= 32'b00000000010000010000000100010011;
ROM[6294] <= 32'b00000001010000000000001110010011;
ROM[6295] <= 32'b00000000100000111000001110010011;
ROM[6296] <= 32'b01000000011100010000001110110011;
ROM[6297] <= 32'b00000000011100000000001000110011;
ROM[6298] <= 32'b00000000001000000000000110110011;
ROM[6299] <= 32'b01011100000000001011000011101111;
ROM[6300] <= 32'b11111111110000010000000100010011;
ROM[6301] <= 32'b00000000000000010010001110000011;
ROM[6302] <= 32'b11111111110000010000000100010011;
ROM[6303] <= 32'b00000000000000010010010000000011;
ROM[6304] <= 32'b00000000011101000000001110110011;
ROM[6305] <= 32'b00000000011100010010000000100011;
ROM[6306] <= 32'b00000000010000010000000100010011;
ROM[6307] <= 32'b11111111110000010000000100010011;
ROM[6308] <= 32'b00000000000000010010001110000011;
ROM[6309] <= 32'b00000000000000111000001100010011;
ROM[6310] <= 32'b11111111110000010000000100010011;
ROM[6311] <= 32'b00000000000000010010001110000011;
ROM[6312] <= 32'b00000000110100110000010000110011;
ROM[6313] <= 32'b00000000011101000010000000100011;
ROM[6314] <= 32'b00000000101100000000001110010011;
ROM[6315] <= 32'b00000000011100010010000000100011;
ROM[6316] <= 32'b00000000010000010000000100010011;
ROM[6317] <= 32'b00000011110000011010001110000011;
ROM[6318] <= 32'b00000000011100010010000000100011;
ROM[6319] <= 32'b00000000010000010000000100010011;
ROM[6320] <= 32'b00000000000100000000001110010011;
ROM[6321] <= 32'b00000000011100010010000000100011;
ROM[6322] <= 32'b00000000010000010000000100010011;
ROM[6323] <= 32'b00000000010000000000001110010011;
ROM[6324] <= 32'b00000000011100010010000000100011;
ROM[6325] <= 32'b00000000010000010000000100010011;
ROM[6326] <= 32'b00000000000000000110001110110111;
ROM[6327] <= 32'b00110010010000111000001110010011;
ROM[6328] <= 32'b00000000111000111000001110110011;
ROM[6329] <= 32'b00000000011100010010000000100011;
ROM[6330] <= 32'b00000000010000010000000100010011;
ROM[6331] <= 32'b00000000001100010010000000100011;
ROM[6332] <= 32'b00000000010000010000000100010011;
ROM[6333] <= 32'b00000000010000010010000000100011;
ROM[6334] <= 32'b00000000010000010000000100010011;
ROM[6335] <= 32'b00000000010100010010000000100011;
ROM[6336] <= 32'b00000000010000010000000100010011;
ROM[6337] <= 32'b00000000011000010010000000100011;
ROM[6338] <= 32'b00000000010000010000000100010011;
ROM[6339] <= 32'b00000001010000000000001110010011;
ROM[6340] <= 32'b00000000100000111000001110010011;
ROM[6341] <= 32'b01000000011100010000001110110011;
ROM[6342] <= 32'b00000000011100000000001000110011;
ROM[6343] <= 32'b00000000001000000000000110110011;
ROM[6344] <= 32'b01010000110000001011000011101111;
ROM[6345] <= 32'b11111111110000010000000100010011;
ROM[6346] <= 32'b00000000000000010010001110000011;
ROM[6347] <= 32'b11111111110000010000000100010011;
ROM[6348] <= 32'b00000000000000010010010000000011;
ROM[6349] <= 32'b00000000011101000000001110110011;
ROM[6350] <= 32'b00000000011100010010000000100011;
ROM[6351] <= 32'b00000000010000010000000100010011;
ROM[6352] <= 32'b11111111110000010000000100010011;
ROM[6353] <= 32'b00000000000000010010001110000011;
ROM[6354] <= 32'b00000000000000111000001100010011;
ROM[6355] <= 32'b11111111110000010000000100010011;
ROM[6356] <= 32'b00000000000000010010001110000011;
ROM[6357] <= 32'b00000000110100110000010000110011;
ROM[6358] <= 32'b00000000011101000010000000100011;
ROM[6359] <= 32'b00000000100000000000001110010011;
ROM[6360] <= 32'b00000000011100010010000000100011;
ROM[6361] <= 32'b00000000010000010000000100010011;
ROM[6362] <= 32'b00000011110000011010001110000011;
ROM[6363] <= 32'b00000000011100010010000000100011;
ROM[6364] <= 32'b00000000010000010000000100010011;
ROM[6365] <= 32'b00000000001000000000001110010011;
ROM[6366] <= 32'b00000000011100010010000000100011;
ROM[6367] <= 32'b00000000010000010000000100010011;
ROM[6368] <= 32'b00000000010000000000001110010011;
ROM[6369] <= 32'b00000000011100010010000000100011;
ROM[6370] <= 32'b00000000010000010000000100010011;
ROM[6371] <= 32'b00000000000000000110001110110111;
ROM[6372] <= 32'b00111101100000111000001110010011;
ROM[6373] <= 32'b00000000111000111000001110110011;
ROM[6374] <= 32'b00000000011100010010000000100011;
ROM[6375] <= 32'b00000000010000010000000100010011;
ROM[6376] <= 32'b00000000001100010010000000100011;
ROM[6377] <= 32'b00000000010000010000000100010011;
ROM[6378] <= 32'b00000000010000010010000000100011;
ROM[6379] <= 32'b00000000010000010000000100010011;
ROM[6380] <= 32'b00000000010100010010000000100011;
ROM[6381] <= 32'b00000000010000010000000100010011;
ROM[6382] <= 32'b00000000011000010010000000100011;
ROM[6383] <= 32'b00000000010000010000000100010011;
ROM[6384] <= 32'b00000001010000000000001110010011;
ROM[6385] <= 32'b00000000100000111000001110010011;
ROM[6386] <= 32'b01000000011100010000001110110011;
ROM[6387] <= 32'b00000000011100000000001000110011;
ROM[6388] <= 32'b00000000001000000000000110110011;
ROM[6389] <= 32'b01000101100000001011000011101111;
ROM[6390] <= 32'b11111111110000010000000100010011;
ROM[6391] <= 32'b00000000000000010010001110000011;
ROM[6392] <= 32'b11111111110000010000000100010011;
ROM[6393] <= 32'b00000000000000010010010000000011;
ROM[6394] <= 32'b00000000011101000000001110110011;
ROM[6395] <= 32'b00000000011100010010000000100011;
ROM[6396] <= 32'b00000000010000010000000100010011;
ROM[6397] <= 32'b11111111110000010000000100010011;
ROM[6398] <= 32'b00000000000000010010001110000011;
ROM[6399] <= 32'b00000000000000111000001100010011;
ROM[6400] <= 32'b11111111110000010000000100010011;
ROM[6401] <= 32'b00000000000000010010001110000011;
ROM[6402] <= 32'b00000000110100110000010000110011;
ROM[6403] <= 32'b00000000011101000010000000100011;
ROM[6404] <= 32'b00000000100000000000001110010011;
ROM[6405] <= 32'b00000000011100010010000000100011;
ROM[6406] <= 32'b00000000010000010000000100010011;
ROM[6407] <= 32'b00000011110000011010001110000011;
ROM[6408] <= 32'b00000000011100010010000000100011;
ROM[6409] <= 32'b00000000010000010000000100010011;
ROM[6410] <= 32'b00000000001100000000001110010011;
ROM[6411] <= 32'b00000000011100010010000000100011;
ROM[6412] <= 32'b00000000010000010000000100010011;
ROM[6413] <= 32'b00000000010000000000001110010011;
ROM[6414] <= 32'b00000000011100010010000000100011;
ROM[6415] <= 32'b00000000010000010000000100010011;
ROM[6416] <= 32'b00000000000000000110001110110111;
ROM[6417] <= 32'b01001000110000111000001110010011;
ROM[6418] <= 32'b00000000111000111000001110110011;
ROM[6419] <= 32'b00000000011100010010000000100011;
ROM[6420] <= 32'b00000000010000010000000100010011;
ROM[6421] <= 32'b00000000001100010010000000100011;
ROM[6422] <= 32'b00000000010000010000000100010011;
ROM[6423] <= 32'b00000000010000010010000000100011;
ROM[6424] <= 32'b00000000010000010000000100010011;
ROM[6425] <= 32'b00000000010100010010000000100011;
ROM[6426] <= 32'b00000000010000010000000100010011;
ROM[6427] <= 32'b00000000011000010010000000100011;
ROM[6428] <= 32'b00000000010000010000000100010011;
ROM[6429] <= 32'b00000001010000000000001110010011;
ROM[6430] <= 32'b00000000100000111000001110010011;
ROM[6431] <= 32'b01000000011100010000001110110011;
ROM[6432] <= 32'b00000000011100000000001000110011;
ROM[6433] <= 32'b00000000001000000000000110110011;
ROM[6434] <= 32'b00111010010000001011000011101111;
ROM[6435] <= 32'b11111111110000010000000100010011;
ROM[6436] <= 32'b00000000000000010010001110000011;
ROM[6437] <= 32'b11111111110000010000000100010011;
ROM[6438] <= 32'b00000000000000010010010000000011;
ROM[6439] <= 32'b00000000011101000000001110110011;
ROM[6440] <= 32'b00000000011100010010000000100011;
ROM[6441] <= 32'b00000000010000010000000100010011;
ROM[6442] <= 32'b11111111110000010000000100010011;
ROM[6443] <= 32'b00000000000000010010001110000011;
ROM[6444] <= 32'b00000000000000111000001100010011;
ROM[6445] <= 32'b11111111110000010000000100010011;
ROM[6446] <= 32'b00000000000000010010001110000011;
ROM[6447] <= 32'b00000000110100110000010000110011;
ROM[6448] <= 32'b00000000011101000010000000100011;
ROM[6449] <= 32'b00000000011100000000001110010011;
ROM[6450] <= 32'b00000000011100010010000000100011;
ROM[6451] <= 32'b00000000010000010000000100010011;
ROM[6452] <= 32'b00000011110000011010001110000011;
ROM[6453] <= 32'b00000000011100010010000000100011;
ROM[6454] <= 32'b00000000010000010000000100010011;
ROM[6455] <= 32'b00000000010000000000001110010011;
ROM[6456] <= 32'b00000000011100010010000000100011;
ROM[6457] <= 32'b00000000010000010000000100010011;
ROM[6458] <= 32'b00000000010000000000001110010011;
ROM[6459] <= 32'b00000000011100010010000000100011;
ROM[6460] <= 32'b00000000010000010000000100010011;
ROM[6461] <= 32'b00000000000000000110001110110111;
ROM[6462] <= 32'b01010100000000111000001110010011;
ROM[6463] <= 32'b00000000111000111000001110110011;
ROM[6464] <= 32'b00000000011100010010000000100011;
ROM[6465] <= 32'b00000000010000010000000100010011;
ROM[6466] <= 32'b00000000001100010010000000100011;
ROM[6467] <= 32'b00000000010000010000000100010011;
ROM[6468] <= 32'b00000000010000010010000000100011;
ROM[6469] <= 32'b00000000010000010000000100010011;
ROM[6470] <= 32'b00000000010100010010000000100011;
ROM[6471] <= 32'b00000000010000010000000100010011;
ROM[6472] <= 32'b00000000011000010010000000100011;
ROM[6473] <= 32'b00000000010000010000000100010011;
ROM[6474] <= 32'b00000001010000000000001110010011;
ROM[6475] <= 32'b00000000100000111000001110010011;
ROM[6476] <= 32'b01000000011100010000001110110011;
ROM[6477] <= 32'b00000000011100000000001000110011;
ROM[6478] <= 32'b00000000001000000000000110110011;
ROM[6479] <= 32'b00101111000000001011000011101111;
ROM[6480] <= 32'b11111111110000010000000100010011;
ROM[6481] <= 32'b00000000000000010010001110000011;
ROM[6482] <= 32'b11111111110000010000000100010011;
ROM[6483] <= 32'b00000000000000010010010000000011;
ROM[6484] <= 32'b00000000011101000000001110110011;
ROM[6485] <= 32'b00000000011100010010000000100011;
ROM[6486] <= 32'b00000000010000010000000100010011;
ROM[6487] <= 32'b11111111110000010000000100010011;
ROM[6488] <= 32'b00000000000000010010001110000011;
ROM[6489] <= 32'b00000000000000111000001100010011;
ROM[6490] <= 32'b11111111110000010000000100010011;
ROM[6491] <= 32'b00000000000000010010001110000011;
ROM[6492] <= 32'b00000000110100110000010000110011;
ROM[6493] <= 32'b00000000011101000010000000100011;
ROM[6494] <= 32'b00000000000000000000001110010011;
ROM[6495] <= 32'b00000000011100010010000000100011;
ROM[6496] <= 32'b00000000010000010000000100010011;
ROM[6497] <= 32'b11111111110000010000000100010011;
ROM[6498] <= 32'b00000000000000010010001110000011;
ROM[6499] <= 32'b00000000011100011010010000100011;
ROM[6500] <= 32'b00000101111100000000001110010011;
ROM[6501] <= 32'b00000000011100010010000000100011;
ROM[6502] <= 32'b00000000010000010000000100010011;
ROM[6503] <= 32'b11111111110000010000000100010011;
ROM[6504] <= 32'b00000000000000010010001110000011;
ROM[6505] <= 32'b00000010011100011010011000100011;
ROM[6506] <= 32'b00000000100000011010001110000011;
ROM[6507] <= 32'b00000000011100010010000000100011;
ROM[6508] <= 32'b00000000010000010000000100010011;
ROM[6509] <= 32'b00000000010100000000001110010011;
ROM[6510] <= 32'b00000000011100010010000000100011;
ROM[6511] <= 32'b00000000010000010000000100010011;
ROM[6512] <= 32'b11111111110000010000000100010011;
ROM[6513] <= 32'b00000000000000010010001110000011;
ROM[6514] <= 32'b11111111110000010000000100010011;
ROM[6515] <= 32'b00000000000000010010010000000011;
ROM[6516] <= 32'b00000000011101000010001110110011;
ROM[6517] <= 32'b00000000011100010010000000100011;
ROM[6518] <= 32'b00000000010000010000000100010011;
ROM[6519] <= 32'b11111111110000010000000100010011;
ROM[6520] <= 32'b00000000000000010010001110000011;
ROM[6521] <= 32'b01000000011100000000001110110011;
ROM[6522] <= 32'b00000000000100111000001110010011;
ROM[6523] <= 32'b00000000011100010010000000100011;
ROM[6524] <= 32'b00000000010000010000000100010011;
ROM[6525] <= 32'b11111111110000010000000100010011;
ROM[6526] <= 32'b00000000000000010010001110000011;
ROM[6527] <= 32'b00000000000000111000101001100011;
ROM[6528] <= 32'b00000000000000001101001110110111;
ROM[6529] <= 32'b01110010010000111000001110010011;
ROM[6530] <= 32'b00000000111000111000001110110011;
ROM[6531] <= 32'b00000000000000111000000011100111;
ROM[6532] <= 32'b00000000011000000000001110010011;
ROM[6533] <= 32'b00000000011100010010000000100011;
ROM[6534] <= 32'b00000000010000010000000100010011;
ROM[6535] <= 32'b11111111110000010000000100010011;
ROM[6536] <= 32'b00000000000000010010001110000011;
ROM[6537] <= 32'b00000000011100011010101000100011;
ROM[6538] <= 32'b00000001101000000000001110010011;
ROM[6539] <= 32'b00000000011100010010000000100011;
ROM[6540] <= 32'b00000000010000010000000100010011;
ROM[6541] <= 32'b00000000000000000110001110110111;
ROM[6542] <= 32'b01101000000000111000001110010011;
ROM[6543] <= 32'b00000000111000111000001110110011;
ROM[6544] <= 32'b00000000011100010010000000100011;
ROM[6545] <= 32'b00000000010000010000000100010011;
ROM[6546] <= 32'b00000000001100010010000000100011;
ROM[6547] <= 32'b00000000010000010000000100010011;
ROM[6548] <= 32'b00000000010000010010000000100011;
ROM[6549] <= 32'b00000000010000010000000100010011;
ROM[6550] <= 32'b00000000010100010010000000100011;
ROM[6551] <= 32'b00000000010000010000000100010011;
ROM[6552] <= 32'b00000000011000010010000000100011;
ROM[6553] <= 32'b00000000010000010000000100010011;
ROM[6554] <= 32'b00000001010000000000001110010011;
ROM[6555] <= 32'b00000000010000111000001110010011;
ROM[6556] <= 32'b01000000011100010000001110110011;
ROM[6557] <= 32'b00000000011100000000001000110011;
ROM[6558] <= 32'b00000000001000000000000110110011;
ROM[6559] <= 32'b10100000010111111001000011101111;
ROM[6560] <= 32'b11111111110000010000000100010011;
ROM[6561] <= 32'b00000000000000010010001110000011;
ROM[6562] <= 32'b00000000011100011010001000100011;
ROM[6563] <= 32'b00000000000000000000001110010011;
ROM[6564] <= 32'b00000000011100010010000000100011;
ROM[6565] <= 32'b00000000010000010000000100010011;
ROM[6566] <= 32'b11111111110000010000000100010011;
ROM[6567] <= 32'b00000000000000010010001110000011;
ROM[6568] <= 32'b00000000011100011010011000100011;
ROM[6569] <= 32'b00000000110000011010001110000011;
ROM[6570] <= 32'b00000000011100010010000000100011;
ROM[6571] <= 32'b00000000010000010000000100010011;
ROM[6572] <= 32'b00000001101000000000001110010011;
ROM[6573] <= 32'b00000000011100010010000000100011;
ROM[6574] <= 32'b00000000010000010000000100010011;
ROM[6575] <= 32'b11111111110000010000000100010011;
ROM[6576] <= 32'b00000000000000010010001110000011;
ROM[6577] <= 32'b11111111110000010000000100010011;
ROM[6578] <= 32'b00000000000000010010010000000011;
ROM[6579] <= 32'b00000000011101000010001110110011;
ROM[6580] <= 32'b00000000011100010010000000100011;
ROM[6581] <= 32'b00000000010000010000000100010011;
ROM[6582] <= 32'b11111111110000010000000100010011;
ROM[6583] <= 32'b00000000000000010010001110000011;
ROM[6584] <= 32'b01000000011100000000001110110011;
ROM[6585] <= 32'b00000000000100111000001110010011;
ROM[6586] <= 32'b00000000011100010010000000100011;
ROM[6587] <= 32'b00000000010000010000000100010011;
ROM[6588] <= 32'b11111111110000010000000100010011;
ROM[6589] <= 32'b00000000000000010010001110000011;
ROM[6590] <= 32'b00000000000000111000101001100011;
ROM[6591] <= 32'b00000000000000000111001110110111;
ROM[6592] <= 32'b10000000010000111000001110010011;
ROM[6593] <= 32'b00000000111000111000001110110011;
ROM[6594] <= 32'b00000000000000111000000011100111;
ROM[6595] <= 32'b00000000000000000000001110010011;
ROM[6596] <= 32'b00000000011100010010000000100011;
ROM[6597] <= 32'b00000000010000010000000100010011;
ROM[6598] <= 32'b00000000010000011010001110000011;
ROM[6599] <= 32'b00000000011100010010000000100011;
ROM[6600] <= 32'b00000000010000010000000100010011;
ROM[6601] <= 32'b00000000110000011010001110000011;
ROM[6602] <= 32'b00000000011100010010000000100011;
ROM[6603] <= 32'b00000000010000010000000100010011;
ROM[6604] <= 32'b00000000010000000000001110010011;
ROM[6605] <= 32'b00000000011100010010000000100011;
ROM[6606] <= 32'b00000000010000010000000100010011;
ROM[6607] <= 32'b00000000000000000110001110110111;
ROM[6608] <= 32'b01111000100000111000001110010011;
ROM[6609] <= 32'b00000000111000111000001110110011;
ROM[6610] <= 32'b00000000011100010010000000100011;
ROM[6611] <= 32'b00000000010000010000000100010011;
ROM[6612] <= 32'b00000000001100010010000000100011;
ROM[6613] <= 32'b00000000010000010000000100010011;
ROM[6614] <= 32'b00000000010000010010000000100011;
ROM[6615] <= 32'b00000000010000010000000100010011;
ROM[6616] <= 32'b00000000010100010010000000100011;
ROM[6617] <= 32'b00000000010000010000000100010011;
ROM[6618] <= 32'b00000000011000010010000000100011;
ROM[6619] <= 32'b00000000010000010000000100010011;
ROM[6620] <= 32'b00000001010000000000001110010011;
ROM[6621] <= 32'b00000000100000111000001110010011;
ROM[6622] <= 32'b01000000011100010000001110110011;
ROM[6623] <= 32'b00000000011100000000001000110011;
ROM[6624] <= 32'b00000000001000000000000110110011;
ROM[6625] <= 32'b00001010100000001011000011101111;
ROM[6626] <= 32'b11111111110000010000000100010011;
ROM[6627] <= 32'b00000000000000010010001110000011;
ROM[6628] <= 32'b11111111110000010000000100010011;
ROM[6629] <= 32'b00000000000000010010010000000011;
ROM[6630] <= 32'b00000000011101000000001110110011;
ROM[6631] <= 32'b00000000011100010010000000100011;
ROM[6632] <= 32'b00000000010000010000000100010011;
ROM[6633] <= 32'b11111111110000010000000100010011;
ROM[6634] <= 32'b00000000000000010010001110000011;
ROM[6635] <= 32'b00000000000000111000001100010011;
ROM[6636] <= 32'b11111111110000010000000100010011;
ROM[6637] <= 32'b00000000000000010010001110000011;
ROM[6638] <= 32'b00000000110100110000010000110011;
ROM[6639] <= 32'b00000000011101000010000000100011;
ROM[6640] <= 32'b00000000110000011010001110000011;
ROM[6641] <= 32'b00000000011100010010000000100011;
ROM[6642] <= 32'b00000000010000010000000100010011;
ROM[6643] <= 32'b00000000000100000000001110010011;
ROM[6644] <= 32'b00000000011100010010000000100011;
ROM[6645] <= 32'b00000000010000010000000100010011;
ROM[6646] <= 32'b11111111110000010000000100010011;
ROM[6647] <= 32'b00000000000000010010001110000011;
ROM[6648] <= 32'b11111111110000010000000100010011;
ROM[6649] <= 32'b00000000000000010010010000000011;
ROM[6650] <= 32'b00000000011101000000001110110011;
ROM[6651] <= 32'b00000000011100010010000000100011;
ROM[6652] <= 32'b00000000010000010000000100010011;
ROM[6653] <= 32'b11111111110000010000000100010011;
ROM[6654] <= 32'b00000000000000010010001110000011;
ROM[6655] <= 32'b00000000011100011010011000100011;
ROM[6656] <= 32'b11101010010111111111000011101111;
ROM[6657] <= 32'b00000011110000011010001110000011;
ROM[6658] <= 32'b00000000011100010010000000100011;
ROM[6659] <= 32'b00000000010000010000000100010011;
ROM[6660] <= 32'b00000000100000011010001110000011;
ROM[6661] <= 32'b00000000011100010010000000100011;
ROM[6662] <= 32'b00000000010000010000000100010011;
ROM[6663] <= 32'b00000000010000000000001110010011;
ROM[6664] <= 32'b00000000011100010010000000100011;
ROM[6665] <= 32'b00000000010000010000000100010011;
ROM[6666] <= 32'b00000000000000000111001110110111;
ROM[6667] <= 32'b10000111010000111000001110010011;
ROM[6668] <= 32'b00000000111000111000001110110011;
ROM[6669] <= 32'b00000000011100010010000000100011;
ROM[6670] <= 32'b00000000010000010000000100010011;
ROM[6671] <= 32'b00000000001100010010000000100011;
ROM[6672] <= 32'b00000000010000010000000100010011;
ROM[6673] <= 32'b00000000010000010010000000100011;
ROM[6674] <= 32'b00000000010000010000000100010011;
ROM[6675] <= 32'b00000000010100010010000000100011;
ROM[6676] <= 32'b00000000010000010000000100010011;
ROM[6677] <= 32'b00000000011000010010000000100011;
ROM[6678] <= 32'b00000000010000010000000100010011;
ROM[6679] <= 32'b00000001010000000000001110010011;
ROM[6680] <= 32'b00000000100000111000001110010011;
ROM[6681] <= 32'b01000000011100010000001110110011;
ROM[6682] <= 32'b00000000011100000000001000110011;
ROM[6683] <= 32'b00000000001000000000000110110011;
ROM[6684] <= 32'b01111011110100001010000011101111;
ROM[6685] <= 32'b11111111110000010000000100010011;
ROM[6686] <= 32'b00000000000000010010001110000011;
ROM[6687] <= 32'b11111111110000010000000100010011;
ROM[6688] <= 32'b00000000000000010010010000000011;
ROM[6689] <= 32'b00000000011101000000001110110011;
ROM[6690] <= 32'b00000000011100010010000000100011;
ROM[6691] <= 32'b00000000010000010000000100010011;
ROM[6692] <= 32'b11111111110000010000000100010011;
ROM[6693] <= 32'b00000000000000010010001110000011;
ROM[6694] <= 32'b00000000000000111000001100010011;
ROM[6695] <= 32'b00000000110100110000010000110011;
ROM[6696] <= 32'b00000000000001000010001110000011;
ROM[6697] <= 32'b00000000011100010010000000100011;
ROM[6698] <= 32'b00000000010000010000000100010011;
ROM[6699] <= 32'b11111111110000010000000100010011;
ROM[6700] <= 32'b00000000000000010010001110000011;
ROM[6701] <= 32'b00000000011100011010100000100011;
ROM[6702] <= 32'b00000000100000011010001110000011;
ROM[6703] <= 32'b00000000011100010010000000100011;
ROM[6704] <= 32'b00000000010000010000000100010011;
ROM[6705] <= 32'b00000000000000000000001110010011;
ROM[6706] <= 32'b00000000011100010010000000100011;
ROM[6707] <= 32'b00000000010000010000000100010011;
ROM[6708] <= 32'b11111111110000010000000100010011;
ROM[6709] <= 32'b00000000000000010010001110000011;
ROM[6710] <= 32'b11111111110000010000000100010011;
ROM[6711] <= 32'b00000000000000010010010000000011;
ROM[6712] <= 32'b00000000011101000010010010110011;
ROM[6713] <= 32'b00000000100000111010010100110011;
ROM[6714] <= 32'b00000000101001001000001110110011;
ROM[6715] <= 32'b00000000000100111000001110010011;
ROM[6716] <= 32'b00000000000100111111001110010011;
ROM[6717] <= 32'b00000000011100010010000000100011;
ROM[6718] <= 32'b00000000010000010000000100010011;
ROM[6719] <= 32'b11111111110000010000000100010011;
ROM[6720] <= 32'b00000000000000010010001110000011;
ROM[6721] <= 32'b00000000000000111000101001100011;
ROM[6722] <= 32'b00000000000000000111001110110111;
ROM[6723] <= 32'b01111000100000111000001110010011;
ROM[6724] <= 32'b00000000111000111000001110110011;
ROM[6725] <= 32'b00000000000000111000000011100111;
ROM[6726] <= 32'b00000000100000011010001110000011;
ROM[6727] <= 32'b00000000011100010010000000100011;
ROM[6728] <= 32'b00000000010000010000000100010011;
ROM[6729] <= 32'b00000000000100000000001110010011;
ROM[6730] <= 32'b00000000011100010010000000100011;
ROM[6731] <= 32'b00000000010000010000000100010011;
ROM[6732] <= 32'b11111111110000010000000100010011;
ROM[6733] <= 32'b00000000000000010010001110000011;
ROM[6734] <= 32'b11111111110000010000000100010011;
ROM[6735] <= 32'b00000000000000010010010000000011;
ROM[6736] <= 32'b00000000011101000010010010110011;
ROM[6737] <= 32'b00000000100000111010010100110011;
ROM[6738] <= 32'b00000000101001001000001110110011;
ROM[6739] <= 32'b00000000000100111000001110010011;
ROM[6740] <= 32'b00000000000100111111001110010011;
ROM[6741] <= 32'b00000000011100010010000000100011;
ROM[6742] <= 32'b00000000010000010000000100010011;
ROM[6743] <= 32'b11111111110000010000000100010011;
ROM[6744] <= 32'b00000000000000010010001110000011;
ROM[6745] <= 32'b00000000000000111000101001100011;
ROM[6746] <= 32'b00000000000000000111001110110111;
ROM[6747] <= 32'b00110101100000111000001110010011;
ROM[6748] <= 32'b00000000111000111000001110110011;
ROM[6749] <= 32'b00000000000000111000000011100111;
ROM[6750] <= 32'b00000000100000011010001110000011;
ROM[6751] <= 32'b00000000011100010010000000100011;
ROM[6752] <= 32'b00000000010000010000000100010011;
ROM[6753] <= 32'b00000000001000000000001110010011;
ROM[6754] <= 32'b00000000011100010010000000100011;
ROM[6755] <= 32'b00000000010000010000000100010011;
ROM[6756] <= 32'b11111111110000010000000100010011;
ROM[6757] <= 32'b00000000000000010010001110000011;
ROM[6758] <= 32'b11111111110000010000000100010011;
ROM[6759] <= 32'b00000000000000010010010000000011;
ROM[6760] <= 32'b00000000011101000010010010110011;
ROM[6761] <= 32'b00000000100000111010010100110011;
ROM[6762] <= 32'b00000000101001001000001110110011;
ROM[6763] <= 32'b00000000000100111000001110010011;
ROM[6764] <= 32'b00000000000100111111001110010011;
ROM[6765] <= 32'b00000000011100010010000000100011;
ROM[6766] <= 32'b00000000010000010000000100010011;
ROM[6767] <= 32'b11111111110000010000000100010011;
ROM[6768] <= 32'b00000000000000010010001110000011;
ROM[6769] <= 32'b00000000000000111000101001100011;
ROM[6770] <= 32'b00000000000000000111001110110111;
ROM[6771] <= 32'b00000011000000111000001110010011;
ROM[6772] <= 32'b00000000111000111000001110110011;
ROM[6773] <= 32'b00000000000000111000000011100111;
ROM[6774] <= 32'b00000000100000011010001110000011;
ROM[6775] <= 32'b00000000011100010010000000100011;
ROM[6776] <= 32'b00000000010000010000000100010011;
ROM[6777] <= 32'b00000000001100000000001110010011;
ROM[6778] <= 32'b00000000011100010010000000100011;
ROM[6779] <= 32'b00000000010000010000000100010011;
ROM[6780] <= 32'b11111111110000010000000100010011;
ROM[6781] <= 32'b00000000000000010010001110000011;
ROM[6782] <= 32'b11111111110000010000000100010011;
ROM[6783] <= 32'b00000000000000010010010000000011;
ROM[6784] <= 32'b00000000011101000010010010110011;
ROM[6785] <= 32'b00000000100000111010010100110011;
ROM[6786] <= 32'b00000000101001001000001110110011;
ROM[6787] <= 32'b00000000000100111000001110010011;
ROM[6788] <= 32'b00000000000100111111001110010011;
ROM[6789] <= 32'b00000000011100010010000000100011;
ROM[6790] <= 32'b00000000010000010000000100010011;
ROM[6791] <= 32'b11111111110000010000000100010011;
ROM[6792] <= 32'b00000000000000010010001110000011;
ROM[6793] <= 32'b00000000000000111000101001100011;
ROM[6794] <= 32'b00000000000000000111001110110111;
ROM[6795] <= 32'b11010000100000111000001110010011;
ROM[6796] <= 32'b00000000111000111000001110110011;
ROM[6797] <= 32'b00000000000000111000000011100111;
ROM[6798] <= 32'b00000000011100000000001110010011;
ROM[6799] <= 32'b00000000011100010010000000100011;
ROM[6800] <= 32'b00000000010000010000000100010011;
ROM[6801] <= 32'b00000000000000000111001110110111;
ROM[6802] <= 32'b10101001000000111000001110010011;
ROM[6803] <= 32'b00000000111000111000001110110011;
ROM[6804] <= 32'b00000000011100010010000000100011;
ROM[6805] <= 32'b00000000010000010000000100010011;
ROM[6806] <= 32'b00000000001100010010000000100011;
ROM[6807] <= 32'b00000000010000010000000100010011;
ROM[6808] <= 32'b00000000010000010010000000100011;
ROM[6809] <= 32'b00000000010000010000000100010011;
ROM[6810] <= 32'b00000000010100010010000000100011;
ROM[6811] <= 32'b00000000010000010000000100010011;
ROM[6812] <= 32'b00000000011000010010000000100011;
ROM[6813] <= 32'b00000000010000010000000100010011;
ROM[6814] <= 32'b00000001010000000000001110010011;
ROM[6815] <= 32'b00000000010000111000001110010011;
ROM[6816] <= 32'b01000000011100010000001110110011;
ROM[6817] <= 32'b00000000011100000000001000110011;
ROM[6818] <= 32'b00000000001000000000000110110011;
ROM[6819] <= 32'b01001011000100100010000011101111;
ROM[6820] <= 32'b00000101111100000000001110010011;
ROM[6821] <= 32'b00000000011100010010000000100011;
ROM[6822] <= 32'b00000000010000010000000100010011;
ROM[6823] <= 32'b00000000000000000111001110110111;
ROM[6824] <= 32'b10101110100000111000001110010011;
ROM[6825] <= 32'b00000000111000111000001110110011;
ROM[6826] <= 32'b00000000011100010010000000100011;
ROM[6827] <= 32'b00000000010000010000000100010011;
ROM[6828] <= 32'b00000000001100010010000000100011;
ROM[6829] <= 32'b00000000010000010000000100010011;
ROM[6830] <= 32'b00000000010000010010000000100011;
ROM[6831] <= 32'b00000000010000010000000100010011;
ROM[6832] <= 32'b00000000010100010010000000100011;
ROM[6833] <= 32'b00000000010000010000000100010011;
ROM[6834] <= 32'b00000000011000010010000000100011;
ROM[6835] <= 32'b00000000010000010000000100010011;
ROM[6836] <= 32'b00000001010000000000001110010011;
ROM[6837] <= 32'b00000000100000111000001110010011;
ROM[6838] <= 32'b01000000011100010000001110110011;
ROM[6839] <= 32'b00000000011100000000001000110011;
ROM[6840] <= 32'b00000000001000000000000110110011;
ROM[6841] <= 32'b00001100100000100011000011101111;
ROM[6842] <= 32'b00000101111100000000001110010011;
ROM[6843] <= 32'b00000000011100010010000000100011;
ROM[6844] <= 32'b00000000010000010000000100010011;
ROM[6845] <= 32'b00000000000000000111001110110111;
ROM[6846] <= 32'b10110100000000111000001110010011;
ROM[6847] <= 32'b00000000111000111000001110110011;
ROM[6848] <= 32'b00000000011100010010000000100011;
ROM[6849] <= 32'b00000000010000010000000100010011;
ROM[6850] <= 32'b00000000001100010010000000100011;
ROM[6851] <= 32'b00000000010000010000000100010011;
ROM[6852] <= 32'b00000000010000010010000000100011;
ROM[6853] <= 32'b00000000010000010000000100010011;
ROM[6854] <= 32'b00000000010100010010000000100011;
ROM[6855] <= 32'b00000000010000010000000100010011;
ROM[6856] <= 32'b00000000011000010010000000100011;
ROM[6857] <= 32'b00000000010000010000000100010011;
ROM[6858] <= 32'b00000001010000000000001110010011;
ROM[6859] <= 32'b00000000100000111000001110010011;
ROM[6860] <= 32'b01000000011100010000001110110011;
ROM[6861] <= 32'b00000000011100000000001000110011;
ROM[6862] <= 32'b00000000001000000000000110110011;
ROM[6863] <= 32'b00000111000000100011000011101111;
ROM[6864] <= 32'b00000101111100000000001110010011;
ROM[6865] <= 32'b00000000011100010010000000100011;
ROM[6866] <= 32'b00000000010000010000000100010011;
ROM[6867] <= 32'b00000000000000000111001110110111;
ROM[6868] <= 32'b10111001100000111000001110010011;
ROM[6869] <= 32'b00000000111000111000001110110011;
ROM[6870] <= 32'b00000000011100010010000000100011;
ROM[6871] <= 32'b00000000010000010000000100010011;
ROM[6872] <= 32'b00000000001100010010000000100011;
ROM[6873] <= 32'b00000000010000010000000100010011;
ROM[6874] <= 32'b00000000010000010010000000100011;
ROM[6875] <= 32'b00000000010000010000000100010011;
ROM[6876] <= 32'b00000000010100010010000000100011;
ROM[6877] <= 32'b00000000010000010000000100010011;
ROM[6878] <= 32'b00000000011000010010000000100011;
ROM[6879] <= 32'b00000000010000010000000100010011;
ROM[6880] <= 32'b00000001010000000000001110010011;
ROM[6881] <= 32'b00000000100000111000001110010011;
ROM[6882] <= 32'b01000000011100010000001110110011;
ROM[6883] <= 32'b00000000011100000000001000110011;
ROM[6884] <= 32'b00000000001000000000000110110011;
ROM[6885] <= 32'b00000001100000100011000011101111;
ROM[6886] <= 32'b00000101111100000000001110010011;
ROM[6887] <= 32'b00000000011100010010000000100011;
ROM[6888] <= 32'b00000000010000010000000100010011;
ROM[6889] <= 32'b00000000000000000111001110110111;
ROM[6890] <= 32'b10111111000000111000001110010011;
ROM[6891] <= 32'b00000000111000111000001110110011;
ROM[6892] <= 32'b00000000011100010010000000100011;
ROM[6893] <= 32'b00000000010000010000000100010011;
ROM[6894] <= 32'b00000000001100010010000000100011;
ROM[6895] <= 32'b00000000010000010000000100010011;
ROM[6896] <= 32'b00000000010000010010000000100011;
ROM[6897] <= 32'b00000000010000010000000100010011;
ROM[6898] <= 32'b00000000010100010010000000100011;
ROM[6899] <= 32'b00000000010000010000000100010011;
ROM[6900] <= 32'b00000000011000010010000000100011;
ROM[6901] <= 32'b00000000010000010000000100010011;
ROM[6902] <= 32'b00000001010000000000001110010011;
ROM[6903] <= 32'b00000000100000111000001110010011;
ROM[6904] <= 32'b01000000011100010000001110110011;
ROM[6905] <= 32'b00000000011100000000001000110011;
ROM[6906] <= 32'b00000000001000000000000110110011;
ROM[6907] <= 32'b01111100000100100010000011101111;
ROM[6908] <= 32'b00000101111100000000001110010011;
ROM[6909] <= 32'b00000000011100010010000000100011;
ROM[6910] <= 32'b00000000010000010000000100010011;
ROM[6911] <= 32'b00000000000000000111001110110111;
ROM[6912] <= 32'b11000100100000111000001110010011;
ROM[6913] <= 32'b00000000111000111000001110110011;
ROM[6914] <= 32'b00000000011100010010000000100011;
ROM[6915] <= 32'b00000000010000010000000100010011;
ROM[6916] <= 32'b00000000001100010010000000100011;
ROM[6917] <= 32'b00000000010000010000000100010011;
ROM[6918] <= 32'b00000000010000010010000000100011;
ROM[6919] <= 32'b00000000010000010000000100010011;
ROM[6920] <= 32'b00000000010100010010000000100011;
ROM[6921] <= 32'b00000000010000010000000100010011;
ROM[6922] <= 32'b00000000011000010010000000100011;
ROM[6923] <= 32'b00000000010000010000000100010011;
ROM[6924] <= 32'b00000001010000000000001110010011;
ROM[6925] <= 32'b00000000100000111000001110010011;
ROM[6926] <= 32'b01000000011100010000001110110011;
ROM[6927] <= 32'b00000000011100000000001000110011;
ROM[6928] <= 32'b00000000001000000000000110110011;
ROM[6929] <= 32'b01110110100100100010000011101111;
ROM[6930] <= 32'b00000101111100000000001110010011;
ROM[6931] <= 32'b00000000011100010010000000100011;
ROM[6932] <= 32'b00000000010000010000000100010011;
ROM[6933] <= 32'b00000000000000000111001110110111;
ROM[6934] <= 32'b11001010000000111000001110010011;
ROM[6935] <= 32'b00000000111000111000001110110011;
ROM[6936] <= 32'b00000000011100010010000000100011;
ROM[6937] <= 32'b00000000010000010000000100010011;
ROM[6938] <= 32'b00000000001100010010000000100011;
ROM[6939] <= 32'b00000000010000010000000100010011;
ROM[6940] <= 32'b00000000010000010010000000100011;
ROM[6941] <= 32'b00000000010000010000000100010011;
ROM[6942] <= 32'b00000000010100010010000000100011;
ROM[6943] <= 32'b00000000010000010000000100010011;
ROM[6944] <= 32'b00000000011000010010000000100011;
ROM[6945] <= 32'b00000000010000010000000100010011;
ROM[6946] <= 32'b00000001010000000000001110010011;
ROM[6947] <= 32'b00000000100000111000001110010011;
ROM[6948] <= 32'b01000000011100010000001110110011;
ROM[6949] <= 32'b00000000011100000000001000110011;
ROM[6950] <= 32'b00000000001000000000000110110011;
ROM[6951] <= 32'b01110001000100100010000011101111;
ROM[6952] <= 32'b00000101111100000000001110010011;
ROM[6953] <= 32'b00000000011100010010000000100011;
ROM[6954] <= 32'b00000000010000010000000100010011;
ROM[6955] <= 32'b00000000000000000111001110110111;
ROM[6956] <= 32'b11001111100000111000001110010011;
ROM[6957] <= 32'b00000000111000111000001110110011;
ROM[6958] <= 32'b00000000011100010010000000100011;
ROM[6959] <= 32'b00000000010000010000000100010011;
ROM[6960] <= 32'b00000000001100010010000000100011;
ROM[6961] <= 32'b00000000010000010000000100010011;
ROM[6962] <= 32'b00000000010000010010000000100011;
ROM[6963] <= 32'b00000000010000010000000100010011;
ROM[6964] <= 32'b00000000010100010010000000100011;
ROM[6965] <= 32'b00000000010000010000000100010011;
ROM[6966] <= 32'b00000000011000010010000000100011;
ROM[6967] <= 32'b00000000010000010000000100010011;
ROM[6968] <= 32'b00000001010000000000001110010011;
ROM[6969] <= 32'b00000000100000111000001110010011;
ROM[6970] <= 32'b01000000011100010000001110110011;
ROM[6971] <= 32'b00000000011100000000001000110011;
ROM[6972] <= 32'b00000000001000000000000110110011;
ROM[6973] <= 32'b01101011100100100010000011101111;
ROM[6974] <= 32'b11111111110000010000000100010011;
ROM[6975] <= 32'b00000000000000010010001110000011;
ROM[6976] <= 32'b00000000011100011010110000100011;
ROM[6977] <= 32'b00110010100000000000000011101111;
ROM[6978] <= 32'b00000000100000000000001110010011;
ROM[6979] <= 32'b00000000011100010010000000100011;
ROM[6980] <= 32'b00000000010000010000000100010011;
ROM[6981] <= 32'b00000000000000000111001110110111;
ROM[6982] <= 32'b11010110000000111000001110010011;
ROM[6983] <= 32'b00000000111000111000001110110011;
ROM[6984] <= 32'b00000000011100010010000000100011;
ROM[6985] <= 32'b00000000010000010000000100010011;
ROM[6986] <= 32'b00000000001100010010000000100011;
ROM[6987] <= 32'b00000000010000010000000100010011;
ROM[6988] <= 32'b00000000010000010010000000100011;
ROM[6989] <= 32'b00000000010000010000000100010011;
ROM[6990] <= 32'b00000000010100010010000000100011;
ROM[6991] <= 32'b00000000010000010000000100010011;
ROM[6992] <= 32'b00000000011000010010000000100011;
ROM[6993] <= 32'b00000000010000010000000100010011;
ROM[6994] <= 32'b00000001010000000000001110010011;
ROM[6995] <= 32'b00000000010000111000001110010011;
ROM[6996] <= 32'b01000000011100010000001110110011;
ROM[6997] <= 32'b00000000011100000000001000110011;
ROM[6998] <= 32'b00000000001000000000000110110011;
ROM[6999] <= 32'b00011110000100100010000011101111;
ROM[7000] <= 32'b00000101111100000000001110010011;
ROM[7001] <= 32'b00000000011100010010000000100011;
ROM[7002] <= 32'b00000000010000010000000100010011;
ROM[7003] <= 32'b00000000000000000111001110110111;
ROM[7004] <= 32'b11011011100000111000001110010011;
ROM[7005] <= 32'b00000000111000111000001110110011;
ROM[7006] <= 32'b00000000011100010010000000100011;
ROM[7007] <= 32'b00000000010000010000000100010011;
ROM[7008] <= 32'b00000000001100010010000000100011;
ROM[7009] <= 32'b00000000010000010000000100010011;
ROM[7010] <= 32'b00000000010000010010000000100011;
ROM[7011] <= 32'b00000000010000010000000100010011;
ROM[7012] <= 32'b00000000010100010010000000100011;
ROM[7013] <= 32'b00000000010000010000000100010011;
ROM[7014] <= 32'b00000000011000010010000000100011;
ROM[7015] <= 32'b00000000010000010000000100010011;
ROM[7016] <= 32'b00000001010000000000001110010011;
ROM[7017] <= 32'b00000000100000111000001110010011;
ROM[7018] <= 32'b01000000011100010000001110110011;
ROM[7019] <= 32'b00000000011100000000001000110011;
ROM[7020] <= 32'b00000000001000000000000110110011;
ROM[7021] <= 32'b01011111100100100010000011101111;
ROM[7022] <= 32'b00000101111100000000001110010011;
ROM[7023] <= 32'b00000000011100010010000000100011;
ROM[7024] <= 32'b00000000010000010000000100010011;
ROM[7025] <= 32'b00000000000000000111001110110111;
ROM[7026] <= 32'b11100001000000111000001110010011;
ROM[7027] <= 32'b00000000111000111000001110110011;
ROM[7028] <= 32'b00000000011100010010000000100011;
ROM[7029] <= 32'b00000000010000010000000100010011;
ROM[7030] <= 32'b00000000001100010010000000100011;
ROM[7031] <= 32'b00000000010000010000000100010011;
ROM[7032] <= 32'b00000000010000010010000000100011;
ROM[7033] <= 32'b00000000010000010000000100010011;
ROM[7034] <= 32'b00000000010100010010000000100011;
ROM[7035] <= 32'b00000000010000010000000100010011;
ROM[7036] <= 32'b00000000011000010010000000100011;
ROM[7037] <= 32'b00000000010000010000000100010011;
ROM[7038] <= 32'b00000001010000000000001110010011;
ROM[7039] <= 32'b00000000100000111000001110010011;
ROM[7040] <= 32'b01000000011100010000001110110011;
ROM[7041] <= 32'b00000000011100000000001000110011;
ROM[7042] <= 32'b00000000001000000000000110110011;
ROM[7043] <= 32'b01011010000100100010000011101111;
ROM[7044] <= 32'b00000101111100000000001110010011;
ROM[7045] <= 32'b00000000011100010010000000100011;
ROM[7046] <= 32'b00000000010000010000000100010011;
ROM[7047] <= 32'b00000000000000000111001110110111;
ROM[7048] <= 32'b11100110100000111000001110010011;
ROM[7049] <= 32'b00000000111000111000001110110011;
ROM[7050] <= 32'b00000000011100010010000000100011;
ROM[7051] <= 32'b00000000010000010000000100010011;
ROM[7052] <= 32'b00000000001100010010000000100011;
ROM[7053] <= 32'b00000000010000010000000100010011;
ROM[7054] <= 32'b00000000010000010010000000100011;
ROM[7055] <= 32'b00000000010000010000000100010011;
ROM[7056] <= 32'b00000000010100010010000000100011;
ROM[7057] <= 32'b00000000010000010000000100010011;
ROM[7058] <= 32'b00000000011000010010000000100011;
ROM[7059] <= 32'b00000000010000010000000100010011;
ROM[7060] <= 32'b00000001010000000000001110010011;
ROM[7061] <= 32'b00000000100000111000001110010011;
ROM[7062] <= 32'b01000000011100010000001110110011;
ROM[7063] <= 32'b00000000011100000000001000110011;
ROM[7064] <= 32'b00000000001000000000000110110011;
ROM[7065] <= 32'b01010100100100100010000011101111;
ROM[7066] <= 32'b00000101111100000000001110010011;
ROM[7067] <= 32'b00000000011100010010000000100011;
ROM[7068] <= 32'b00000000010000010000000100010011;
ROM[7069] <= 32'b00000000000000000111001110110111;
ROM[7070] <= 32'b11101100000000111000001110010011;
ROM[7071] <= 32'b00000000111000111000001110110011;
ROM[7072] <= 32'b00000000011100010010000000100011;
ROM[7073] <= 32'b00000000010000010000000100010011;
ROM[7074] <= 32'b00000000001100010010000000100011;
ROM[7075] <= 32'b00000000010000010000000100010011;
ROM[7076] <= 32'b00000000010000010010000000100011;
ROM[7077] <= 32'b00000000010000010000000100010011;
ROM[7078] <= 32'b00000000010100010010000000100011;
ROM[7079] <= 32'b00000000010000010000000100010011;
ROM[7080] <= 32'b00000000011000010010000000100011;
ROM[7081] <= 32'b00000000010000010000000100010011;
ROM[7082] <= 32'b00000001010000000000001110010011;
ROM[7083] <= 32'b00000000100000111000001110010011;
ROM[7084] <= 32'b01000000011100010000001110110011;
ROM[7085] <= 32'b00000000011100000000001000110011;
ROM[7086] <= 32'b00000000001000000000000110110011;
ROM[7087] <= 32'b01001111000100100010000011101111;
ROM[7088] <= 32'b00000101111100000000001110010011;
ROM[7089] <= 32'b00000000011100010010000000100011;
ROM[7090] <= 32'b00000000010000010000000100010011;
ROM[7091] <= 32'b00000000000000000111001110110111;
ROM[7092] <= 32'b11110001100000111000001110010011;
ROM[7093] <= 32'b00000000111000111000001110110011;
ROM[7094] <= 32'b00000000011100010010000000100011;
ROM[7095] <= 32'b00000000010000010000000100010011;
ROM[7096] <= 32'b00000000001100010010000000100011;
ROM[7097] <= 32'b00000000010000010000000100010011;
ROM[7098] <= 32'b00000000010000010010000000100011;
ROM[7099] <= 32'b00000000010000010000000100010011;
ROM[7100] <= 32'b00000000010100010010000000100011;
ROM[7101] <= 32'b00000000010000010000000100010011;
ROM[7102] <= 32'b00000000011000010010000000100011;
ROM[7103] <= 32'b00000000010000010000000100010011;
ROM[7104] <= 32'b00000001010000000000001110010011;
ROM[7105] <= 32'b00000000100000111000001110010011;
ROM[7106] <= 32'b01000000011100010000001110110011;
ROM[7107] <= 32'b00000000011100000000001000110011;
ROM[7108] <= 32'b00000000001000000000000110110011;
ROM[7109] <= 32'b01001001100100100010000011101111;
ROM[7110] <= 32'b00000101111100000000001110010011;
ROM[7111] <= 32'b00000000011100010010000000100011;
ROM[7112] <= 32'b00000000010000010000000100010011;
ROM[7113] <= 32'b00000000000000000111001110110111;
ROM[7114] <= 32'b11110111000000111000001110010011;
ROM[7115] <= 32'b00000000111000111000001110110011;
ROM[7116] <= 32'b00000000011100010010000000100011;
ROM[7117] <= 32'b00000000010000010000000100010011;
ROM[7118] <= 32'b00000000001100010010000000100011;
ROM[7119] <= 32'b00000000010000010000000100010011;
ROM[7120] <= 32'b00000000010000010010000000100011;
ROM[7121] <= 32'b00000000010000010000000100010011;
ROM[7122] <= 32'b00000000010100010010000000100011;
ROM[7123] <= 32'b00000000010000010000000100010011;
ROM[7124] <= 32'b00000000011000010010000000100011;
ROM[7125] <= 32'b00000000010000010000000100010011;
ROM[7126] <= 32'b00000001010000000000001110010011;
ROM[7127] <= 32'b00000000100000111000001110010011;
ROM[7128] <= 32'b01000000011100010000001110110011;
ROM[7129] <= 32'b00000000011100000000001000110011;
ROM[7130] <= 32'b00000000001000000000000110110011;
ROM[7131] <= 32'b01000100000100100010000011101111;
ROM[7132] <= 32'b00000101111100000000001110010011;
ROM[7133] <= 32'b00000000011100010010000000100011;
ROM[7134] <= 32'b00000000010000010000000100010011;
ROM[7135] <= 32'b00000000000000000111001110110111;
ROM[7136] <= 32'b11111100100000111000001110010011;
ROM[7137] <= 32'b00000000111000111000001110110011;
ROM[7138] <= 32'b00000000011100010010000000100011;
ROM[7139] <= 32'b00000000010000010000000100010011;
ROM[7140] <= 32'b00000000001100010010000000100011;
ROM[7141] <= 32'b00000000010000010000000100010011;
ROM[7142] <= 32'b00000000010000010010000000100011;
ROM[7143] <= 32'b00000000010000010000000100010011;
ROM[7144] <= 32'b00000000010100010010000000100011;
ROM[7145] <= 32'b00000000010000010000000100010011;
ROM[7146] <= 32'b00000000011000010010000000100011;
ROM[7147] <= 32'b00000000010000010000000100010011;
ROM[7148] <= 32'b00000001010000000000001110010011;
ROM[7149] <= 32'b00000000100000111000001110010011;
ROM[7150] <= 32'b01000000011100010000001110110011;
ROM[7151] <= 32'b00000000011100000000001000110011;
ROM[7152] <= 32'b00000000001000000000000110110011;
ROM[7153] <= 32'b00111110100100100010000011101111;
ROM[7154] <= 32'b00000101111100000000001110010011;
ROM[7155] <= 32'b00000000011100010010000000100011;
ROM[7156] <= 32'b00000000010000010000000100010011;
ROM[7157] <= 32'b00000000000000000111001110110111;
ROM[7158] <= 32'b00000010000000111000001110010011;
ROM[7159] <= 32'b00000000111000111000001110110011;
ROM[7160] <= 32'b00000000011100010010000000100011;
ROM[7161] <= 32'b00000000010000010000000100010011;
ROM[7162] <= 32'b00000000001100010010000000100011;
ROM[7163] <= 32'b00000000010000010000000100010011;
ROM[7164] <= 32'b00000000010000010010000000100011;
ROM[7165] <= 32'b00000000010000010000000100010011;
ROM[7166] <= 32'b00000000010100010010000000100011;
ROM[7167] <= 32'b00000000010000010000000100010011;
ROM[7168] <= 32'b00000000011000010010000000100011;
ROM[7169] <= 32'b00000000010000010000000100010011;
ROM[7170] <= 32'b00000001010000000000001110010011;
ROM[7171] <= 32'b00000000100000111000001110010011;
ROM[7172] <= 32'b01000000011100010000001110110011;
ROM[7173] <= 32'b00000000011100000000001000110011;
ROM[7174] <= 32'b00000000001000000000000110110011;
ROM[7175] <= 32'b00111001000100100010000011101111;
ROM[7176] <= 32'b11111111110000010000000100010011;
ROM[7177] <= 32'b00000000000000010010001110000011;
ROM[7178] <= 32'b00000000011100011010110000100011;
ROM[7179] <= 32'b00110010100000000000000011101111;
ROM[7180] <= 32'b00000000100000000000001110010011;
ROM[7181] <= 32'b00000000011100010010000000100011;
ROM[7182] <= 32'b00000000010000010000000100010011;
ROM[7183] <= 32'b00000000000000000111001110110111;
ROM[7184] <= 32'b00001000100000111000001110010011;
ROM[7185] <= 32'b00000000111000111000001110110011;
ROM[7186] <= 32'b00000000011100010010000000100011;
ROM[7187] <= 32'b00000000010000010000000100010011;
ROM[7188] <= 32'b00000000001100010010000000100011;
ROM[7189] <= 32'b00000000010000010000000100010011;
ROM[7190] <= 32'b00000000010000010010000000100011;
ROM[7191] <= 32'b00000000010000010000000100010011;
ROM[7192] <= 32'b00000000010100010010000000100011;
ROM[7193] <= 32'b00000000010000010000000100010011;
ROM[7194] <= 32'b00000000011000010010000000100011;
ROM[7195] <= 32'b00000000010000010000000100010011;
ROM[7196] <= 32'b00000001010000000000001110010011;
ROM[7197] <= 32'b00000000010000111000001110010011;
ROM[7198] <= 32'b01000000011100010000001110110011;
ROM[7199] <= 32'b00000000011100000000001000110011;
ROM[7200] <= 32'b00000000001000000000000110110011;
ROM[7201] <= 32'b01101011100000100010000011101111;
ROM[7202] <= 32'b00000101111100000000001110010011;
ROM[7203] <= 32'b00000000011100010010000000100011;
ROM[7204] <= 32'b00000000010000010000000100010011;
ROM[7205] <= 32'b00000000000000000111001110110111;
ROM[7206] <= 32'b00001110000000111000001110010011;
ROM[7207] <= 32'b00000000111000111000001110110011;
ROM[7208] <= 32'b00000000011100010010000000100011;
ROM[7209] <= 32'b00000000010000010000000100010011;
ROM[7210] <= 32'b00000000001100010010000000100011;
ROM[7211] <= 32'b00000000010000010000000100010011;
ROM[7212] <= 32'b00000000010000010010000000100011;
ROM[7213] <= 32'b00000000010000010000000100010011;
ROM[7214] <= 32'b00000000010100010010000000100011;
ROM[7215] <= 32'b00000000010000010000000100010011;
ROM[7216] <= 32'b00000000011000010010000000100011;
ROM[7217] <= 32'b00000000010000010000000100010011;
ROM[7218] <= 32'b00000001010000000000001110010011;
ROM[7219] <= 32'b00000000100000111000001110010011;
ROM[7220] <= 32'b01000000011100010000001110110011;
ROM[7221] <= 32'b00000000011100000000001000110011;
ROM[7222] <= 32'b00000000001000000000000110110011;
ROM[7223] <= 32'b00101101000100100010000011101111;
ROM[7224] <= 32'b00000101111100000000001110010011;
ROM[7225] <= 32'b00000000011100010010000000100011;
ROM[7226] <= 32'b00000000010000010000000100010011;
ROM[7227] <= 32'b00000000000000000111001110110111;
ROM[7228] <= 32'b00010011100000111000001110010011;
ROM[7229] <= 32'b00000000111000111000001110110011;
ROM[7230] <= 32'b00000000011100010010000000100011;
ROM[7231] <= 32'b00000000010000010000000100010011;
ROM[7232] <= 32'b00000000001100010010000000100011;
ROM[7233] <= 32'b00000000010000010000000100010011;
ROM[7234] <= 32'b00000000010000010010000000100011;
ROM[7235] <= 32'b00000000010000010000000100010011;
ROM[7236] <= 32'b00000000010100010010000000100011;
ROM[7237] <= 32'b00000000010000010000000100010011;
ROM[7238] <= 32'b00000000011000010010000000100011;
ROM[7239] <= 32'b00000000010000010000000100010011;
ROM[7240] <= 32'b00000001010000000000001110010011;
ROM[7241] <= 32'b00000000100000111000001110010011;
ROM[7242] <= 32'b01000000011100010000001110110011;
ROM[7243] <= 32'b00000000011100000000001000110011;
ROM[7244] <= 32'b00000000001000000000000110110011;
ROM[7245] <= 32'b00100111100100100010000011101111;
ROM[7246] <= 32'b00000101111100000000001110010011;
ROM[7247] <= 32'b00000000011100010010000000100011;
ROM[7248] <= 32'b00000000010000010000000100010011;
ROM[7249] <= 32'b00000000000000000111001110110111;
ROM[7250] <= 32'b00011001000000111000001110010011;
ROM[7251] <= 32'b00000000111000111000001110110011;
ROM[7252] <= 32'b00000000011100010010000000100011;
ROM[7253] <= 32'b00000000010000010000000100010011;
ROM[7254] <= 32'b00000000001100010010000000100011;
ROM[7255] <= 32'b00000000010000010000000100010011;
ROM[7256] <= 32'b00000000010000010010000000100011;
ROM[7257] <= 32'b00000000010000010000000100010011;
ROM[7258] <= 32'b00000000010100010010000000100011;
ROM[7259] <= 32'b00000000010000010000000100010011;
ROM[7260] <= 32'b00000000011000010010000000100011;
ROM[7261] <= 32'b00000000010000010000000100010011;
ROM[7262] <= 32'b00000001010000000000001110010011;
ROM[7263] <= 32'b00000000100000111000001110010011;
ROM[7264] <= 32'b01000000011100010000001110110011;
ROM[7265] <= 32'b00000000011100000000001000110011;
ROM[7266] <= 32'b00000000001000000000000110110011;
ROM[7267] <= 32'b00100010000100100010000011101111;
ROM[7268] <= 32'b00000101111100000000001110010011;
ROM[7269] <= 32'b00000000011100010010000000100011;
ROM[7270] <= 32'b00000000010000010000000100010011;
ROM[7271] <= 32'b00000000000000000111001110110111;
ROM[7272] <= 32'b00011110100000111000001110010011;
ROM[7273] <= 32'b00000000111000111000001110110011;
ROM[7274] <= 32'b00000000011100010010000000100011;
ROM[7275] <= 32'b00000000010000010000000100010011;
ROM[7276] <= 32'b00000000001100010010000000100011;
ROM[7277] <= 32'b00000000010000010000000100010011;
ROM[7278] <= 32'b00000000010000010010000000100011;
ROM[7279] <= 32'b00000000010000010000000100010011;
ROM[7280] <= 32'b00000000010100010010000000100011;
ROM[7281] <= 32'b00000000010000010000000100010011;
ROM[7282] <= 32'b00000000011000010010000000100011;
ROM[7283] <= 32'b00000000010000010000000100010011;
ROM[7284] <= 32'b00000001010000000000001110010011;
ROM[7285] <= 32'b00000000100000111000001110010011;
ROM[7286] <= 32'b01000000011100010000001110110011;
ROM[7287] <= 32'b00000000011100000000001000110011;
ROM[7288] <= 32'b00000000001000000000000110110011;
ROM[7289] <= 32'b00011100100100100010000011101111;
ROM[7290] <= 32'b00000101111100000000001110010011;
ROM[7291] <= 32'b00000000011100010010000000100011;
ROM[7292] <= 32'b00000000010000010000000100010011;
ROM[7293] <= 32'b00000000000000000111001110110111;
ROM[7294] <= 32'b00100100000000111000001110010011;
ROM[7295] <= 32'b00000000111000111000001110110011;
ROM[7296] <= 32'b00000000011100010010000000100011;
ROM[7297] <= 32'b00000000010000010000000100010011;
ROM[7298] <= 32'b00000000001100010010000000100011;
ROM[7299] <= 32'b00000000010000010000000100010011;
ROM[7300] <= 32'b00000000010000010010000000100011;
ROM[7301] <= 32'b00000000010000010000000100010011;
ROM[7302] <= 32'b00000000010100010010000000100011;
ROM[7303] <= 32'b00000000010000010000000100010011;
ROM[7304] <= 32'b00000000011000010010000000100011;
ROM[7305] <= 32'b00000000010000010000000100010011;
ROM[7306] <= 32'b00000001010000000000001110010011;
ROM[7307] <= 32'b00000000100000111000001110010011;
ROM[7308] <= 32'b01000000011100010000001110110011;
ROM[7309] <= 32'b00000000011100000000001000110011;
ROM[7310] <= 32'b00000000001000000000000110110011;
ROM[7311] <= 32'b00010111000100100010000011101111;
ROM[7312] <= 32'b00000101111100000000001110010011;
ROM[7313] <= 32'b00000000011100010010000000100011;
ROM[7314] <= 32'b00000000010000010000000100010011;
ROM[7315] <= 32'b00000000000000000111001110110111;
ROM[7316] <= 32'b00101001100000111000001110010011;
ROM[7317] <= 32'b00000000111000111000001110110011;
ROM[7318] <= 32'b00000000011100010010000000100011;
ROM[7319] <= 32'b00000000010000010000000100010011;
ROM[7320] <= 32'b00000000001100010010000000100011;
ROM[7321] <= 32'b00000000010000010000000100010011;
ROM[7322] <= 32'b00000000010000010010000000100011;
ROM[7323] <= 32'b00000000010000010000000100010011;
ROM[7324] <= 32'b00000000010100010010000000100011;
ROM[7325] <= 32'b00000000010000010000000100010011;
ROM[7326] <= 32'b00000000011000010010000000100011;
ROM[7327] <= 32'b00000000010000010000000100010011;
ROM[7328] <= 32'b00000001010000000000001110010011;
ROM[7329] <= 32'b00000000100000111000001110010011;
ROM[7330] <= 32'b01000000011100010000001110110011;
ROM[7331] <= 32'b00000000011100000000001000110011;
ROM[7332] <= 32'b00000000001000000000000110110011;
ROM[7333] <= 32'b00010001100100100010000011101111;
ROM[7334] <= 32'b00000101111100000000001110010011;
ROM[7335] <= 32'b00000000011100010010000000100011;
ROM[7336] <= 32'b00000000010000010000000100010011;
ROM[7337] <= 32'b00000000000000000111001110110111;
ROM[7338] <= 32'b00101111000000111000001110010011;
ROM[7339] <= 32'b00000000111000111000001110110011;
ROM[7340] <= 32'b00000000011100010010000000100011;
ROM[7341] <= 32'b00000000010000010000000100010011;
ROM[7342] <= 32'b00000000001100010010000000100011;
ROM[7343] <= 32'b00000000010000010000000100010011;
ROM[7344] <= 32'b00000000010000010010000000100011;
ROM[7345] <= 32'b00000000010000010000000100010011;
ROM[7346] <= 32'b00000000010100010010000000100011;
ROM[7347] <= 32'b00000000010000010000000100010011;
ROM[7348] <= 32'b00000000011000010010000000100011;
ROM[7349] <= 32'b00000000010000010000000100010011;
ROM[7350] <= 32'b00000001010000000000001110010011;
ROM[7351] <= 32'b00000000100000111000001110010011;
ROM[7352] <= 32'b01000000011100010000001110110011;
ROM[7353] <= 32'b00000000011100000000001000110011;
ROM[7354] <= 32'b00000000001000000000000110110011;
ROM[7355] <= 32'b00001100000100100010000011101111;
ROM[7356] <= 32'b00000101111100000000001110010011;
ROM[7357] <= 32'b00000000011100010010000000100011;
ROM[7358] <= 32'b00000000010000010000000100010011;
ROM[7359] <= 32'b00000000000000000111001110110111;
ROM[7360] <= 32'b00110100100000111000001110010011;
ROM[7361] <= 32'b00000000111000111000001110110011;
ROM[7362] <= 32'b00000000011100010010000000100011;
ROM[7363] <= 32'b00000000010000010000000100010011;
ROM[7364] <= 32'b00000000001100010010000000100011;
ROM[7365] <= 32'b00000000010000010000000100010011;
ROM[7366] <= 32'b00000000010000010010000000100011;
ROM[7367] <= 32'b00000000010000010000000100010011;
ROM[7368] <= 32'b00000000010100010010000000100011;
ROM[7369] <= 32'b00000000010000010000000100010011;
ROM[7370] <= 32'b00000000011000010010000000100011;
ROM[7371] <= 32'b00000000010000010000000100010011;
ROM[7372] <= 32'b00000001010000000000001110010011;
ROM[7373] <= 32'b00000000100000111000001110010011;
ROM[7374] <= 32'b01000000011100010000001110110011;
ROM[7375] <= 32'b00000000011100000000001000110011;
ROM[7376] <= 32'b00000000001000000000000110110011;
ROM[7377] <= 32'b00000110100100100010000011101111;
ROM[7378] <= 32'b11111111110000010000000100010011;
ROM[7379] <= 32'b00000000000000010010001110000011;
ROM[7380] <= 32'b00000000011100011010110000100011;
ROM[7381] <= 32'b01000011000000000000000011101111;
ROM[7382] <= 32'b00000000101100000000001110010011;
ROM[7383] <= 32'b00000000011100010010000000100011;
ROM[7384] <= 32'b00000000010000010000000100010011;
ROM[7385] <= 32'b00000000000000000111001110110111;
ROM[7386] <= 32'b00111011000000111000001110010011;
ROM[7387] <= 32'b00000000111000111000001110110011;
ROM[7388] <= 32'b00000000011100010010000000100011;
ROM[7389] <= 32'b00000000010000010000000100010011;
ROM[7390] <= 32'b00000000001100010010000000100011;
ROM[7391] <= 32'b00000000010000010000000100010011;
ROM[7392] <= 32'b00000000010000010010000000100011;
ROM[7393] <= 32'b00000000010000010000000100010011;
ROM[7394] <= 32'b00000000010100010010000000100011;
ROM[7395] <= 32'b00000000010000010000000100010011;
ROM[7396] <= 32'b00000000011000010010000000100011;
ROM[7397] <= 32'b00000000010000010000000100010011;
ROM[7398] <= 32'b00000001010000000000001110010011;
ROM[7399] <= 32'b00000000010000111000001110010011;
ROM[7400] <= 32'b01000000011100010000001110110011;
ROM[7401] <= 32'b00000000011100000000001000110011;
ROM[7402] <= 32'b00000000001000000000000110110011;
ROM[7403] <= 32'b00111001000000100010000011101111;
ROM[7404] <= 32'b00000101111100000000001110010011;
ROM[7405] <= 32'b00000000011100010010000000100011;
ROM[7406] <= 32'b00000000010000010000000100010011;
ROM[7407] <= 32'b00000000000000000111001110110111;
ROM[7408] <= 32'b01000000100000111000001110010011;
ROM[7409] <= 32'b00000000111000111000001110110011;
ROM[7410] <= 32'b00000000011100010010000000100011;
ROM[7411] <= 32'b00000000010000010000000100010011;
ROM[7412] <= 32'b00000000001100010010000000100011;
ROM[7413] <= 32'b00000000010000010000000100010011;
ROM[7414] <= 32'b00000000010000010010000000100011;
ROM[7415] <= 32'b00000000010000010000000100010011;
ROM[7416] <= 32'b00000000010100010010000000100011;
ROM[7417] <= 32'b00000000010000010000000100010011;
ROM[7418] <= 32'b00000000011000010010000000100011;
ROM[7419] <= 32'b00000000010000010000000100010011;
ROM[7420] <= 32'b00000001010000000000001110010011;
ROM[7421] <= 32'b00000000100000111000001110010011;
ROM[7422] <= 32'b01000000011100010000001110110011;
ROM[7423] <= 32'b00000000011100000000001000110011;
ROM[7424] <= 32'b00000000001000000000000110110011;
ROM[7425] <= 32'b01111010100000100010000011101111;
ROM[7426] <= 32'b00000101111100000000001110010011;
ROM[7427] <= 32'b00000000011100010010000000100011;
ROM[7428] <= 32'b00000000010000010000000100010011;
ROM[7429] <= 32'b00000000000000000111001110110111;
ROM[7430] <= 32'b01000110000000111000001110010011;
ROM[7431] <= 32'b00000000111000111000001110110011;
ROM[7432] <= 32'b00000000011100010010000000100011;
ROM[7433] <= 32'b00000000010000010000000100010011;
ROM[7434] <= 32'b00000000001100010010000000100011;
ROM[7435] <= 32'b00000000010000010000000100010011;
ROM[7436] <= 32'b00000000010000010010000000100011;
ROM[7437] <= 32'b00000000010000010000000100010011;
ROM[7438] <= 32'b00000000010100010010000000100011;
ROM[7439] <= 32'b00000000010000010000000100010011;
ROM[7440] <= 32'b00000000011000010010000000100011;
ROM[7441] <= 32'b00000000010000010000000100010011;
ROM[7442] <= 32'b00000001010000000000001110010011;
ROM[7443] <= 32'b00000000100000111000001110010011;
ROM[7444] <= 32'b01000000011100010000001110110011;
ROM[7445] <= 32'b00000000011100000000001000110011;
ROM[7446] <= 32'b00000000001000000000000110110011;
ROM[7447] <= 32'b01110101000000100010000011101111;
ROM[7448] <= 32'b00000101111100000000001110010011;
ROM[7449] <= 32'b00000000011100010010000000100011;
ROM[7450] <= 32'b00000000010000010000000100010011;
ROM[7451] <= 32'b00000000000000000111001110110111;
ROM[7452] <= 32'b01001011100000111000001110010011;
ROM[7453] <= 32'b00000000111000111000001110110011;
ROM[7454] <= 32'b00000000011100010010000000100011;
ROM[7455] <= 32'b00000000010000010000000100010011;
ROM[7456] <= 32'b00000000001100010010000000100011;
ROM[7457] <= 32'b00000000010000010000000100010011;
ROM[7458] <= 32'b00000000010000010010000000100011;
ROM[7459] <= 32'b00000000010000010000000100010011;
ROM[7460] <= 32'b00000000010100010010000000100011;
ROM[7461] <= 32'b00000000010000010000000100010011;
ROM[7462] <= 32'b00000000011000010010000000100011;
ROM[7463] <= 32'b00000000010000010000000100010011;
ROM[7464] <= 32'b00000001010000000000001110010011;
ROM[7465] <= 32'b00000000100000111000001110010011;
ROM[7466] <= 32'b01000000011100010000001110110011;
ROM[7467] <= 32'b00000000011100000000001000110011;
ROM[7468] <= 32'b00000000001000000000000110110011;
ROM[7469] <= 32'b01101111100000100010000011101111;
ROM[7470] <= 32'b00000101111100000000001110010011;
ROM[7471] <= 32'b00000000011100010010000000100011;
ROM[7472] <= 32'b00000000010000010000000100010011;
ROM[7473] <= 32'b00000000000000000111001110110111;
ROM[7474] <= 32'b01010001000000111000001110010011;
ROM[7475] <= 32'b00000000111000111000001110110011;
ROM[7476] <= 32'b00000000011100010010000000100011;
ROM[7477] <= 32'b00000000010000010000000100010011;
ROM[7478] <= 32'b00000000001100010010000000100011;
ROM[7479] <= 32'b00000000010000010000000100010011;
ROM[7480] <= 32'b00000000010000010010000000100011;
ROM[7481] <= 32'b00000000010000010000000100010011;
ROM[7482] <= 32'b00000000010100010010000000100011;
ROM[7483] <= 32'b00000000010000010000000100010011;
ROM[7484] <= 32'b00000000011000010010000000100011;
ROM[7485] <= 32'b00000000010000010000000100010011;
ROM[7486] <= 32'b00000001010000000000001110010011;
ROM[7487] <= 32'b00000000100000111000001110010011;
ROM[7488] <= 32'b01000000011100010000001110110011;
ROM[7489] <= 32'b00000000011100000000001000110011;
ROM[7490] <= 32'b00000000001000000000000110110011;
ROM[7491] <= 32'b01101010000000100010000011101111;
ROM[7492] <= 32'b00000101111100000000001110010011;
ROM[7493] <= 32'b00000000011100010010000000100011;
ROM[7494] <= 32'b00000000010000010000000100010011;
ROM[7495] <= 32'b00000000000000000111001110110111;
ROM[7496] <= 32'b01010110100000111000001110010011;
ROM[7497] <= 32'b00000000111000111000001110110011;
ROM[7498] <= 32'b00000000011100010010000000100011;
ROM[7499] <= 32'b00000000010000010000000100010011;
ROM[7500] <= 32'b00000000001100010010000000100011;
ROM[7501] <= 32'b00000000010000010000000100010011;
ROM[7502] <= 32'b00000000010000010010000000100011;
ROM[7503] <= 32'b00000000010000010000000100010011;
ROM[7504] <= 32'b00000000010100010010000000100011;
ROM[7505] <= 32'b00000000010000010000000100010011;
ROM[7506] <= 32'b00000000011000010010000000100011;
ROM[7507] <= 32'b00000000010000010000000100010011;
ROM[7508] <= 32'b00000001010000000000001110010011;
ROM[7509] <= 32'b00000000100000111000001110010011;
ROM[7510] <= 32'b01000000011100010000001110110011;
ROM[7511] <= 32'b00000000011100000000001000110011;
ROM[7512] <= 32'b00000000001000000000000110110011;
ROM[7513] <= 32'b01100100100000100010000011101111;
ROM[7514] <= 32'b00000101111100000000001110010011;
ROM[7515] <= 32'b00000000011100010010000000100011;
ROM[7516] <= 32'b00000000010000010000000100010011;
ROM[7517] <= 32'b00000000000000000111001110110111;
ROM[7518] <= 32'b01011100000000111000001110010011;
ROM[7519] <= 32'b00000000111000111000001110110011;
ROM[7520] <= 32'b00000000011100010010000000100011;
ROM[7521] <= 32'b00000000010000010000000100010011;
ROM[7522] <= 32'b00000000001100010010000000100011;
ROM[7523] <= 32'b00000000010000010000000100010011;
ROM[7524] <= 32'b00000000010000010010000000100011;
ROM[7525] <= 32'b00000000010000010000000100010011;
ROM[7526] <= 32'b00000000010100010010000000100011;
ROM[7527] <= 32'b00000000010000010000000100010011;
ROM[7528] <= 32'b00000000011000010010000000100011;
ROM[7529] <= 32'b00000000010000010000000100010011;
ROM[7530] <= 32'b00000001010000000000001110010011;
ROM[7531] <= 32'b00000000100000111000001110010011;
ROM[7532] <= 32'b01000000011100010000001110110011;
ROM[7533] <= 32'b00000000011100000000001000110011;
ROM[7534] <= 32'b00000000001000000000000110110011;
ROM[7535] <= 32'b01011111000000100010000011101111;
ROM[7536] <= 32'b00000101111100000000001110010011;
ROM[7537] <= 32'b00000000011100010010000000100011;
ROM[7538] <= 32'b00000000010000010000000100010011;
ROM[7539] <= 32'b00000000000000000111001110110111;
ROM[7540] <= 32'b01100001100000111000001110010011;
ROM[7541] <= 32'b00000000111000111000001110110011;
ROM[7542] <= 32'b00000000011100010010000000100011;
ROM[7543] <= 32'b00000000010000010000000100010011;
ROM[7544] <= 32'b00000000001100010010000000100011;
ROM[7545] <= 32'b00000000010000010000000100010011;
ROM[7546] <= 32'b00000000010000010010000000100011;
ROM[7547] <= 32'b00000000010000010000000100010011;
ROM[7548] <= 32'b00000000010100010010000000100011;
ROM[7549] <= 32'b00000000010000010000000100010011;
ROM[7550] <= 32'b00000000011000010010000000100011;
ROM[7551] <= 32'b00000000010000010000000100010011;
ROM[7552] <= 32'b00000001010000000000001110010011;
ROM[7553] <= 32'b00000000100000111000001110010011;
ROM[7554] <= 32'b01000000011100010000001110110011;
ROM[7555] <= 32'b00000000011100000000001000110011;
ROM[7556] <= 32'b00000000001000000000000110110011;
ROM[7557] <= 32'b01011001100000100010000011101111;
ROM[7558] <= 32'b00000101111100000000001110010011;
ROM[7559] <= 32'b00000000011100010010000000100011;
ROM[7560] <= 32'b00000000010000010000000100010011;
ROM[7561] <= 32'b00000000000000000111001110110111;
ROM[7562] <= 32'b01100111000000111000001110010011;
ROM[7563] <= 32'b00000000111000111000001110110011;
ROM[7564] <= 32'b00000000011100010010000000100011;
ROM[7565] <= 32'b00000000010000010000000100010011;
ROM[7566] <= 32'b00000000001100010010000000100011;
ROM[7567] <= 32'b00000000010000010000000100010011;
ROM[7568] <= 32'b00000000010000010010000000100011;
ROM[7569] <= 32'b00000000010000010000000100010011;
ROM[7570] <= 32'b00000000010100010010000000100011;
ROM[7571] <= 32'b00000000010000010000000100010011;
ROM[7572] <= 32'b00000000011000010010000000100011;
ROM[7573] <= 32'b00000000010000010000000100010011;
ROM[7574] <= 32'b00000001010000000000001110010011;
ROM[7575] <= 32'b00000000100000111000001110010011;
ROM[7576] <= 32'b01000000011100010000001110110011;
ROM[7577] <= 32'b00000000011100000000001000110011;
ROM[7578] <= 32'b00000000001000000000000110110011;
ROM[7579] <= 32'b01010100000000100010000011101111;
ROM[7580] <= 32'b00000101111100000000001110010011;
ROM[7581] <= 32'b00000000011100010010000000100011;
ROM[7582] <= 32'b00000000010000010000000100010011;
ROM[7583] <= 32'b00000000000000000111001110110111;
ROM[7584] <= 32'b01101100100000111000001110010011;
ROM[7585] <= 32'b00000000111000111000001110110011;
ROM[7586] <= 32'b00000000011100010010000000100011;
ROM[7587] <= 32'b00000000010000010000000100010011;
ROM[7588] <= 32'b00000000001100010010000000100011;
ROM[7589] <= 32'b00000000010000010000000100010011;
ROM[7590] <= 32'b00000000010000010010000000100011;
ROM[7591] <= 32'b00000000010000010000000100010011;
ROM[7592] <= 32'b00000000010100010010000000100011;
ROM[7593] <= 32'b00000000010000010000000100010011;
ROM[7594] <= 32'b00000000011000010010000000100011;
ROM[7595] <= 32'b00000000010000010000000100010011;
ROM[7596] <= 32'b00000001010000000000001110010011;
ROM[7597] <= 32'b00000000100000111000001110010011;
ROM[7598] <= 32'b01000000011100010000001110110011;
ROM[7599] <= 32'b00000000011100000000001000110011;
ROM[7600] <= 32'b00000000001000000000000110110011;
ROM[7601] <= 32'b01001110100000100010000011101111;
ROM[7602] <= 32'b00000101111100000000001110010011;
ROM[7603] <= 32'b00000000011100010010000000100011;
ROM[7604] <= 32'b00000000010000010000000100010011;
ROM[7605] <= 32'b00000000000000000111001110110111;
ROM[7606] <= 32'b01110010000000111000001110010011;
ROM[7607] <= 32'b00000000111000111000001110110011;
ROM[7608] <= 32'b00000000011100010010000000100011;
ROM[7609] <= 32'b00000000010000010000000100010011;
ROM[7610] <= 32'b00000000001100010010000000100011;
ROM[7611] <= 32'b00000000010000010000000100010011;
ROM[7612] <= 32'b00000000010000010010000000100011;
ROM[7613] <= 32'b00000000010000010000000100010011;
ROM[7614] <= 32'b00000000010100010010000000100011;
ROM[7615] <= 32'b00000000010000010000000100010011;
ROM[7616] <= 32'b00000000011000010010000000100011;
ROM[7617] <= 32'b00000000010000010000000100010011;
ROM[7618] <= 32'b00000001010000000000001110010011;
ROM[7619] <= 32'b00000000100000111000001110010011;
ROM[7620] <= 32'b01000000011100010000001110110011;
ROM[7621] <= 32'b00000000011100000000001000110011;
ROM[7622] <= 32'b00000000001000000000000110110011;
ROM[7623] <= 32'b01001001000000100010000011101111;
ROM[7624] <= 32'b00000101111100000000001110010011;
ROM[7625] <= 32'b00000000011100010010000000100011;
ROM[7626] <= 32'b00000000010000010000000100010011;
ROM[7627] <= 32'b00000000000000000111001110110111;
ROM[7628] <= 32'b01110111100000111000001110010011;
ROM[7629] <= 32'b00000000111000111000001110110011;
ROM[7630] <= 32'b00000000011100010010000000100011;
ROM[7631] <= 32'b00000000010000010000000100010011;
ROM[7632] <= 32'b00000000001100010010000000100011;
ROM[7633] <= 32'b00000000010000010000000100010011;
ROM[7634] <= 32'b00000000010000010010000000100011;
ROM[7635] <= 32'b00000000010000010000000100010011;
ROM[7636] <= 32'b00000000010100010010000000100011;
ROM[7637] <= 32'b00000000010000010000000100010011;
ROM[7638] <= 32'b00000000011000010010000000100011;
ROM[7639] <= 32'b00000000010000010000000100010011;
ROM[7640] <= 32'b00000001010000000000001110010011;
ROM[7641] <= 32'b00000000100000111000001110010011;
ROM[7642] <= 32'b01000000011100010000001110110011;
ROM[7643] <= 32'b00000000011100000000001000110011;
ROM[7644] <= 32'b00000000001000000000000110110011;
ROM[7645] <= 32'b01000011100000100010000011101111;
ROM[7646] <= 32'b11111111110000010000000100010011;
ROM[7647] <= 32'b00000000000000010010001110000011;
ROM[7648] <= 32'b00000000011100011010110000100011;
ROM[7649] <= 32'b00011100100000000000000011101111;
ROM[7650] <= 32'b00000000010000000000001110010011;
ROM[7651] <= 32'b00000000011100010010000000100011;
ROM[7652] <= 32'b00000000010000010000000100010011;
ROM[7653] <= 32'b00000000000000000111001110110111;
ROM[7654] <= 32'b01111110000000111000001110010011;
ROM[7655] <= 32'b00000000111000111000001110110011;
ROM[7656] <= 32'b00000000011100010010000000100011;
ROM[7657] <= 32'b00000000010000010000000100010011;
ROM[7658] <= 32'b00000000001100010010000000100011;
ROM[7659] <= 32'b00000000010000010000000100010011;
ROM[7660] <= 32'b00000000010000010010000000100011;
ROM[7661] <= 32'b00000000010000010000000100010011;
ROM[7662] <= 32'b00000000010100010010000000100011;
ROM[7663] <= 32'b00000000010000010000000100010011;
ROM[7664] <= 32'b00000000011000010010000000100011;
ROM[7665] <= 32'b00000000010000010000000100010011;
ROM[7666] <= 32'b00000001010000000000001110010011;
ROM[7667] <= 32'b00000000010000111000001110010011;
ROM[7668] <= 32'b01000000011100010000001110110011;
ROM[7669] <= 32'b00000000011100000000001000110011;
ROM[7670] <= 32'b00000000001000000000000110110011;
ROM[7671] <= 32'b01110110000100100001000011101111;
ROM[7672] <= 32'b00000101111100000000001110010011;
ROM[7673] <= 32'b00000000011100010010000000100011;
ROM[7674] <= 32'b00000000010000010000000100010011;
ROM[7675] <= 32'b00000000000000001000001110110111;
ROM[7676] <= 32'b10000011100000111000001110010011;
ROM[7677] <= 32'b00000000111000111000001110110011;
ROM[7678] <= 32'b00000000011100010010000000100011;
ROM[7679] <= 32'b00000000010000010000000100010011;
ROM[7680] <= 32'b00000000001100010010000000100011;
ROM[7681] <= 32'b00000000010000010000000100010011;
ROM[7682] <= 32'b00000000010000010010000000100011;
ROM[7683] <= 32'b00000000010000010000000100010011;
ROM[7684] <= 32'b00000000010100010010000000100011;
ROM[7685] <= 32'b00000000010000010000000100010011;
ROM[7686] <= 32'b00000000011000010010000000100011;
ROM[7687] <= 32'b00000000010000010000000100010011;
ROM[7688] <= 32'b00000001010000000000001110010011;
ROM[7689] <= 32'b00000000100000111000001110010011;
ROM[7690] <= 32'b01000000011100010000001110110011;
ROM[7691] <= 32'b00000000011100000000001000110011;
ROM[7692] <= 32'b00000000001000000000000110110011;
ROM[7693] <= 32'b00110111100000100010000011101111;
ROM[7694] <= 32'b00000101111100000000001110010011;
ROM[7695] <= 32'b00000000011100010010000000100011;
ROM[7696] <= 32'b00000000010000010000000100010011;
ROM[7697] <= 32'b00000000000000001000001110110111;
ROM[7698] <= 32'b10001001000000111000001110010011;
ROM[7699] <= 32'b00000000111000111000001110110011;
ROM[7700] <= 32'b00000000011100010010000000100011;
ROM[7701] <= 32'b00000000010000010000000100010011;
ROM[7702] <= 32'b00000000001100010010000000100011;
ROM[7703] <= 32'b00000000010000010000000100010011;
ROM[7704] <= 32'b00000000010000010010000000100011;
ROM[7705] <= 32'b00000000010000010000000100010011;
ROM[7706] <= 32'b00000000010100010010000000100011;
ROM[7707] <= 32'b00000000010000010000000100010011;
ROM[7708] <= 32'b00000000011000010010000000100011;
ROM[7709] <= 32'b00000000010000010000000100010011;
ROM[7710] <= 32'b00000001010000000000001110010011;
ROM[7711] <= 32'b00000000100000111000001110010011;
ROM[7712] <= 32'b01000000011100010000001110110011;
ROM[7713] <= 32'b00000000011100000000001000110011;
ROM[7714] <= 32'b00000000001000000000000110110011;
ROM[7715] <= 32'b00110010000000100010000011101111;
ROM[7716] <= 32'b00000101111100000000001110010011;
ROM[7717] <= 32'b00000000011100010010000000100011;
ROM[7718] <= 32'b00000000010000010000000100010011;
ROM[7719] <= 32'b00000000000000001000001110110111;
ROM[7720] <= 32'b10001110100000111000001110010011;
ROM[7721] <= 32'b00000000111000111000001110110011;
ROM[7722] <= 32'b00000000011100010010000000100011;
ROM[7723] <= 32'b00000000010000010000000100010011;
ROM[7724] <= 32'b00000000001100010010000000100011;
ROM[7725] <= 32'b00000000010000010000000100010011;
ROM[7726] <= 32'b00000000010000010010000000100011;
ROM[7727] <= 32'b00000000010000010000000100010011;
ROM[7728] <= 32'b00000000010100010010000000100011;
ROM[7729] <= 32'b00000000010000010000000100010011;
ROM[7730] <= 32'b00000000011000010010000000100011;
ROM[7731] <= 32'b00000000010000010000000100010011;
ROM[7732] <= 32'b00000001010000000000001110010011;
ROM[7733] <= 32'b00000000100000111000001110010011;
ROM[7734] <= 32'b01000000011100010000001110110011;
ROM[7735] <= 32'b00000000011100000000001000110011;
ROM[7736] <= 32'b00000000001000000000000110110011;
ROM[7737] <= 32'b00101100100000100010000011101111;
ROM[7738] <= 32'b00000101111100000000001110010011;
ROM[7739] <= 32'b00000000011100010010000000100011;
ROM[7740] <= 32'b00000000010000010000000100010011;
ROM[7741] <= 32'b00000000000000001000001110110111;
ROM[7742] <= 32'b10010100000000111000001110010011;
ROM[7743] <= 32'b00000000111000111000001110110011;
ROM[7744] <= 32'b00000000011100010010000000100011;
ROM[7745] <= 32'b00000000010000010000000100010011;
ROM[7746] <= 32'b00000000001100010010000000100011;
ROM[7747] <= 32'b00000000010000010000000100010011;
ROM[7748] <= 32'b00000000010000010010000000100011;
ROM[7749] <= 32'b00000000010000010000000100010011;
ROM[7750] <= 32'b00000000010100010010000000100011;
ROM[7751] <= 32'b00000000010000010000000100010011;
ROM[7752] <= 32'b00000000011000010010000000100011;
ROM[7753] <= 32'b00000000010000010000000100010011;
ROM[7754] <= 32'b00000001010000000000001110010011;
ROM[7755] <= 32'b00000000100000111000001110010011;
ROM[7756] <= 32'b01000000011100010000001110110011;
ROM[7757] <= 32'b00000000011100000000001000110011;
ROM[7758] <= 32'b00000000001000000000000110110011;
ROM[7759] <= 32'b00100111000000100010000011101111;
ROM[7760] <= 32'b11111111110000010000000100010011;
ROM[7761] <= 32'b00000000000000010010001110000011;
ROM[7762] <= 32'b00000000011100011010110000100011;
ROM[7763] <= 32'b00000000000000000000001110010011;
ROM[7764] <= 32'b00000000011100010010000000100011;
ROM[7765] <= 32'b00000000010000010000000100010011;
ROM[7766] <= 32'b11111111110000010000000100010011;
ROM[7767] <= 32'b00000000000000010010001110000011;
ROM[7768] <= 32'b00000010011100011010000000100011;
ROM[7769] <= 32'b00000010000000011010001110000011;
ROM[7770] <= 32'b00000000011100010010000000100011;
ROM[7771] <= 32'b00000000010000010000000100010011;
ROM[7772] <= 32'b00000000000000000000001110010011;
ROM[7773] <= 32'b00000000011100010010000000100011;
ROM[7774] <= 32'b00000000010000010000000100010011;
ROM[7775] <= 32'b11111111110000010000000100010011;
ROM[7776] <= 32'b00000000000000010010001110000011;
ROM[7777] <= 32'b11111111110000010000000100010011;
ROM[7778] <= 32'b00000000000000010010010000000011;
ROM[7779] <= 32'b00000000011101000010010010110011;
ROM[7780] <= 32'b00000000100000111010010100110011;
ROM[7781] <= 32'b00000000101001001000001110110011;
ROM[7782] <= 32'b00000000000100111000001110010011;
ROM[7783] <= 32'b00000000000100111111001110010011;
ROM[7784] <= 32'b00000000011100010010000000100011;
ROM[7785] <= 32'b00000000010000010000000100010011;
ROM[7786] <= 32'b00000001010000011010001110000011;
ROM[7787] <= 32'b00000000011100010010000000100011;
ROM[7788] <= 32'b00000000010000010000000100010011;
ROM[7789] <= 32'b11111111110000010000000100010011;
ROM[7790] <= 32'b00000000000000010010001110000011;
ROM[7791] <= 32'b11111111110000010000000100010011;
ROM[7792] <= 32'b00000000000000010010010000000011;
ROM[7793] <= 32'b00000000011101000111001110110011;
ROM[7794] <= 32'b00000000011100010010000000100011;
ROM[7795] <= 32'b00000000010000010000000100010011;
ROM[7796] <= 32'b00000000000000000000001110010011;
ROM[7797] <= 32'b00000000011100010010000000100011;
ROM[7798] <= 32'b00000000010000010000000100010011;
ROM[7799] <= 32'b11111111110000010000000100010011;
ROM[7800] <= 32'b00000000000000010010001110000011;
ROM[7801] <= 32'b11111111110000010000000100010011;
ROM[7802] <= 32'b00000000000000010010010000000011;
ROM[7803] <= 32'b00000000100000111010001110110011;
ROM[7804] <= 32'b00000000011100010010000000100011;
ROM[7805] <= 32'b00000000010000010000000100010011;
ROM[7806] <= 32'b11111111110000010000000100010011;
ROM[7807] <= 32'b00000000000000010010001110000011;
ROM[7808] <= 32'b01000000011100000000001110110011;
ROM[7809] <= 32'b00000000000100111000001110010011;
ROM[7810] <= 32'b00000000011100010010000000100011;
ROM[7811] <= 32'b00000000010000010000000100010011;
ROM[7812] <= 32'b11111111110000010000000100010011;
ROM[7813] <= 32'b00000000000000010010001110000011;
ROM[7814] <= 32'b00000000000000111000101001100011;
ROM[7815] <= 32'b00000000000000001101001110110111;
ROM[7816] <= 32'b01101110000000111000001110010011;
ROM[7817] <= 32'b00000000111000111000001110110011;
ROM[7818] <= 32'b00000000000000111000000011100111;
ROM[7819] <= 32'b00000000111000000000001110010011;
ROM[7820] <= 32'b00000000011100010010000000100011;
ROM[7821] <= 32'b00000000010000010000000100010011;
ROM[7822] <= 32'b00000000000000001000001110110111;
ROM[7823] <= 32'b10101000010000111000001110010011;
ROM[7824] <= 32'b00000000111000111000001110110011;
ROM[7825] <= 32'b00000000011100010010000000100011;
ROM[7826] <= 32'b00000000010000010000000100010011;
ROM[7827] <= 32'b00000000001100010010000000100011;
ROM[7828] <= 32'b00000000010000010000000100010011;
ROM[7829] <= 32'b00000000010000010010000000100011;
ROM[7830] <= 32'b00000000010000010000000100010011;
ROM[7831] <= 32'b00000000010100010010000000100011;
ROM[7832] <= 32'b00000000010000010000000100010011;
ROM[7833] <= 32'b00000000011000010010000000100011;
ROM[7834] <= 32'b00000000010000010000000100010011;
ROM[7835] <= 32'b00000001010000000000001110010011;
ROM[7836] <= 32'b00000000010000111000001110010011;
ROM[7837] <= 32'b01000000011100010000001110110011;
ROM[7838] <= 32'b00000000011100000000001000110011;
ROM[7839] <= 32'b00000000001000000000000110110011;
ROM[7840] <= 32'b01001011110100100001000011101111;
ROM[7841] <= 32'b00000100001100000000001110010011;
ROM[7842] <= 32'b00000000011100010010000000100011;
ROM[7843] <= 32'b00000000010000010000000100010011;
ROM[7844] <= 32'b00000000000000001000001110110111;
ROM[7845] <= 32'b10101101110000111000001110010011;
ROM[7846] <= 32'b00000000111000111000001110110011;
ROM[7847] <= 32'b00000000011100010010000000100011;
ROM[7848] <= 32'b00000000010000010000000100010011;
ROM[7849] <= 32'b00000000001100010010000000100011;
ROM[7850] <= 32'b00000000010000010000000100010011;
ROM[7851] <= 32'b00000000010000010010000000100011;
ROM[7852] <= 32'b00000000010000010000000100010011;
ROM[7853] <= 32'b00000000010100010010000000100011;
ROM[7854] <= 32'b00000000010000010000000100010011;
ROM[7855] <= 32'b00000000011000010010000000100011;
ROM[7856] <= 32'b00000000010000010000000100010011;
ROM[7857] <= 32'b00000001010000000000001110010011;
ROM[7858] <= 32'b00000000100000111000001110010011;
ROM[7859] <= 32'b01000000011100010000001110110011;
ROM[7860] <= 32'b00000000011100000000001000110011;
ROM[7861] <= 32'b00000000001000000000000110110011;
ROM[7862] <= 32'b00001101010000100010000011101111;
ROM[7863] <= 32'b00000111010100000000001110010011;
ROM[7864] <= 32'b00000000011100010010000000100011;
ROM[7865] <= 32'b00000000010000010000000100010011;
ROM[7866] <= 32'b00000000000000001000001110110111;
ROM[7867] <= 32'b10110011010000111000001110010011;
ROM[7868] <= 32'b00000000111000111000001110110011;
ROM[7869] <= 32'b00000000011100010010000000100011;
ROM[7870] <= 32'b00000000010000010000000100010011;
ROM[7871] <= 32'b00000000001100010010000000100011;
ROM[7872] <= 32'b00000000010000010000000100010011;
ROM[7873] <= 32'b00000000010000010010000000100011;
ROM[7874] <= 32'b00000000010000010000000100010011;
ROM[7875] <= 32'b00000000010100010010000000100011;
ROM[7876] <= 32'b00000000010000010000000100010011;
ROM[7877] <= 32'b00000000011000010010000000100011;
ROM[7878] <= 32'b00000000010000010000000100010011;
ROM[7879] <= 32'b00000001010000000000001110010011;
ROM[7880] <= 32'b00000000100000111000001110010011;
ROM[7881] <= 32'b01000000011100010000001110110011;
ROM[7882] <= 32'b00000000011100000000001000110011;
ROM[7883] <= 32'b00000000001000000000000110110011;
ROM[7884] <= 32'b00000111110000100010000011101111;
ROM[7885] <= 32'b00000111001000000000001110010011;
ROM[7886] <= 32'b00000000011100010010000000100011;
ROM[7887] <= 32'b00000000010000010000000100010011;
ROM[7888] <= 32'b00000000000000001000001110110111;
ROM[7889] <= 32'b10111000110000111000001110010011;
ROM[7890] <= 32'b00000000111000111000001110110011;
ROM[7891] <= 32'b00000000011100010010000000100011;
ROM[7892] <= 32'b00000000010000010000000100010011;
ROM[7893] <= 32'b00000000001100010010000000100011;
ROM[7894] <= 32'b00000000010000010000000100010011;
ROM[7895] <= 32'b00000000010000010010000000100011;
ROM[7896] <= 32'b00000000010000010000000100010011;
ROM[7897] <= 32'b00000000010100010010000000100011;
ROM[7898] <= 32'b00000000010000010000000100010011;
ROM[7899] <= 32'b00000000011000010010000000100011;
ROM[7900] <= 32'b00000000010000010000000100010011;
ROM[7901] <= 32'b00000001010000000000001110010011;
ROM[7902] <= 32'b00000000100000111000001110010011;
ROM[7903] <= 32'b01000000011100010000001110110011;
ROM[7904] <= 32'b00000000011100000000001000110011;
ROM[7905] <= 32'b00000000001000000000000110110011;
ROM[7906] <= 32'b00000010010000100010000011101111;
ROM[7907] <= 32'b00000111001000000000001110010011;
ROM[7908] <= 32'b00000000011100010010000000100011;
ROM[7909] <= 32'b00000000010000010000000100010011;
ROM[7910] <= 32'b00000000000000001000001110110111;
ROM[7911] <= 32'b10111110010000111000001110010011;
ROM[7912] <= 32'b00000000111000111000001110110011;
ROM[7913] <= 32'b00000000011100010010000000100011;
ROM[7914] <= 32'b00000000010000010000000100010011;
ROM[7915] <= 32'b00000000001100010010000000100011;
ROM[7916] <= 32'b00000000010000010000000100010011;
ROM[7917] <= 32'b00000000010000010010000000100011;
ROM[7918] <= 32'b00000000010000010000000100010011;
ROM[7919] <= 32'b00000000010100010010000000100011;
ROM[7920] <= 32'b00000000010000010000000100010011;
ROM[7921] <= 32'b00000000011000010010000000100011;
ROM[7922] <= 32'b00000000010000010000000100010011;
ROM[7923] <= 32'b00000001010000000000001110010011;
ROM[7924] <= 32'b00000000100000111000001110010011;
ROM[7925] <= 32'b01000000011100010000001110110011;
ROM[7926] <= 32'b00000000011100000000001000110011;
ROM[7927] <= 32'b00000000001000000000000110110011;
ROM[7928] <= 32'b01111100110100100001000011101111;
ROM[7929] <= 32'b00000110010100000000001110010011;
ROM[7930] <= 32'b00000000011100010010000000100011;
ROM[7931] <= 32'b00000000010000010000000100010011;
ROM[7932] <= 32'b00000000000000001000001110110111;
ROM[7933] <= 32'b11000011110000111000001110010011;
ROM[7934] <= 32'b00000000111000111000001110110011;
ROM[7935] <= 32'b00000000011100010010000000100011;
ROM[7936] <= 32'b00000000010000010000000100010011;
ROM[7937] <= 32'b00000000001100010010000000100011;
ROM[7938] <= 32'b00000000010000010000000100010011;
ROM[7939] <= 32'b00000000010000010010000000100011;
ROM[7940] <= 32'b00000000010000010000000100010011;
ROM[7941] <= 32'b00000000010100010010000000100011;
ROM[7942] <= 32'b00000000010000010000000100010011;
ROM[7943] <= 32'b00000000011000010010000000100011;
ROM[7944] <= 32'b00000000010000010000000100010011;
ROM[7945] <= 32'b00000001010000000000001110010011;
ROM[7946] <= 32'b00000000100000111000001110010011;
ROM[7947] <= 32'b01000000011100010000001110110011;
ROM[7948] <= 32'b00000000011100000000001000110011;
ROM[7949] <= 32'b00000000001000000000000110110011;
ROM[7950] <= 32'b01110111010100100001000011101111;
ROM[7951] <= 32'b00000110111000000000001110010011;
ROM[7952] <= 32'b00000000011100010010000000100011;
ROM[7953] <= 32'b00000000010000010000000100010011;
ROM[7954] <= 32'b00000000000000001000001110110111;
ROM[7955] <= 32'b11001001010000111000001110010011;
ROM[7956] <= 32'b00000000111000111000001110110011;
ROM[7957] <= 32'b00000000011100010010000000100011;
ROM[7958] <= 32'b00000000010000010000000100010011;
ROM[7959] <= 32'b00000000001100010010000000100011;
ROM[7960] <= 32'b00000000010000010000000100010011;
ROM[7961] <= 32'b00000000010000010010000000100011;
ROM[7962] <= 32'b00000000010000010000000100010011;
ROM[7963] <= 32'b00000000010100010010000000100011;
ROM[7964] <= 32'b00000000010000010000000100010011;
ROM[7965] <= 32'b00000000011000010010000000100011;
ROM[7966] <= 32'b00000000010000010000000100010011;
ROM[7967] <= 32'b00000001010000000000001110010011;
ROM[7968] <= 32'b00000000100000111000001110010011;
ROM[7969] <= 32'b01000000011100010000001110110011;
ROM[7970] <= 32'b00000000011100000000001000110011;
ROM[7971] <= 32'b00000000001000000000000110110011;
ROM[7972] <= 32'b01110001110100100001000011101111;
ROM[7973] <= 32'b00000111010000000000001110010011;
ROM[7974] <= 32'b00000000011100010010000000100011;
ROM[7975] <= 32'b00000000010000010000000100010011;
ROM[7976] <= 32'b00000000000000001000001110110111;
ROM[7977] <= 32'b11001110110000111000001110010011;
ROM[7978] <= 32'b00000000111000111000001110110011;
ROM[7979] <= 32'b00000000011100010010000000100011;
ROM[7980] <= 32'b00000000010000010000000100010011;
ROM[7981] <= 32'b00000000001100010010000000100011;
ROM[7982] <= 32'b00000000010000010000000100010011;
ROM[7983] <= 32'b00000000010000010010000000100011;
ROM[7984] <= 32'b00000000010000010000000100010011;
ROM[7985] <= 32'b00000000010100010010000000100011;
ROM[7986] <= 32'b00000000010000010000000100010011;
ROM[7987] <= 32'b00000000011000010010000000100011;
ROM[7988] <= 32'b00000000010000010000000100010011;
ROM[7989] <= 32'b00000001010000000000001110010011;
ROM[7990] <= 32'b00000000100000111000001110010011;
ROM[7991] <= 32'b01000000011100010000001110110011;
ROM[7992] <= 32'b00000000011100000000001000110011;
ROM[7993] <= 32'b00000000001000000000000110110011;
ROM[7994] <= 32'b01101100010100100001000011101111;
ROM[7995] <= 32'b00000010000000000000001110010011;
ROM[7996] <= 32'b00000000011100010010000000100011;
ROM[7997] <= 32'b00000000010000010000000100010011;
ROM[7998] <= 32'b00000000000000001000001110110111;
ROM[7999] <= 32'b11010100010000111000001110010011;
ROM[8000] <= 32'b00000000111000111000001110110011;
ROM[8001] <= 32'b00000000011100010010000000100011;
ROM[8002] <= 32'b00000000010000010000000100010011;
ROM[8003] <= 32'b00000000001100010010000000100011;
ROM[8004] <= 32'b00000000010000010000000100010011;
ROM[8005] <= 32'b00000000010000010010000000100011;
ROM[8006] <= 32'b00000000010000010000000100010011;
ROM[8007] <= 32'b00000000010100010010000000100011;
ROM[8008] <= 32'b00000000010000010000000100010011;
ROM[8009] <= 32'b00000000011000010010000000100011;
ROM[8010] <= 32'b00000000010000010000000100010011;
ROM[8011] <= 32'b00000001010000000000001110010011;
ROM[8012] <= 32'b00000000100000111000001110010011;
ROM[8013] <= 32'b01000000011100010000001110110011;
ROM[8014] <= 32'b00000000011100000000001000110011;
ROM[8015] <= 32'b00000000001000000000000110110011;
ROM[8016] <= 32'b01100110110100100001000011101111;
ROM[8017] <= 32'b00000111011100000000001110010011;
ROM[8018] <= 32'b00000000011100010010000000100011;
ROM[8019] <= 32'b00000000010000010000000100010011;
ROM[8020] <= 32'b00000000000000001000001110110111;
ROM[8021] <= 32'b11011001110000111000001110010011;
ROM[8022] <= 32'b00000000111000111000001110110011;
ROM[8023] <= 32'b00000000011100010010000000100011;
ROM[8024] <= 32'b00000000010000010000000100010011;
ROM[8025] <= 32'b00000000001100010010000000100011;
ROM[8026] <= 32'b00000000010000010000000100010011;
ROM[8027] <= 32'b00000000010000010010000000100011;
ROM[8028] <= 32'b00000000010000010000000100010011;
ROM[8029] <= 32'b00000000010100010010000000100011;
ROM[8030] <= 32'b00000000010000010000000100010011;
ROM[8031] <= 32'b00000000011000010010000000100011;
ROM[8032] <= 32'b00000000010000010000000100010011;
ROM[8033] <= 32'b00000001010000000000001110010011;
ROM[8034] <= 32'b00000000100000111000001110010011;
ROM[8035] <= 32'b01000000011100010000001110110011;
ROM[8036] <= 32'b00000000011100000000001000110011;
ROM[8037] <= 32'b00000000001000000000000110110011;
ROM[8038] <= 32'b01100001010100100001000011101111;
ROM[8039] <= 32'b00000110111100000000001110010011;
ROM[8040] <= 32'b00000000011100010010000000100011;
ROM[8041] <= 32'b00000000010000010000000100010011;
ROM[8042] <= 32'b00000000000000001000001110110111;
ROM[8043] <= 32'b11011111010000111000001110010011;
ROM[8044] <= 32'b00000000111000111000001110110011;
ROM[8045] <= 32'b00000000011100010010000000100011;
ROM[8046] <= 32'b00000000010000010000000100010011;
ROM[8047] <= 32'b00000000001100010010000000100011;
ROM[8048] <= 32'b00000000010000010000000100010011;
ROM[8049] <= 32'b00000000010000010010000000100011;
ROM[8050] <= 32'b00000000010000010000000100010011;
ROM[8051] <= 32'b00000000010100010010000000100011;
ROM[8052] <= 32'b00000000010000010000000100010011;
ROM[8053] <= 32'b00000000011000010010000000100011;
ROM[8054] <= 32'b00000000010000010000000100010011;
ROM[8055] <= 32'b00000001010000000000001110010011;
ROM[8056] <= 32'b00000000100000111000001110010011;
ROM[8057] <= 32'b01000000011100010000001110110011;
ROM[8058] <= 32'b00000000011100000000001000110011;
ROM[8059] <= 32'b00000000001000000000000110110011;
ROM[8060] <= 32'b01011011110100100001000011101111;
ROM[8061] <= 32'b00000111001000000000001110010011;
ROM[8062] <= 32'b00000000011100010010000000100011;
ROM[8063] <= 32'b00000000010000010000000100010011;
ROM[8064] <= 32'b00000000000000001000001110110111;
ROM[8065] <= 32'b11100100110000111000001110010011;
ROM[8066] <= 32'b00000000111000111000001110110011;
ROM[8067] <= 32'b00000000011100010010000000100011;
ROM[8068] <= 32'b00000000010000010000000100010011;
ROM[8069] <= 32'b00000000001100010010000000100011;
ROM[8070] <= 32'b00000000010000010000000100010011;
ROM[8071] <= 32'b00000000010000010010000000100011;
ROM[8072] <= 32'b00000000010000010000000100010011;
ROM[8073] <= 32'b00000000010100010010000000100011;
ROM[8074] <= 32'b00000000010000010000000100010011;
ROM[8075] <= 32'b00000000011000010010000000100011;
ROM[8076] <= 32'b00000000010000010000000100010011;
ROM[8077] <= 32'b00000001010000000000001110010011;
ROM[8078] <= 32'b00000000100000111000001110010011;
ROM[8079] <= 32'b01000000011100010000001110110011;
ROM[8080] <= 32'b00000000011100000000001000110011;
ROM[8081] <= 32'b00000000001000000000000110110011;
ROM[8082] <= 32'b01010110010100100001000011101111;
ROM[8083] <= 32'b00000110010000000000001110010011;
ROM[8084] <= 32'b00000000011100010010000000100011;
ROM[8085] <= 32'b00000000010000010000000100010011;
ROM[8086] <= 32'b00000000000000001000001110110111;
ROM[8087] <= 32'b11101010010000111000001110010011;
ROM[8088] <= 32'b00000000111000111000001110110011;
ROM[8089] <= 32'b00000000011100010010000000100011;
ROM[8090] <= 32'b00000000010000010000000100010011;
ROM[8091] <= 32'b00000000001100010010000000100011;
ROM[8092] <= 32'b00000000010000010000000100010011;
ROM[8093] <= 32'b00000000010000010010000000100011;
ROM[8094] <= 32'b00000000010000010000000100010011;
ROM[8095] <= 32'b00000000010100010010000000100011;
ROM[8096] <= 32'b00000000010000010000000100010011;
ROM[8097] <= 32'b00000000011000010010000000100011;
ROM[8098] <= 32'b00000000010000010000000100010011;
ROM[8099] <= 32'b00000001010000000000001110010011;
ROM[8100] <= 32'b00000000100000111000001110010011;
ROM[8101] <= 32'b01000000011100010000001110110011;
ROM[8102] <= 32'b00000000011100000000001000110011;
ROM[8103] <= 32'b00000000001000000000000110110011;
ROM[8104] <= 32'b01010000110100100001000011101111;
ROM[8105] <= 32'b00000011101000000000001110010011;
ROM[8106] <= 32'b00000000011100010010000000100011;
ROM[8107] <= 32'b00000000010000010000000100010011;
ROM[8108] <= 32'b00000000000000001000001110110111;
ROM[8109] <= 32'b11101111110000111000001110010011;
ROM[8110] <= 32'b00000000111000111000001110110011;
ROM[8111] <= 32'b00000000011100010010000000100011;
ROM[8112] <= 32'b00000000010000010000000100010011;
ROM[8113] <= 32'b00000000001100010010000000100011;
ROM[8114] <= 32'b00000000010000010000000100010011;
ROM[8115] <= 32'b00000000010000010010000000100011;
ROM[8116] <= 32'b00000000010000010000000100010011;
ROM[8117] <= 32'b00000000010100010010000000100011;
ROM[8118] <= 32'b00000000010000010000000100010011;
ROM[8119] <= 32'b00000000011000010010000000100011;
ROM[8120] <= 32'b00000000010000010000000100010011;
ROM[8121] <= 32'b00000001010000000000001110010011;
ROM[8122] <= 32'b00000000100000111000001110010011;
ROM[8123] <= 32'b01000000011100010000001110110011;
ROM[8124] <= 32'b00000000011100000000001000110011;
ROM[8125] <= 32'b00000000001000000000000110110011;
ROM[8126] <= 32'b01001011010100100001000011101111;
ROM[8127] <= 32'b00000010000000000000001110010011;
ROM[8128] <= 32'b00000000011100010010000000100011;
ROM[8129] <= 32'b00000000010000010000000100010011;
ROM[8130] <= 32'b00000000000000001000001110110111;
ROM[8131] <= 32'b11110101010000111000001110010011;
ROM[8132] <= 32'b00000000111000111000001110110011;
ROM[8133] <= 32'b00000000011100010010000000100011;
ROM[8134] <= 32'b00000000010000010000000100010011;
ROM[8135] <= 32'b00000000001100010010000000100011;
ROM[8136] <= 32'b00000000010000010000000100010011;
ROM[8137] <= 32'b00000000010000010010000000100011;
ROM[8138] <= 32'b00000000010000010000000100010011;
ROM[8139] <= 32'b00000000010100010010000000100011;
ROM[8140] <= 32'b00000000010000010000000100010011;
ROM[8141] <= 32'b00000000011000010010000000100011;
ROM[8142] <= 32'b00000000010000010000000100010011;
ROM[8143] <= 32'b00000001010000000000001110010011;
ROM[8144] <= 32'b00000000100000111000001110010011;
ROM[8145] <= 32'b01000000011100010000001110110011;
ROM[8146] <= 32'b00000000011100000000001000110011;
ROM[8147] <= 32'b00000000001000000000000110110011;
ROM[8148] <= 32'b01000101110100100001000011101111;
ROM[8149] <= 32'b00000000000000001000001110110111;
ROM[8150] <= 32'b11111010000000111000001110010011;
ROM[8151] <= 32'b00000000111000111000001110110011;
ROM[8152] <= 32'b00000000011100010010000000100011;
ROM[8153] <= 32'b00000000010000010000000100010011;
ROM[8154] <= 32'b00000000001100010010000000100011;
ROM[8155] <= 32'b00000000010000010000000100010011;
ROM[8156] <= 32'b00000000010000010010000000100011;
ROM[8157] <= 32'b00000000010000010000000100010011;
ROM[8158] <= 32'b00000000010100010010000000100011;
ROM[8159] <= 32'b00000000010000010000000100010011;
ROM[8160] <= 32'b00000000011000010010000000100011;
ROM[8161] <= 32'b00000000010000010000000100010011;
ROM[8162] <= 32'b00000001010000000000001110010011;
ROM[8163] <= 32'b00000000010000111000001110010011;
ROM[8164] <= 32'b01000000011100010000001110110011;
ROM[8165] <= 32'b00000000011100000000001000110011;
ROM[8166] <= 32'b00000000001000000000000110110011;
ROM[8167] <= 32'b01111100110100001110000011101111;
ROM[8168] <= 32'b11111111110000010000000100010011;
ROM[8169] <= 32'b00000000000000010010001110000011;
ROM[8170] <= 32'b00000000011101100010000000100011;
ROM[8171] <= 32'b00000001100000011010001110000011;
ROM[8172] <= 32'b00000000011100010010000000100011;
ROM[8173] <= 32'b00000000010000010000000100010011;
ROM[8174] <= 32'b00000000000000001000001110110111;
ROM[8175] <= 32'b00000000010000111000001110010011;
ROM[8176] <= 32'b00000000111000111000001110110011;
ROM[8177] <= 32'b00000000011100010010000000100011;
ROM[8178] <= 32'b00000000010000010000000100010011;
ROM[8179] <= 32'b00000000001100010010000000100011;
ROM[8180] <= 32'b00000000010000010000000100010011;
ROM[8181] <= 32'b00000000010000010010000000100011;
ROM[8182] <= 32'b00000000010000010000000100010011;
ROM[8183] <= 32'b00000000010100010010000000100011;
ROM[8184] <= 32'b00000000010000010000000100010011;
ROM[8185] <= 32'b00000000011000010010000000100011;
ROM[8186] <= 32'b00000000010000010000000100010011;
ROM[8187] <= 32'b00000001010000000000001110010011;
ROM[8188] <= 32'b00000000010000111000001110010011;
ROM[8189] <= 32'b01000000011100010000001110110011;
ROM[8190] <= 32'b00000000011100000000001000110011;
ROM[8191] <= 32'b00000000001000000000000110110011;
ROM[8192] <= 32'b01110110100100001110000011101111;
ROM[8193] <= 32'b11111111110000010000000100010011;
ROM[8194] <= 32'b00000000000000010010001110000011;
ROM[8195] <= 32'b00000000011101100010000000100011;
ROM[8196] <= 32'b00000000000000001000001110110111;
ROM[8197] <= 32'b00000101110000111000001110010011;
ROM[8198] <= 32'b00000000111000111000001110110011;
ROM[8199] <= 32'b00000000011100010010000000100011;
ROM[8200] <= 32'b00000000010000010000000100010011;
ROM[8201] <= 32'b00000000001100010010000000100011;
ROM[8202] <= 32'b00000000010000010000000100010011;
ROM[8203] <= 32'b00000000010000010010000000100011;
ROM[8204] <= 32'b00000000010000010000000100010011;
ROM[8205] <= 32'b00000000010100010010000000100011;
ROM[8206] <= 32'b00000000010000010000000100010011;
ROM[8207] <= 32'b00000000011000010010000000100011;
ROM[8208] <= 32'b00000000010000010000000100010011;
ROM[8209] <= 32'b00000001010000000000001110010011;
ROM[8210] <= 32'b00000000000000111000001110010011;
ROM[8211] <= 32'b01000000011100010000001110110011;
ROM[8212] <= 32'b00000000011100000000001000110011;
ROM[8213] <= 32'b00000000001000000000000110110011;
ROM[8214] <= 32'b00110001000000001111000011101111;
ROM[8215] <= 32'b11111111110000010000000100010011;
ROM[8216] <= 32'b00000000000000010010001110000011;
ROM[8217] <= 32'b00000000011101100010000000100011;
ROM[8218] <= 32'b00000001101000000000001110010011;
ROM[8219] <= 32'b00000000011100010010000000100011;
ROM[8220] <= 32'b00000000010000010000000100010011;
ROM[8221] <= 32'b00000000000000001000001110110111;
ROM[8222] <= 32'b00001100000000111000001110010011;
ROM[8223] <= 32'b00000000111000111000001110110011;
ROM[8224] <= 32'b00000000011100010010000000100011;
ROM[8225] <= 32'b00000000010000010000000100010011;
ROM[8226] <= 32'b00000000001100010010000000100011;
ROM[8227] <= 32'b00000000010000010000000100010011;
ROM[8228] <= 32'b00000000010000010010000000100011;
ROM[8229] <= 32'b00000000010000010000000100010011;
ROM[8230] <= 32'b00000000010100010010000000100011;
ROM[8231] <= 32'b00000000010000010000000100010011;
ROM[8232] <= 32'b00000000011000010010000000100011;
ROM[8233] <= 32'b00000000010000010000000100010011;
ROM[8234] <= 32'b00000001010000000000001110010011;
ROM[8235] <= 32'b00000000010000111000001110010011;
ROM[8236] <= 32'b01000000011100010000001110110011;
ROM[8237] <= 32'b00000000011100000000001000110011;
ROM[8238] <= 32'b00000000001000000000000110110011;
ROM[8239] <= 32'b01101000000000100001000011101111;
ROM[8240] <= 32'b00000100010100000000001110010011;
ROM[8241] <= 32'b00000000011100010010000000100011;
ROM[8242] <= 32'b00000000010000010000000100010011;
ROM[8243] <= 32'b00000000000000001000001110110111;
ROM[8244] <= 32'b00010001100000111000001110010011;
ROM[8245] <= 32'b00000000111000111000001110110011;
ROM[8246] <= 32'b00000000011100010010000000100011;
ROM[8247] <= 32'b00000000010000010000000100010011;
ROM[8248] <= 32'b00000000001100010010000000100011;
ROM[8249] <= 32'b00000000010000010000000100010011;
ROM[8250] <= 32'b00000000010000010010000000100011;
ROM[8251] <= 32'b00000000010000010000000100010011;
ROM[8252] <= 32'b00000000010100010010000000100011;
ROM[8253] <= 32'b00000000010000010000000100010011;
ROM[8254] <= 32'b00000000011000010010000000100011;
ROM[8255] <= 32'b00000000010000010000000100010011;
ROM[8256] <= 32'b00000001010000000000001110010011;
ROM[8257] <= 32'b00000000100000111000001110010011;
ROM[8258] <= 32'b01000000011100010000001110110011;
ROM[8259] <= 32'b00000000011100000000001000110011;
ROM[8260] <= 32'b00000000001000000000000110110011;
ROM[8261] <= 32'b00101001100100100001000011101111;
ROM[8262] <= 32'b00000110111000000000001110010011;
ROM[8263] <= 32'b00000000011100010010000000100011;
ROM[8264] <= 32'b00000000010000010000000100010011;
ROM[8265] <= 32'b00000000000000001000001110110111;
ROM[8266] <= 32'b00010111000000111000001110010011;
ROM[8267] <= 32'b00000000111000111000001110110011;
ROM[8268] <= 32'b00000000011100010010000000100011;
ROM[8269] <= 32'b00000000010000010000000100010011;
ROM[8270] <= 32'b00000000001100010010000000100011;
ROM[8271] <= 32'b00000000010000010000000100010011;
ROM[8272] <= 32'b00000000010000010010000000100011;
ROM[8273] <= 32'b00000000010000010000000100010011;
ROM[8274] <= 32'b00000000010100010010000000100011;
ROM[8275] <= 32'b00000000010000010000000100010011;
ROM[8276] <= 32'b00000000011000010010000000100011;
ROM[8277] <= 32'b00000000010000010000000100010011;
ROM[8278] <= 32'b00000001010000000000001110010011;
ROM[8279] <= 32'b00000000100000111000001110010011;
ROM[8280] <= 32'b01000000011100010000001110110011;
ROM[8281] <= 32'b00000000011100000000001000110011;
ROM[8282] <= 32'b00000000001000000000000110110011;
ROM[8283] <= 32'b00100100000100100001000011101111;
ROM[8284] <= 32'b00000111010000000000001110010011;
ROM[8285] <= 32'b00000000011100010010000000100011;
ROM[8286] <= 32'b00000000010000010000000100010011;
ROM[8287] <= 32'b00000000000000001000001110110111;
ROM[8288] <= 32'b00011100100000111000001110010011;
ROM[8289] <= 32'b00000000111000111000001110110011;
ROM[8290] <= 32'b00000000011100010010000000100011;
ROM[8291] <= 32'b00000000010000010000000100010011;
ROM[8292] <= 32'b00000000001100010010000000100011;
ROM[8293] <= 32'b00000000010000010000000100010011;
ROM[8294] <= 32'b00000000010000010010000000100011;
ROM[8295] <= 32'b00000000010000010000000100010011;
ROM[8296] <= 32'b00000000010100010010000000100011;
ROM[8297] <= 32'b00000000010000010000000100010011;
ROM[8298] <= 32'b00000000011000010010000000100011;
ROM[8299] <= 32'b00000000010000010000000100010011;
ROM[8300] <= 32'b00000001010000000000001110010011;
ROM[8301] <= 32'b00000000100000111000001110010011;
ROM[8302] <= 32'b01000000011100010000001110110011;
ROM[8303] <= 32'b00000000011100000000001000110011;
ROM[8304] <= 32'b00000000001000000000000110110011;
ROM[8305] <= 32'b00011110100100100001000011101111;
ROM[8306] <= 32'b00000110010100000000001110010011;
ROM[8307] <= 32'b00000000011100010010000000100011;
ROM[8308] <= 32'b00000000010000010000000100010011;
ROM[8309] <= 32'b00000000000000001000001110110111;
ROM[8310] <= 32'b00100010000000111000001110010011;
ROM[8311] <= 32'b00000000111000111000001110110011;
ROM[8312] <= 32'b00000000011100010010000000100011;
ROM[8313] <= 32'b00000000010000010000000100010011;
ROM[8314] <= 32'b00000000001100010010000000100011;
ROM[8315] <= 32'b00000000010000010000000100010011;
ROM[8316] <= 32'b00000000010000010010000000100011;
ROM[8317] <= 32'b00000000010000010000000100010011;
ROM[8318] <= 32'b00000000010100010010000000100011;
ROM[8319] <= 32'b00000000010000010000000100010011;
ROM[8320] <= 32'b00000000011000010010000000100011;
ROM[8321] <= 32'b00000000010000010000000100010011;
ROM[8322] <= 32'b00000001010000000000001110010011;
ROM[8323] <= 32'b00000000100000111000001110010011;
ROM[8324] <= 32'b01000000011100010000001110110011;
ROM[8325] <= 32'b00000000011100000000001000110011;
ROM[8326] <= 32'b00000000001000000000000110110011;
ROM[8327] <= 32'b00011001000100100001000011101111;
ROM[8328] <= 32'b00000111001000000000001110010011;
ROM[8329] <= 32'b00000000011100010010000000100011;
ROM[8330] <= 32'b00000000010000010000000100010011;
ROM[8331] <= 32'b00000000000000001000001110110111;
ROM[8332] <= 32'b00100111100000111000001110010011;
ROM[8333] <= 32'b00000000111000111000001110110011;
ROM[8334] <= 32'b00000000011100010010000000100011;
ROM[8335] <= 32'b00000000010000010000000100010011;
ROM[8336] <= 32'b00000000001100010010000000100011;
ROM[8337] <= 32'b00000000010000010000000100010011;
ROM[8338] <= 32'b00000000010000010010000000100011;
ROM[8339] <= 32'b00000000010000010000000100010011;
ROM[8340] <= 32'b00000000010100010010000000100011;
ROM[8341] <= 32'b00000000010000010000000100010011;
ROM[8342] <= 32'b00000000011000010010000000100011;
ROM[8343] <= 32'b00000000010000010000000100010011;
ROM[8344] <= 32'b00000001010000000000001110010011;
ROM[8345] <= 32'b00000000100000111000001110010011;
ROM[8346] <= 32'b01000000011100010000001110110011;
ROM[8347] <= 32'b00000000011100000000001000110011;
ROM[8348] <= 32'b00000000001000000000000110110011;
ROM[8349] <= 32'b00010011100100100001000011101111;
ROM[8350] <= 32'b00000010000000000000001110010011;
ROM[8351] <= 32'b00000000011100010010000000100011;
ROM[8352] <= 32'b00000000010000010000000100010011;
ROM[8353] <= 32'b00000000000000001000001110110111;
ROM[8354] <= 32'b00101101000000111000001110010011;
ROM[8355] <= 32'b00000000111000111000001110110011;
ROM[8356] <= 32'b00000000011100010010000000100011;
ROM[8357] <= 32'b00000000010000010000000100010011;
ROM[8358] <= 32'b00000000001100010010000000100011;
ROM[8359] <= 32'b00000000010000010000000100010011;
ROM[8360] <= 32'b00000000010000010010000000100011;
ROM[8361] <= 32'b00000000010000010000000100010011;
ROM[8362] <= 32'b00000000010100010010000000100011;
ROM[8363] <= 32'b00000000010000010000000100010011;
ROM[8364] <= 32'b00000000011000010010000000100011;
ROM[8365] <= 32'b00000000010000010000000100010011;
ROM[8366] <= 32'b00000001010000000000001110010011;
ROM[8367] <= 32'b00000000100000111000001110010011;
ROM[8368] <= 32'b01000000011100010000001110110011;
ROM[8369] <= 32'b00000000011100000000001000110011;
ROM[8370] <= 32'b00000000001000000000000110110011;
ROM[8371] <= 32'b00001110000100100001000011101111;
ROM[8372] <= 32'b00000110000100000000001110010011;
ROM[8373] <= 32'b00000000011100010010000000100011;
ROM[8374] <= 32'b00000000010000010000000100010011;
ROM[8375] <= 32'b00000000000000001000001110110111;
ROM[8376] <= 32'b00110010100000111000001110010011;
ROM[8377] <= 32'b00000000111000111000001110110011;
ROM[8378] <= 32'b00000000011100010010000000100011;
ROM[8379] <= 32'b00000000010000010000000100010011;
ROM[8380] <= 32'b00000000001100010010000000100011;
ROM[8381] <= 32'b00000000010000010000000100010011;
ROM[8382] <= 32'b00000000010000010010000000100011;
ROM[8383] <= 32'b00000000010000010000000100010011;
ROM[8384] <= 32'b00000000010100010010000000100011;
ROM[8385] <= 32'b00000000010000010000000100010011;
ROM[8386] <= 32'b00000000011000010010000000100011;
ROM[8387] <= 32'b00000000010000010000000100010011;
ROM[8388] <= 32'b00000001010000000000001110010011;
ROM[8389] <= 32'b00000000100000111000001110010011;
ROM[8390] <= 32'b01000000011100010000001110110011;
ROM[8391] <= 32'b00000000011100000000001000110011;
ROM[8392] <= 32'b00000000001000000000000110110011;
ROM[8393] <= 32'b00001000100100100001000011101111;
ROM[8394] <= 32'b00000010000000000000001110010011;
ROM[8395] <= 32'b00000000011100010010000000100011;
ROM[8396] <= 32'b00000000010000010000000100010011;
ROM[8397] <= 32'b00000000000000001000001110110111;
ROM[8398] <= 32'b00111000000000111000001110010011;
ROM[8399] <= 32'b00000000111000111000001110110011;
ROM[8400] <= 32'b00000000011100010010000000100011;
ROM[8401] <= 32'b00000000010000010000000100010011;
ROM[8402] <= 32'b00000000001100010010000000100011;
ROM[8403] <= 32'b00000000010000010000000100010011;
ROM[8404] <= 32'b00000000010000010010000000100011;
ROM[8405] <= 32'b00000000010000010000000100010011;
ROM[8406] <= 32'b00000000010100010010000000100011;
ROM[8407] <= 32'b00000000010000010000000100010011;
ROM[8408] <= 32'b00000000011000010010000000100011;
ROM[8409] <= 32'b00000000010000010000000100010011;
ROM[8410] <= 32'b00000001010000000000001110010011;
ROM[8411] <= 32'b00000000100000111000001110010011;
ROM[8412] <= 32'b01000000011100010000001110110011;
ROM[8413] <= 32'b00000000011100000000001000110011;
ROM[8414] <= 32'b00000000001000000000000110110011;
ROM[8415] <= 32'b00000011000100100001000011101111;
ROM[8416] <= 32'b00000110110000000000001110010011;
ROM[8417] <= 32'b00000000011100010010000000100011;
ROM[8418] <= 32'b00000000010000010000000100010011;
ROM[8419] <= 32'b00000000000000001000001110110111;
ROM[8420] <= 32'b00111101100000111000001110010011;
ROM[8421] <= 32'b00000000111000111000001110110011;
ROM[8422] <= 32'b00000000011100010010000000100011;
ROM[8423] <= 32'b00000000010000010000000100010011;
ROM[8424] <= 32'b00000000001100010010000000100011;
ROM[8425] <= 32'b00000000010000010000000100010011;
ROM[8426] <= 32'b00000000010000010010000000100011;
ROM[8427] <= 32'b00000000010000010000000100010011;
ROM[8428] <= 32'b00000000010100010010000000100011;
ROM[8429] <= 32'b00000000010000010000000100010011;
ROM[8430] <= 32'b00000000011000010010000000100011;
ROM[8431] <= 32'b00000000010000010000000100010011;
ROM[8432] <= 32'b00000001010000000000001110010011;
ROM[8433] <= 32'b00000000100000111000001110010011;
ROM[8434] <= 32'b01000000011100010000001110110011;
ROM[8435] <= 32'b00000000011100000000001000110011;
ROM[8436] <= 32'b00000000001000000000000110110011;
ROM[8437] <= 32'b01111101100000100001000011101111;
ROM[8438] <= 32'b00000110010100000000001110010011;
ROM[8439] <= 32'b00000000011100010010000000100011;
ROM[8440] <= 32'b00000000010000010000000100010011;
ROM[8441] <= 32'b00000000000000001000001110110111;
ROM[8442] <= 32'b01000011000000111000001110010011;
ROM[8443] <= 32'b00000000111000111000001110110011;
ROM[8444] <= 32'b00000000011100010010000000100011;
ROM[8445] <= 32'b00000000010000010000000100010011;
ROM[8446] <= 32'b00000000001100010010000000100011;
ROM[8447] <= 32'b00000000010000010000000100010011;
ROM[8448] <= 32'b00000000010000010010000000100011;
ROM[8449] <= 32'b00000000010000010000000100010011;
ROM[8450] <= 32'b00000000010100010010000000100011;
ROM[8451] <= 32'b00000000010000010000000100010011;
ROM[8452] <= 32'b00000000011000010010000000100011;
ROM[8453] <= 32'b00000000010000010000000100010011;
ROM[8454] <= 32'b00000001010000000000001110010011;
ROM[8455] <= 32'b00000000100000111000001110010011;
ROM[8456] <= 32'b01000000011100010000001110110011;
ROM[8457] <= 32'b00000000011100000000001000110011;
ROM[8458] <= 32'b00000000001000000000000110110011;
ROM[8459] <= 32'b01111000000000100001000011101111;
ROM[8460] <= 32'b00000111010000000000001110010011;
ROM[8461] <= 32'b00000000011100010010000000100011;
ROM[8462] <= 32'b00000000010000010000000100010011;
ROM[8463] <= 32'b00000000000000001000001110110111;
ROM[8464] <= 32'b01001000100000111000001110010011;
ROM[8465] <= 32'b00000000111000111000001110110011;
ROM[8466] <= 32'b00000000011100010010000000100011;
ROM[8467] <= 32'b00000000010000010000000100010011;
ROM[8468] <= 32'b00000000001100010010000000100011;
ROM[8469] <= 32'b00000000010000010000000100010011;
ROM[8470] <= 32'b00000000010000010010000000100011;
ROM[8471] <= 32'b00000000010000010000000100010011;
ROM[8472] <= 32'b00000000010100010010000000100011;
ROM[8473] <= 32'b00000000010000010000000100010011;
ROM[8474] <= 32'b00000000011000010010000000100011;
ROM[8475] <= 32'b00000000010000010000000100010011;
ROM[8476] <= 32'b00000001010000000000001110010011;
ROM[8477] <= 32'b00000000100000111000001110010011;
ROM[8478] <= 32'b01000000011100010000001110110011;
ROM[8479] <= 32'b00000000011100000000001000110011;
ROM[8480] <= 32'b00000000001000000000000110110011;
ROM[8481] <= 32'b01110010100000100001000011101111;
ROM[8482] <= 32'b00000111010000000000001110010011;
ROM[8483] <= 32'b00000000011100010010000000100011;
ROM[8484] <= 32'b00000000010000010000000100010011;
ROM[8485] <= 32'b00000000000000001000001110110111;
ROM[8486] <= 32'b01001110000000111000001110010011;
ROM[8487] <= 32'b00000000111000111000001110110011;
ROM[8488] <= 32'b00000000011100010010000000100011;
ROM[8489] <= 32'b00000000010000010000000100010011;
ROM[8490] <= 32'b00000000001100010010000000100011;
ROM[8491] <= 32'b00000000010000010000000100010011;
ROM[8492] <= 32'b00000000010000010010000000100011;
ROM[8493] <= 32'b00000000010000010000000100010011;
ROM[8494] <= 32'b00000000010100010010000000100011;
ROM[8495] <= 32'b00000000010000010000000100010011;
ROM[8496] <= 32'b00000000011000010010000000100011;
ROM[8497] <= 32'b00000000010000010000000100010011;
ROM[8498] <= 32'b00000001010000000000001110010011;
ROM[8499] <= 32'b00000000100000111000001110010011;
ROM[8500] <= 32'b01000000011100010000001110110011;
ROM[8501] <= 32'b00000000011100000000001000110011;
ROM[8502] <= 32'b00000000001000000000000110110011;
ROM[8503] <= 32'b01101101000000100001000011101111;
ROM[8504] <= 32'b00000110010100000000001110010011;
ROM[8505] <= 32'b00000000011100010010000000100011;
ROM[8506] <= 32'b00000000010000010000000100010011;
ROM[8507] <= 32'b00000000000000001000001110110111;
ROM[8508] <= 32'b01010011100000111000001110010011;
ROM[8509] <= 32'b00000000111000111000001110110011;
ROM[8510] <= 32'b00000000011100010010000000100011;
ROM[8511] <= 32'b00000000010000010000000100010011;
ROM[8512] <= 32'b00000000001100010010000000100011;
ROM[8513] <= 32'b00000000010000010000000100010011;
ROM[8514] <= 32'b00000000010000010010000000100011;
ROM[8515] <= 32'b00000000010000010000000100010011;
ROM[8516] <= 32'b00000000010100010010000000100011;
ROM[8517] <= 32'b00000000010000010000000100010011;
ROM[8518] <= 32'b00000000011000010010000000100011;
ROM[8519] <= 32'b00000000010000010000000100010011;
ROM[8520] <= 32'b00000001010000000000001110010011;
ROM[8521] <= 32'b00000000100000111000001110010011;
ROM[8522] <= 32'b01000000011100010000001110110011;
ROM[8523] <= 32'b00000000011100000000001000110011;
ROM[8524] <= 32'b00000000001000000000000110110011;
ROM[8525] <= 32'b01100111100000100001000011101111;
ROM[8526] <= 32'b00000111001000000000001110010011;
ROM[8527] <= 32'b00000000011100010010000000100011;
ROM[8528] <= 32'b00000000010000010000000100010011;
ROM[8529] <= 32'b00000000000000001000001110110111;
ROM[8530] <= 32'b01011001000000111000001110010011;
ROM[8531] <= 32'b00000000111000111000001110110011;
ROM[8532] <= 32'b00000000011100010010000000100011;
ROM[8533] <= 32'b00000000010000010000000100010011;
ROM[8534] <= 32'b00000000001100010010000000100011;
ROM[8535] <= 32'b00000000010000010000000100010011;
ROM[8536] <= 32'b00000000010000010010000000100011;
ROM[8537] <= 32'b00000000010000010000000100010011;
ROM[8538] <= 32'b00000000010100010010000000100011;
ROM[8539] <= 32'b00000000010000010000000100010011;
ROM[8540] <= 32'b00000000011000010010000000100011;
ROM[8541] <= 32'b00000000010000010000000100010011;
ROM[8542] <= 32'b00000001010000000000001110010011;
ROM[8543] <= 32'b00000000100000111000001110010011;
ROM[8544] <= 32'b01000000011100010000001110110011;
ROM[8545] <= 32'b00000000011100000000001000110011;
ROM[8546] <= 32'b00000000001000000000000110110011;
ROM[8547] <= 32'b01100010000000100001000011101111;
ROM[8548] <= 32'b00000010100000000000001110010011;
ROM[8549] <= 32'b00000000011100010010000000100011;
ROM[8550] <= 32'b00000000010000010000000100010011;
ROM[8551] <= 32'b00000000000000001000001110110111;
ROM[8552] <= 32'b01011110100000111000001110010011;
ROM[8553] <= 32'b00000000111000111000001110110011;
ROM[8554] <= 32'b00000000011100010010000000100011;
ROM[8555] <= 32'b00000000010000010000000100010011;
ROM[8556] <= 32'b00000000001100010010000000100011;
ROM[8557] <= 32'b00000000010000010000000100010011;
ROM[8558] <= 32'b00000000010000010010000000100011;
ROM[8559] <= 32'b00000000010000010000000100010011;
ROM[8560] <= 32'b00000000010100010010000000100011;
ROM[8561] <= 32'b00000000010000010000000100010011;
ROM[8562] <= 32'b00000000011000010010000000100011;
ROM[8563] <= 32'b00000000010000010000000100010011;
ROM[8564] <= 32'b00000001010000000000001110010011;
ROM[8565] <= 32'b00000000100000111000001110010011;
ROM[8566] <= 32'b01000000011100010000001110110011;
ROM[8567] <= 32'b00000000011100000000001000110011;
ROM[8568] <= 32'b00000000001000000000000110110011;
ROM[8569] <= 32'b01011100100000100001000011101111;
ROM[8570] <= 32'b00000110110000000000001110010011;
ROM[8571] <= 32'b00000000011100010010000000100011;
ROM[8572] <= 32'b00000000010000010000000100010011;
ROM[8573] <= 32'b00000000000000001000001110110111;
ROM[8574] <= 32'b01100100000000111000001110010011;
ROM[8575] <= 32'b00000000111000111000001110110011;
ROM[8576] <= 32'b00000000011100010010000000100011;
ROM[8577] <= 32'b00000000010000010000000100010011;
ROM[8578] <= 32'b00000000001100010010000000100011;
ROM[8579] <= 32'b00000000010000010000000100010011;
ROM[8580] <= 32'b00000000010000010010000000100011;
ROM[8581] <= 32'b00000000010000010000000100010011;
ROM[8582] <= 32'b00000000010100010010000000100011;
ROM[8583] <= 32'b00000000010000010000000100010011;
ROM[8584] <= 32'b00000000011000010010000000100011;
ROM[8585] <= 32'b00000000010000010000000100010011;
ROM[8586] <= 32'b00000001010000000000001110010011;
ROM[8587] <= 32'b00000000100000111000001110010011;
ROM[8588] <= 32'b01000000011100010000001110110011;
ROM[8589] <= 32'b00000000011100000000001000110011;
ROM[8590] <= 32'b00000000001000000000000110110011;
ROM[8591] <= 32'b01010111000000100001000011101111;
ROM[8592] <= 32'b00000110111100000000001110010011;
ROM[8593] <= 32'b00000000011100010010000000100011;
ROM[8594] <= 32'b00000000010000010000000100010011;
ROM[8595] <= 32'b00000000000000001000001110110111;
ROM[8596] <= 32'b01101001100000111000001110010011;
ROM[8597] <= 32'b00000000111000111000001110110011;
ROM[8598] <= 32'b00000000011100010010000000100011;
ROM[8599] <= 32'b00000000010000010000000100010011;
ROM[8600] <= 32'b00000000001100010010000000100011;
ROM[8601] <= 32'b00000000010000010000000100010011;
ROM[8602] <= 32'b00000000010000010010000000100011;
ROM[8603] <= 32'b00000000010000010000000100010011;
ROM[8604] <= 32'b00000000010100010010000000100011;
ROM[8605] <= 32'b00000000010000010000000100010011;
ROM[8606] <= 32'b00000000011000010010000000100011;
ROM[8607] <= 32'b00000000010000010000000100010011;
ROM[8608] <= 32'b00000001010000000000001110010011;
ROM[8609] <= 32'b00000000100000111000001110010011;
ROM[8610] <= 32'b01000000011100010000001110110011;
ROM[8611] <= 32'b00000000011100000000001000110011;
ROM[8612] <= 32'b00000000001000000000000110110011;
ROM[8613] <= 32'b01010001100000100001000011101111;
ROM[8614] <= 32'b00000111011100000000001110010011;
ROM[8615] <= 32'b00000000011100010010000000100011;
ROM[8616] <= 32'b00000000010000010000000100010011;
ROM[8617] <= 32'b00000000000000001000001110110111;
ROM[8618] <= 32'b01101111000000111000001110010011;
ROM[8619] <= 32'b00000000111000111000001110110011;
ROM[8620] <= 32'b00000000011100010010000000100011;
ROM[8621] <= 32'b00000000010000010000000100010011;
ROM[8622] <= 32'b00000000001100010010000000100011;
ROM[8623] <= 32'b00000000010000010000000100010011;
ROM[8624] <= 32'b00000000010000010010000000100011;
ROM[8625] <= 32'b00000000010000010000000100010011;
ROM[8626] <= 32'b00000000010100010010000000100011;
ROM[8627] <= 32'b00000000010000010000000100010011;
ROM[8628] <= 32'b00000000011000010010000000100011;
ROM[8629] <= 32'b00000000010000010000000100010011;
ROM[8630] <= 32'b00000001010000000000001110010011;
ROM[8631] <= 32'b00000000100000111000001110010011;
ROM[8632] <= 32'b01000000011100010000001110110011;
ROM[8633] <= 32'b00000000011100000000001000110011;
ROM[8634] <= 32'b00000000001000000000000110110011;
ROM[8635] <= 32'b01001100000000100001000011101111;
ROM[8636] <= 32'b00000110010100000000001110010011;
ROM[8637] <= 32'b00000000011100010010000000100011;
ROM[8638] <= 32'b00000000010000010000000100010011;
ROM[8639] <= 32'b00000000000000001000001110110111;
ROM[8640] <= 32'b01110100100000111000001110010011;
ROM[8641] <= 32'b00000000111000111000001110110011;
ROM[8642] <= 32'b00000000011100010010000000100011;
ROM[8643] <= 32'b00000000010000010000000100010011;
ROM[8644] <= 32'b00000000001100010010000000100011;
ROM[8645] <= 32'b00000000010000010000000100010011;
ROM[8646] <= 32'b00000000010000010010000000100011;
ROM[8647] <= 32'b00000000010000010000000100010011;
ROM[8648] <= 32'b00000000010100010010000000100011;
ROM[8649] <= 32'b00000000010000010000000100010011;
ROM[8650] <= 32'b00000000011000010010000000100011;
ROM[8651] <= 32'b00000000010000010000000100010011;
ROM[8652] <= 32'b00000001010000000000001110010011;
ROM[8653] <= 32'b00000000100000111000001110010011;
ROM[8654] <= 32'b01000000011100010000001110110011;
ROM[8655] <= 32'b00000000011100000000001000110011;
ROM[8656] <= 32'b00000000001000000000000110110011;
ROM[8657] <= 32'b01000110100000100001000011101111;
ROM[8658] <= 32'b00000111001000000000001110010011;
ROM[8659] <= 32'b00000000011100010010000000100011;
ROM[8660] <= 32'b00000000010000010000000100010011;
ROM[8661] <= 32'b00000000000000001000001110110111;
ROM[8662] <= 32'b01111010000000111000001110010011;
ROM[8663] <= 32'b00000000111000111000001110110011;
ROM[8664] <= 32'b00000000011100010010000000100011;
ROM[8665] <= 32'b00000000010000010000000100010011;
ROM[8666] <= 32'b00000000001100010010000000100011;
ROM[8667] <= 32'b00000000010000010000000100010011;
ROM[8668] <= 32'b00000000010000010010000000100011;
ROM[8669] <= 32'b00000000010000010000000100010011;
ROM[8670] <= 32'b00000000010100010010000000100011;
ROM[8671] <= 32'b00000000010000010000000100010011;
ROM[8672] <= 32'b00000000011000010010000000100011;
ROM[8673] <= 32'b00000000010000010000000100010011;
ROM[8674] <= 32'b00000001010000000000001110010011;
ROM[8675] <= 32'b00000000100000111000001110010011;
ROM[8676] <= 32'b01000000011100010000001110110011;
ROM[8677] <= 32'b00000000011100000000001000110011;
ROM[8678] <= 32'b00000000001000000000000110110011;
ROM[8679] <= 32'b01000001000000100001000011101111;
ROM[8680] <= 32'b00000010000000000000001110010011;
ROM[8681] <= 32'b00000000011100010010000000100011;
ROM[8682] <= 32'b00000000010000010000000100010011;
ROM[8683] <= 32'b00000000000000001000001110110111;
ROM[8684] <= 32'b01111111100000111000001110010011;
ROM[8685] <= 32'b00000000111000111000001110110011;
ROM[8686] <= 32'b00000000011100010010000000100011;
ROM[8687] <= 32'b00000000010000010000000100010011;
ROM[8688] <= 32'b00000000001100010010000000100011;
ROM[8689] <= 32'b00000000010000010000000100010011;
ROM[8690] <= 32'b00000000010000010010000000100011;
ROM[8691] <= 32'b00000000010000010000000100010011;
ROM[8692] <= 32'b00000000010100010010000000100011;
ROM[8693] <= 32'b00000000010000010000000100010011;
ROM[8694] <= 32'b00000000011000010010000000100011;
ROM[8695] <= 32'b00000000010000010000000100010011;
ROM[8696] <= 32'b00000001010000000000001110010011;
ROM[8697] <= 32'b00000000100000111000001110010011;
ROM[8698] <= 32'b01000000011100010000001110110011;
ROM[8699] <= 32'b00000000011100000000001000110011;
ROM[8700] <= 32'b00000000001000000000000110110011;
ROM[8701] <= 32'b00111011100000100001000011101111;
ROM[8702] <= 32'b00000110001100000000001110010011;
ROM[8703] <= 32'b00000000011100010010000000100011;
ROM[8704] <= 32'b00000000010000010000000100010011;
ROM[8705] <= 32'b00000000000000001001001110110111;
ROM[8706] <= 32'b10000101000000111000001110010011;
ROM[8707] <= 32'b00000000111000111000001110110011;
ROM[8708] <= 32'b00000000011100010010000000100011;
ROM[8709] <= 32'b00000000010000010000000100010011;
ROM[8710] <= 32'b00000000001100010010000000100011;
ROM[8711] <= 32'b00000000010000010000000100010011;
ROM[8712] <= 32'b00000000010000010010000000100011;
ROM[8713] <= 32'b00000000010000010000000100010011;
ROM[8714] <= 32'b00000000010100010010000000100011;
ROM[8715] <= 32'b00000000010000010000000100010011;
ROM[8716] <= 32'b00000000011000010010000000100011;
ROM[8717] <= 32'b00000000010000010000000100010011;
ROM[8718] <= 32'b00000001010000000000001110010011;
ROM[8719] <= 32'b00000000100000111000001110010011;
ROM[8720] <= 32'b01000000011100010000001110110011;
ROM[8721] <= 32'b00000000011100000000001000110011;
ROM[8722] <= 32'b00000000001000000000000110110011;
ROM[8723] <= 32'b00110110000000100001000011101111;
ROM[8724] <= 32'b00000110000100000000001110010011;
ROM[8725] <= 32'b00000000011100010010000000100011;
ROM[8726] <= 32'b00000000010000010000000100010011;
ROM[8727] <= 32'b00000000000000001001001110110111;
ROM[8728] <= 32'b10001010100000111000001110010011;
ROM[8729] <= 32'b00000000111000111000001110110011;
ROM[8730] <= 32'b00000000011100010010000000100011;
ROM[8731] <= 32'b00000000010000010000000100010011;
ROM[8732] <= 32'b00000000001100010010000000100011;
ROM[8733] <= 32'b00000000010000010000000100010011;
ROM[8734] <= 32'b00000000010000010010000000100011;
ROM[8735] <= 32'b00000000010000010000000100010011;
ROM[8736] <= 32'b00000000010100010010000000100011;
ROM[8737] <= 32'b00000000010000010000000100010011;
ROM[8738] <= 32'b00000000011000010010000000100011;
ROM[8739] <= 32'b00000000010000010000000100010011;
ROM[8740] <= 32'b00000001010000000000001110010011;
ROM[8741] <= 32'b00000000100000111000001110010011;
ROM[8742] <= 32'b01000000011100010000001110110011;
ROM[8743] <= 32'b00000000011100000000001000110011;
ROM[8744] <= 32'b00000000001000000000000110110011;
ROM[8745] <= 32'b00110000100000100001000011101111;
ROM[8746] <= 32'b00000111001100000000001110010011;
ROM[8747] <= 32'b00000000011100010010000000100011;
ROM[8748] <= 32'b00000000010000010000000100010011;
ROM[8749] <= 32'b00000000000000001001001110110111;
ROM[8750] <= 32'b10010000000000111000001110010011;
ROM[8751] <= 32'b00000000111000111000001110110011;
ROM[8752] <= 32'b00000000011100010010000000100011;
ROM[8753] <= 32'b00000000010000010000000100010011;
ROM[8754] <= 32'b00000000001100010010000000100011;
ROM[8755] <= 32'b00000000010000010000000100010011;
ROM[8756] <= 32'b00000000010000010010000000100011;
ROM[8757] <= 32'b00000000010000010000000100010011;
ROM[8758] <= 32'b00000000010100010010000000100011;
ROM[8759] <= 32'b00000000010000010000000100010011;
ROM[8760] <= 32'b00000000011000010010000000100011;
ROM[8761] <= 32'b00000000010000010000000100010011;
ROM[8762] <= 32'b00000001010000000000001110010011;
ROM[8763] <= 32'b00000000100000111000001110010011;
ROM[8764] <= 32'b01000000011100010000001110110011;
ROM[8765] <= 32'b00000000011100000000001000110011;
ROM[8766] <= 32'b00000000001000000000000110110011;
ROM[8767] <= 32'b00101011000000100001000011101111;
ROM[8768] <= 32'b00000110010100000000001110010011;
ROM[8769] <= 32'b00000000011100010010000000100011;
ROM[8770] <= 32'b00000000010000010000000100010011;
ROM[8771] <= 32'b00000000000000001001001110110111;
ROM[8772] <= 32'b10010101100000111000001110010011;
ROM[8773] <= 32'b00000000111000111000001110110011;
ROM[8774] <= 32'b00000000011100010010000000100011;
ROM[8775] <= 32'b00000000010000010000000100010011;
ROM[8776] <= 32'b00000000001100010010000000100011;
ROM[8777] <= 32'b00000000010000010000000100010011;
ROM[8778] <= 32'b00000000010000010010000000100011;
ROM[8779] <= 32'b00000000010000010000000100010011;
ROM[8780] <= 32'b00000000010100010010000000100011;
ROM[8781] <= 32'b00000000010000010000000100010011;
ROM[8782] <= 32'b00000000011000010010000000100011;
ROM[8783] <= 32'b00000000010000010000000100010011;
ROM[8784] <= 32'b00000001010000000000001110010011;
ROM[8785] <= 32'b00000000100000111000001110010011;
ROM[8786] <= 32'b01000000011100010000001110110011;
ROM[8787] <= 32'b00000000011100000000001000110011;
ROM[8788] <= 32'b00000000001000000000000110110011;
ROM[8789] <= 32'b00100101100000100001000011101111;
ROM[8790] <= 32'b00000010100100000000001110010011;
ROM[8791] <= 32'b00000000011100010010000000100011;
ROM[8792] <= 32'b00000000010000010000000100010011;
ROM[8793] <= 32'b00000000000000001001001110110111;
ROM[8794] <= 32'b10011011000000111000001110010011;
ROM[8795] <= 32'b00000000111000111000001110110011;
ROM[8796] <= 32'b00000000011100010010000000100011;
ROM[8797] <= 32'b00000000010000010000000100010011;
ROM[8798] <= 32'b00000000001100010010000000100011;
ROM[8799] <= 32'b00000000010000010000000100010011;
ROM[8800] <= 32'b00000000010000010010000000100011;
ROM[8801] <= 32'b00000000010000010000000100010011;
ROM[8802] <= 32'b00000000010100010010000000100011;
ROM[8803] <= 32'b00000000010000010000000100010011;
ROM[8804] <= 32'b00000000011000010010000000100011;
ROM[8805] <= 32'b00000000010000010000000100010011;
ROM[8806] <= 32'b00000001010000000000001110010011;
ROM[8807] <= 32'b00000000100000111000001110010011;
ROM[8808] <= 32'b01000000011100010000001110110011;
ROM[8809] <= 32'b00000000011100000000001000110011;
ROM[8810] <= 32'b00000000001000000000000110110011;
ROM[8811] <= 32'b00100000000000100001000011101111;
ROM[8812] <= 32'b00000000000000001001001110110111;
ROM[8813] <= 32'b10011111110000111000001110010011;
ROM[8814] <= 32'b00000000111000111000001110110011;
ROM[8815] <= 32'b00000000011100010010000000100011;
ROM[8816] <= 32'b00000000010000010000000100010011;
ROM[8817] <= 32'b00000000001100010010000000100011;
ROM[8818] <= 32'b00000000010000010000000100010011;
ROM[8819] <= 32'b00000000010000010010000000100011;
ROM[8820] <= 32'b00000000010000010000000100010011;
ROM[8821] <= 32'b00000000010100010010000000100011;
ROM[8822] <= 32'b00000000010000010000000100010011;
ROM[8823] <= 32'b00000000011000010010000000100011;
ROM[8824] <= 32'b00000000010000010000000100010011;
ROM[8825] <= 32'b00000001010000000000001110010011;
ROM[8826] <= 32'b00000000010000111000001110010011;
ROM[8827] <= 32'b01000000011100010000001110110011;
ROM[8828] <= 32'b00000000011100000000001000110011;
ROM[8829] <= 32'b00000000001000000000000110110011;
ROM[8830] <= 32'b01010111000000001110000011101111;
ROM[8831] <= 32'b11111111110000010000000100010011;
ROM[8832] <= 32'b00000000000000010010001110000011;
ROM[8833] <= 32'b00000000011101100010000000100011;
ROM[8834] <= 32'b00000000000000001001001110110111;
ROM[8835] <= 32'b10100101010000111000001110010011;
ROM[8836] <= 32'b00000000111000111000001110110011;
ROM[8837] <= 32'b00000000011100010010000000100011;
ROM[8838] <= 32'b00000000010000010000000100010011;
ROM[8839] <= 32'b00000000001100010010000000100011;
ROM[8840] <= 32'b00000000010000010000000100010011;
ROM[8841] <= 32'b00000000010000010010000000100011;
ROM[8842] <= 32'b00000000010000010000000100010011;
ROM[8843] <= 32'b00000000010100010010000000100011;
ROM[8844] <= 32'b00000000010000010000000100010011;
ROM[8845] <= 32'b00000000011000010010000000100011;
ROM[8846] <= 32'b00000000010000010000000100010011;
ROM[8847] <= 32'b00000001010000000000001110010011;
ROM[8848] <= 32'b00000000000000111000001110010011;
ROM[8849] <= 32'b01000000011100010000001110110011;
ROM[8850] <= 32'b00000000011100000000001000110011;
ROM[8851] <= 32'b00000000001000000000000110110011;
ROM[8852] <= 32'b01101001000100000100000011101111;
ROM[8853] <= 32'b11111111110000010000000100010011;
ROM[8854] <= 32'b00000000000000010010001110000011;
ROM[8855] <= 32'b00000000011100011010111000100011;
ROM[8856] <= 32'b00000001110000011010001110000011;
ROM[8857] <= 32'b00000000011100010010000000100011;
ROM[8858] <= 32'b00000000010000010000000100010011;
ROM[8859] <= 32'b00000000000000001001001110110111;
ROM[8860] <= 32'b10101011100000111000001110010011;
ROM[8861] <= 32'b00000000111000111000001110110011;
ROM[8862] <= 32'b00000000011100010010000000100011;
ROM[8863] <= 32'b00000000010000010000000100010011;
ROM[8864] <= 32'b00000000001100010010000000100011;
ROM[8865] <= 32'b00000000010000010000000100010011;
ROM[8866] <= 32'b00000000010000010010000000100011;
ROM[8867] <= 32'b00000000010000010000000100010011;
ROM[8868] <= 32'b00000000010100010010000000100011;
ROM[8869] <= 32'b00000000010000010000000100010011;
ROM[8870] <= 32'b00000000011000010010000000100011;
ROM[8871] <= 32'b00000000010000010000000100010011;
ROM[8872] <= 32'b00000001010000000000001110010011;
ROM[8873] <= 32'b00000000010000111000001110010011;
ROM[8874] <= 32'b01000000011100010000001110110011;
ROM[8875] <= 32'b00000000011100000000001000110011;
ROM[8876] <= 32'b00000000001000000000000110110011;
ROM[8877] <= 32'b10101000000011111011000011101111;
ROM[8878] <= 32'b11111111110000010000000100010011;
ROM[8879] <= 32'b00000000000000010010001110000011;
ROM[8880] <= 32'b00000010011100011010001000100011;
ROM[8881] <= 32'b00000000010000011010001110000011;
ROM[8882] <= 32'b00000000011100010010000000100011;
ROM[8883] <= 32'b00000000010000010000000100010011;
ROM[8884] <= 32'b00000010010000011010001110000011;
ROM[8885] <= 32'b00000000011100010010000000100011;
ROM[8886] <= 32'b00000000010000010000000100010011;
ROM[8887] <= 32'b00000000010000000000001110010011;
ROM[8888] <= 32'b00000000011100010010000000100011;
ROM[8889] <= 32'b00000000010000010000000100010011;
ROM[8890] <= 32'b00000000000000001001001110110111;
ROM[8891] <= 32'b10110011010000111000001110010011;
ROM[8892] <= 32'b00000000111000111000001110110011;
ROM[8893] <= 32'b00000000011100010010000000100011;
ROM[8894] <= 32'b00000000010000010000000100010011;
ROM[8895] <= 32'b00000000001100010010000000100011;
ROM[8896] <= 32'b00000000010000010000000100010011;
ROM[8897] <= 32'b00000000010000010010000000100011;
ROM[8898] <= 32'b00000000010000010000000100010011;
ROM[8899] <= 32'b00000000010100010010000000100011;
ROM[8900] <= 32'b00000000010000010000000100010011;
ROM[8901] <= 32'b00000000011000010010000000100011;
ROM[8902] <= 32'b00000000010000010000000100010011;
ROM[8903] <= 32'b00000001010000000000001110010011;
ROM[8904] <= 32'b00000000100000111000001110010011;
ROM[8905] <= 32'b01000000011100010000001110110011;
ROM[8906] <= 32'b00000000011100000000001000110011;
ROM[8907] <= 32'b00000000001000000000000110110011;
ROM[8908] <= 32'b01001111110100001000000011101111;
ROM[8909] <= 32'b11111111110000010000000100010011;
ROM[8910] <= 32'b00000000000000010010001110000011;
ROM[8911] <= 32'b11111111110000010000000100010011;
ROM[8912] <= 32'b00000000000000010010010000000011;
ROM[8913] <= 32'b00000000011101000000001110110011;
ROM[8914] <= 32'b00000000011100010010000000100011;
ROM[8915] <= 32'b00000000010000010000000100010011;
ROM[8916] <= 32'b11111111110000010000000100010011;
ROM[8917] <= 32'b00000000000000010010001110000011;
ROM[8918] <= 32'b00000000000000111000001100010011;
ROM[8919] <= 32'b00000000110100110000010000110011;
ROM[8920] <= 32'b00000000000001000010001110000011;
ROM[8921] <= 32'b00000000011100010010000000100011;
ROM[8922] <= 32'b00000000010000010000000100010011;
ROM[8923] <= 32'b00000000000100000000001110010011;
ROM[8924] <= 32'b00000000011100010010000000100011;
ROM[8925] <= 32'b00000000010000010000000100010011;
ROM[8926] <= 32'b11111111110000010000000100010011;
ROM[8927] <= 32'b00000000000000010010001110000011;
ROM[8928] <= 32'b11111111110000010000000100010011;
ROM[8929] <= 32'b00000000000000010010010000000011;
ROM[8930] <= 32'b00000000011101000010010010110011;
ROM[8931] <= 32'b00000000100000111010010100110011;
ROM[8932] <= 32'b00000000101001001000001110110011;
ROM[8933] <= 32'b00000000000100111000001110010011;
ROM[8934] <= 32'b00000000000100111111001110010011;
ROM[8935] <= 32'b00000000011100010010000000100011;
ROM[8936] <= 32'b00000000010000010000000100010011;
ROM[8937] <= 32'b11111111110000010000000100010011;
ROM[8938] <= 32'b00000000000000010010001110000011;
ROM[8939] <= 32'b00000000000000111000101001100011;
ROM[8940] <= 32'b00000000000000001100001110110111;
ROM[8941] <= 32'b01100101110000111000001110010011;
ROM[8942] <= 32'b00000000111000111000001110110011;
ROM[8943] <= 32'b00000000000000111000000011100111;
ROM[8944] <= 32'b00000000000100000000001110010011;
ROM[8945] <= 32'b00000000011100010010000000100011;
ROM[8946] <= 32'b00000000010000010000000100010011;
ROM[8947] <= 32'b00000000010000011010001110000011;
ROM[8948] <= 32'b00000000011100010010000000100011;
ROM[8949] <= 32'b00000000010000010000000100010011;
ROM[8950] <= 32'b00000010010000011010001110000011;
ROM[8951] <= 32'b00000000011100010010000000100011;
ROM[8952] <= 32'b00000000010000010000000100010011;
ROM[8953] <= 32'b00000000010000000000001110010011;
ROM[8954] <= 32'b00000000011100010010000000100011;
ROM[8955] <= 32'b00000000010000010000000100010011;
ROM[8956] <= 32'b00000000000000001001001110110111;
ROM[8957] <= 32'b11000011110000111000001110010011;
ROM[8958] <= 32'b00000000111000111000001110110011;
ROM[8959] <= 32'b00000000011100010010000000100011;
ROM[8960] <= 32'b00000000010000010000000100010011;
ROM[8961] <= 32'b00000000001100010010000000100011;
ROM[8962] <= 32'b00000000010000010000000100010011;
ROM[8963] <= 32'b00000000010000010010000000100011;
ROM[8964] <= 32'b00000000010000010000000100010011;
ROM[8965] <= 32'b00000000010100010010000000100011;
ROM[8966] <= 32'b00000000010000010000000100010011;
ROM[8967] <= 32'b00000000011000010010000000100011;
ROM[8968] <= 32'b00000000010000010000000100010011;
ROM[8969] <= 32'b00000001010000000000001110010011;
ROM[8970] <= 32'b00000000100000111000001110010011;
ROM[8971] <= 32'b01000000011100010000001110110011;
ROM[8972] <= 32'b00000000011100000000001000110011;
ROM[8973] <= 32'b00000000001000000000000110110011;
ROM[8974] <= 32'b00111111010100001000000011101111;
ROM[8975] <= 32'b11111111110000010000000100010011;
ROM[8976] <= 32'b00000000000000010010001110000011;
ROM[8977] <= 32'b11111111110000010000000100010011;
ROM[8978] <= 32'b00000000000000010010010000000011;
ROM[8979] <= 32'b00000000011101000000001110110011;
ROM[8980] <= 32'b00000000011100010010000000100011;
ROM[8981] <= 32'b00000000010000010000000100010011;
ROM[8982] <= 32'b11111111110000010000000100010011;
ROM[8983] <= 32'b00000000000000010010001110000011;
ROM[8984] <= 32'b00000000000000111000001100010011;
ROM[8985] <= 32'b11111111110000010000000100010011;
ROM[8986] <= 32'b00000000000000010010001110000011;
ROM[8987] <= 32'b00000000110100110000010000110011;
ROM[8988] <= 32'b00000000011101000010000000100011;
ROM[8989] <= 32'b00000000000000000000001110010011;
ROM[8990] <= 32'b00000000011100010010000000100011;
ROM[8991] <= 32'b00000000010000010000000100010011;
ROM[8992] <= 32'b11111111110000010000000100010011;
ROM[8993] <= 32'b00000000000000010010001110000011;
ROM[8994] <= 32'b00000010011100011010100000100011;
ROM[8995] <= 32'b00000000000000000000001110010011;
ROM[8996] <= 32'b00000000011100010010000000100011;
ROM[8997] <= 32'b00000000010000010000000100010011;
ROM[8998] <= 32'b11111111110000010000000100010011;
ROM[8999] <= 32'b00000000000000010010001110000011;
ROM[9000] <= 32'b00000000011100011010011000100011;
ROM[9001] <= 32'b00000000110000011010001110000011;
ROM[9002] <= 32'b00000000011100010010000000100011;
ROM[9003] <= 32'b00000000010000010000000100010011;
ROM[9004] <= 32'b00000001000000011010001110000011;
ROM[9005] <= 32'b00000000011100010010000000100011;
ROM[9006] <= 32'b00000000010000010000000100010011;
ROM[9007] <= 32'b11111111110000010000000100010011;
ROM[9008] <= 32'b00000000000000010010001110000011;
ROM[9009] <= 32'b11111111110000010000000100010011;
ROM[9010] <= 32'b00000000000000010010010000000011;
ROM[9011] <= 32'b00000000011101000010001110110011;
ROM[9012] <= 32'b00000000011100010010000000100011;
ROM[9013] <= 32'b00000000010000010000000100010011;
ROM[9014] <= 32'b11111111110000010000000100010011;
ROM[9015] <= 32'b00000000000000010010001110000011;
ROM[9016] <= 32'b01000000011100000000001110110011;
ROM[9017] <= 32'b00000000000100111000001110010011;
ROM[9018] <= 32'b00000000011100010010000000100011;
ROM[9019] <= 32'b00000000010000010000000100010011;
ROM[9020] <= 32'b11111111110000010000000100010011;
ROM[9021] <= 32'b00000000000000010010001110000011;
ROM[9022] <= 32'b00000000000000111000101001100011;
ROM[9023] <= 32'b00000000000000001001001110110111;
ROM[9024] <= 32'b00000001110000111000001110010011;
ROM[9025] <= 32'b00000000111000111000001110110011;
ROM[9026] <= 32'b00000000000000111000000011100111;
ROM[9027] <= 32'b00000000000000011010001110000011;
ROM[9028] <= 32'b00000000011100010010000000100011;
ROM[9029] <= 32'b00000000010000010000000100010011;
ROM[9030] <= 32'b00000000100000011010001110000011;
ROM[9031] <= 32'b00000000011100010010000000100011;
ROM[9032] <= 32'b00000000010000010000000100010011;
ROM[9033] <= 32'b00000000010000000000001110010011;
ROM[9034] <= 32'b00000000011100010010000000100011;
ROM[9035] <= 32'b00000000010000010000000100010011;
ROM[9036] <= 32'b00000000000000001001001110110111;
ROM[9037] <= 32'b11010111110000111000001110010011;
ROM[9038] <= 32'b00000000111000111000001110110011;
ROM[9039] <= 32'b00000000011100010010000000100011;
ROM[9040] <= 32'b00000000010000010000000100010011;
ROM[9041] <= 32'b00000000001100010010000000100011;
ROM[9042] <= 32'b00000000010000010000000100010011;
ROM[9043] <= 32'b00000000010000010010000000100011;
ROM[9044] <= 32'b00000000010000010000000100010011;
ROM[9045] <= 32'b00000000010100010010000000100011;
ROM[9046] <= 32'b00000000010000010000000100010011;
ROM[9047] <= 32'b00000000011000010010000000100011;
ROM[9048] <= 32'b00000000010000010000000100010011;
ROM[9049] <= 32'b00000001010000000000001110010011;
ROM[9050] <= 32'b00000000100000111000001110010011;
ROM[9051] <= 32'b01000000011100010000001110110011;
ROM[9052] <= 32'b00000000011100000000001000110011;
ROM[9053] <= 32'b00000000001000000000000110110011;
ROM[9054] <= 32'b00101011010100001000000011101111;
ROM[9055] <= 32'b11111111110000010000000100010011;
ROM[9056] <= 32'b00000000000000010010001110000011;
ROM[9057] <= 32'b11111111110000010000000100010011;
ROM[9058] <= 32'b00000000000000010010010000000011;
ROM[9059] <= 32'b00000000011101000000001110110011;
ROM[9060] <= 32'b00000000011100010010000000100011;
ROM[9061] <= 32'b00000000010000010000000100010011;
ROM[9062] <= 32'b11111111110000010000000100010011;
ROM[9063] <= 32'b00000000000000010010001110000011;
ROM[9064] <= 32'b00000000000000111000001100010011;
ROM[9065] <= 32'b00000000110100110000010000110011;
ROM[9066] <= 32'b00000000000001000010001110000011;
ROM[9067] <= 32'b00000000011100010010000000100011;
ROM[9068] <= 32'b00000000010000010000000100010011;
ROM[9069] <= 32'b11111111110000010000000100010011;
ROM[9070] <= 32'b00000000000000010010001110000011;
ROM[9071] <= 32'b00000010011100011010110000100011;
ROM[9072] <= 32'b00000011100000011010001110000011;
ROM[9073] <= 32'b00000000011100010010000000100011;
ROM[9074] <= 32'b00000000010000010000000100010011;
ROM[9075] <= 32'b00000000110000011010001110000011;
ROM[9076] <= 32'b00000000011100010010000000100011;
ROM[9077] <= 32'b00000000010000010000000100010011;
ROM[9078] <= 32'b00000000010000000000001110010011;
ROM[9079] <= 32'b00000000011100010010000000100011;
ROM[9080] <= 32'b00000000010000010000000100010011;
ROM[9081] <= 32'b00000000000000001001001110110111;
ROM[9082] <= 32'b11100011000000111000001110010011;
ROM[9083] <= 32'b00000000111000111000001110110011;
ROM[9084] <= 32'b00000000011100010010000000100011;
ROM[9085] <= 32'b00000000010000010000000100010011;
ROM[9086] <= 32'b00000000001100010010000000100011;
ROM[9087] <= 32'b00000000010000010000000100010011;
ROM[9088] <= 32'b00000000010000010010000000100011;
ROM[9089] <= 32'b00000000010000010000000100010011;
ROM[9090] <= 32'b00000000010100010010000000100011;
ROM[9091] <= 32'b00000000010000010000000100010011;
ROM[9092] <= 32'b00000000011000010010000000100011;
ROM[9093] <= 32'b00000000010000010000000100010011;
ROM[9094] <= 32'b00000001010000000000001110010011;
ROM[9095] <= 32'b00000000100000111000001110010011;
ROM[9096] <= 32'b01000000011100010000001110110011;
ROM[9097] <= 32'b00000000011100000000001000110011;
ROM[9098] <= 32'b00000000001000000000000110110011;
ROM[9099] <= 32'b00100000000100001000000011101111;
ROM[9100] <= 32'b00000000000000001001001110110111;
ROM[9101] <= 32'b11100111110000111000001110010011;
ROM[9102] <= 32'b00000000111000111000001110110011;
ROM[9103] <= 32'b00000000011100010010000000100011;
ROM[9104] <= 32'b00000000010000010000000100010011;
ROM[9105] <= 32'b00000000001100010010000000100011;
ROM[9106] <= 32'b00000000010000010000000100010011;
ROM[9107] <= 32'b00000000010000010010000000100011;
ROM[9108] <= 32'b00000000010000010000000100010011;
ROM[9109] <= 32'b00000000010100010010000000100011;
ROM[9110] <= 32'b00000000010000010000000100010011;
ROM[9111] <= 32'b00000000011000010010000000100011;
ROM[9112] <= 32'b00000000010000010000000100010011;
ROM[9113] <= 32'b00000001010000000000001110010011;
ROM[9114] <= 32'b00000000100000111000001110010011;
ROM[9115] <= 32'b01000000011100010000001110110011;
ROM[9116] <= 32'b00000000011100000000001000110011;
ROM[9117] <= 32'b00000000001000000000000110110011;
ROM[9118] <= 32'b00101110010100100000000011101111;
ROM[9119] <= 32'b11111111110000010000000100010011;
ROM[9120] <= 32'b00000000000000010010001110000011;
ROM[9121] <= 32'b00000010011100011010010000100011;
ROM[9122] <= 32'b00000010100000011010001110000011;
ROM[9123] <= 32'b00000000011100010010000000100011;
ROM[9124] <= 32'b00000000010000010000000100010011;
ROM[9125] <= 32'b00000001110000011010001110000011;
ROM[9126] <= 32'b00000000011100010010000000100011;
ROM[9127] <= 32'b00000000010000010000000100010011;
ROM[9128] <= 32'b11111111110000010000000100010011;
ROM[9129] <= 32'b00000000000000010010001110000011;
ROM[9130] <= 32'b11111111110000010000000100010011;
ROM[9131] <= 32'b00000000000000010010010000000011;
ROM[9132] <= 32'b00000000011101000010010010110011;
ROM[9133] <= 32'b00000000100000111010010100110011;
ROM[9134] <= 32'b00000000101001001000001110110011;
ROM[9135] <= 32'b00000000000100111000001110010011;
ROM[9136] <= 32'b00000000000100111111001110010011;
ROM[9137] <= 32'b00000000011100010010000000100011;
ROM[9138] <= 32'b00000000010000010000000100010011;
ROM[9139] <= 32'b11111111110000010000000100010011;
ROM[9140] <= 32'b00000000000000010010001110000011;
ROM[9141] <= 32'b00000000000000111000101001100011;
ROM[9142] <= 32'b00000000000000001001001110110111;
ROM[9143] <= 32'b11101110110000111000001110010011;
ROM[9144] <= 32'b00000000111000111000001110110011;
ROM[9145] <= 32'b00000000000000111000000011100111;
ROM[9146] <= 32'b00001111000000000000000011101111;
ROM[9147] <= 32'b00000000000100000000001110010011;
ROM[9148] <= 32'b00000000011100010010000000100011;
ROM[9149] <= 32'b00000000010000010000000100010011;
ROM[9150] <= 32'b11111111110000010000000100010011;
ROM[9151] <= 32'b00000000000000010010001110000011;
ROM[9152] <= 32'b00000010011100011010100000100011;
ROM[9153] <= 32'b00000001100000011010001110000011;
ROM[9154] <= 32'b00000000011100010010000000100011;
ROM[9155] <= 32'b00000000010000010000000100010011;
ROM[9156] <= 32'b00000000110000011010001110000011;
ROM[9157] <= 32'b00000000011100010010000000100011;
ROM[9158] <= 32'b00000000010000010000000100010011;
ROM[9159] <= 32'b00000000010000000000001110010011;
ROM[9160] <= 32'b00000000011100010010000000100011;
ROM[9161] <= 32'b00000000010000010000000100010011;
ROM[9162] <= 32'b00000000000000001001001110110111;
ROM[9163] <= 32'b11110111010000111000001110010011;
ROM[9164] <= 32'b00000000111000111000001110110011;
ROM[9165] <= 32'b00000000011100010010000000100011;
ROM[9166] <= 32'b00000000010000010000000100010011;
ROM[9167] <= 32'b00000000001100010010000000100011;
ROM[9168] <= 32'b00000000010000010000000100010011;
ROM[9169] <= 32'b00000000010000010010000000100011;
ROM[9170] <= 32'b00000000010000010000000100010011;
ROM[9171] <= 32'b00000000010100010010000000100011;
ROM[9172] <= 32'b00000000010000010000000100010011;
ROM[9173] <= 32'b00000000011000010010000000100011;
ROM[9174] <= 32'b00000000010000010000000100010011;
ROM[9175] <= 32'b00000001010000000000001110010011;
ROM[9176] <= 32'b00000000100000111000001110010011;
ROM[9177] <= 32'b01000000011100010000001110110011;
ROM[9178] <= 32'b00000000011100000000001000110011;
ROM[9179] <= 32'b00000000001000000000000110110011;
ROM[9180] <= 32'b00001011110100001000000011101111;
ROM[9181] <= 32'b00000001110000011010001110000011;
ROM[9182] <= 32'b00000000011100010010000000100011;
ROM[9183] <= 32'b00000000010000010000000100010011;
ROM[9184] <= 32'b00000000000000001001001110110111;
ROM[9185] <= 32'b11111100110000111000001110010011;
ROM[9186] <= 32'b00000000111000111000001110110011;
ROM[9187] <= 32'b00000000011100010010000000100011;
ROM[9188] <= 32'b00000000010000010000000100010011;
ROM[9189] <= 32'b00000000001100010010000000100011;
ROM[9190] <= 32'b00000000010000010000000100010011;
ROM[9191] <= 32'b00000000010000010010000000100011;
ROM[9192] <= 32'b00000000010000010000000100010011;
ROM[9193] <= 32'b00000000010100010010000000100011;
ROM[9194] <= 32'b00000000010000010000000100010011;
ROM[9195] <= 32'b00000000011000010010000000100011;
ROM[9196] <= 32'b00000000010000010000000100010011;
ROM[9197] <= 32'b00000001010000000000001110010011;
ROM[9198] <= 32'b00000000110000111000001110010011;
ROM[9199] <= 32'b01000000011100010000001110110011;
ROM[9200] <= 32'b00000000011100000000001000110011;
ROM[9201] <= 32'b00000000001000000000000110110011;
ROM[9202] <= 32'b00101011000100100000000011101111;
ROM[9203] <= 32'b11111111110000010000000100010011;
ROM[9204] <= 32'b00000000000000010010001110000011;
ROM[9205] <= 32'b00000000011101100010000000100011;
ROM[9206] <= 32'b00000000110000011010001110000011;
ROM[9207] <= 32'b00000000011100010010000000100011;
ROM[9208] <= 32'b00000000010000010000000100010011;
ROM[9209] <= 32'b00000000000100000000001110010011;
ROM[9210] <= 32'b00000000011100010010000000100011;
ROM[9211] <= 32'b00000000010000010000000100010011;
ROM[9212] <= 32'b11111111110000010000000100010011;
ROM[9213] <= 32'b00000000000000010010001110000011;
ROM[9214] <= 32'b11111111110000010000000100010011;
ROM[9215] <= 32'b00000000000000010010010000000011;
ROM[9216] <= 32'b00000000011101000000001110110011;
ROM[9217] <= 32'b00000000011100010010000000100011;
ROM[9218] <= 32'b00000000010000010000000100010011;
ROM[9219] <= 32'b11111111110000010000000100010011;
ROM[9220] <= 32'b00000000000000010010001110000011;
ROM[9221] <= 32'b00000000011100011010011000100011;
ROM[9222] <= 32'b11001000110111111111000011101111;
ROM[9223] <= 32'b00000011000000011010001110000011;
ROM[9224] <= 32'b00000000011100010010000000100011;
ROM[9225] <= 32'b00000000010000010000000100010011;
ROM[9226] <= 32'b00000000000000000000001110010011;
ROM[9227] <= 32'b00000000011100010010000000100011;
ROM[9228] <= 32'b00000000010000010000000100010011;
ROM[9229] <= 32'b11111111110000010000000100010011;
ROM[9230] <= 32'b00000000000000010010001110000011;
ROM[9231] <= 32'b11111111110000010000000100010011;
ROM[9232] <= 32'b00000000000000010010010000000011;
ROM[9233] <= 32'b00000000011101000010010010110011;
ROM[9234] <= 32'b00000000100000111010010100110011;
ROM[9235] <= 32'b00000000101001001000001110110011;
ROM[9236] <= 32'b00000000000100111000001110010011;
ROM[9237] <= 32'b00000000000100111111001110010011;
ROM[9238] <= 32'b00000000011100010010000000100011;
ROM[9239] <= 32'b00000000010000010000000100010011;
ROM[9240] <= 32'b11111111110000010000000100010011;
ROM[9241] <= 32'b00000000000000010010001110000011;
ROM[9242] <= 32'b00000000000000111000101001100011;
ROM[9243] <= 32'b00000000000000001010001110110111;
ROM[9244] <= 32'b01101100000000111000001110010011;
ROM[9245] <= 32'b00000000111000111000001110110011;
ROM[9246] <= 32'b00000000000000111000000011100111;
ROM[9247] <= 32'b00000000000000000000001110010011;
ROM[9248] <= 32'b00000000011100010010000000100011;
ROM[9249] <= 32'b00000000010000010000000100010011;
ROM[9250] <= 32'b11111111110000010000000100010011;
ROM[9251] <= 32'b00000000000000010010001110000011;
ROM[9252] <= 32'b00000010011100011010101000100011;
ROM[9253] <= 32'b00000000000000000000001110010011;
ROM[9254] <= 32'b00000000011100010010000000100011;
ROM[9255] <= 32'b00000000010000010000000100010011;
ROM[9256] <= 32'b11111111110000010000000100010011;
ROM[9257] <= 32'b00000000000000010010001110000011;
ROM[9258] <= 32'b00000000011100011010011000100011;
ROM[9259] <= 32'b00000000110000011010001110000011;
ROM[9260] <= 32'b00000000011100010010000000100011;
ROM[9261] <= 32'b00000000010000010000000100010011;
ROM[9262] <= 32'b00000001000000011010001110000011;
ROM[9263] <= 32'b00000000011100010010000000100011;
ROM[9264] <= 32'b00000000010000010000000100010011;
ROM[9265] <= 32'b11111111110000010000000100010011;
ROM[9266] <= 32'b00000000000000010010001110000011;
ROM[9267] <= 32'b11111111110000010000000100010011;
ROM[9268] <= 32'b00000000000000010010010000000011;
ROM[9269] <= 32'b00000000011101000010001110110011;
ROM[9270] <= 32'b00000000011100010010000000100011;
ROM[9271] <= 32'b00000000010000010000000100010011;
ROM[9272] <= 32'b11111111110000010000000100010011;
ROM[9273] <= 32'b00000000000000010010001110000011;
ROM[9274] <= 32'b01000000011100000000001110110011;
ROM[9275] <= 32'b00000000000100111000001110010011;
ROM[9276] <= 32'b00000000011100010010000000100011;
ROM[9277] <= 32'b00000000010000010000000100010011;
ROM[9278] <= 32'b11111111110000010000000100010011;
ROM[9279] <= 32'b00000000000000010010001110000011;
ROM[9280] <= 32'b00000000000000111000101001100011;
ROM[9281] <= 32'b00000000000000001001001110110111;
ROM[9282] <= 32'b00101001110000111000001110010011;
ROM[9283] <= 32'b00000000111000111000001110110011;
ROM[9284] <= 32'b00000000000000111000000011100111;
ROM[9285] <= 32'b00000001100000011010001110000011;
ROM[9286] <= 32'b00000000011100010010000000100011;
ROM[9287] <= 32'b00000000010000010000000100010011;
ROM[9288] <= 32'b00000000110000011010001110000011;
ROM[9289] <= 32'b00000000011100010010000000100011;
ROM[9290] <= 32'b00000000010000010000000100010011;
ROM[9291] <= 32'b00000000010000000000001110010011;
ROM[9292] <= 32'b00000000011100010010000000100011;
ROM[9293] <= 32'b00000000010000010000000100010011;
ROM[9294] <= 32'b00000000000000001001001110110111;
ROM[9295] <= 32'b00011000010000111000001110010011;
ROM[9296] <= 32'b00000000111000111000001110110011;
ROM[9297] <= 32'b00000000011100010010000000100011;
ROM[9298] <= 32'b00000000010000010000000100010011;
ROM[9299] <= 32'b00000000001100010010000000100011;
ROM[9300] <= 32'b00000000010000010000000100010011;
ROM[9301] <= 32'b00000000010000010010000000100011;
ROM[9302] <= 32'b00000000010000010000000100010011;
ROM[9303] <= 32'b00000000010100010010000000100011;
ROM[9304] <= 32'b00000000010000010000000100010011;
ROM[9305] <= 32'b00000000011000010010000000100011;
ROM[9306] <= 32'b00000000010000010000000100010011;
ROM[9307] <= 32'b00000001010000000000001110010011;
ROM[9308] <= 32'b00000000100000111000001110010011;
ROM[9309] <= 32'b01000000011100010000001110110011;
ROM[9310] <= 32'b00000000011100000000001000110011;
ROM[9311] <= 32'b00000000001000000000000110110011;
ROM[9312] <= 32'b01101010110000001000000011101111;
ROM[9313] <= 32'b00000000000000001001001110110111;
ROM[9314] <= 32'b00011101000000111000001110010011;
ROM[9315] <= 32'b00000000111000111000001110110011;
ROM[9316] <= 32'b00000000011100010010000000100011;
ROM[9317] <= 32'b00000000010000010000000100010011;
ROM[9318] <= 32'b00000000001100010010000000100011;
ROM[9319] <= 32'b00000000010000010000000100010011;
ROM[9320] <= 32'b00000000010000010010000000100011;
ROM[9321] <= 32'b00000000010000010000000100010011;
ROM[9322] <= 32'b00000000010100010010000000100011;
ROM[9323] <= 32'b00000000010000010000000100010011;
ROM[9324] <= 32'b00000000011000010010000000100011;
ROM[9325] <= 32'b00000000010000010000000100010011;
ROM[9326] <= 32'b00000001010000000000001110010011;
ROM[9327] <= 32'b00000000100000111000001110010011;
ROM[9328] <= 32'b01000000011100010000001110110011;
ROM[9329] <= 32'b00000000011100000000001000110011;
ROM[9330] <= 32'b00000000001000000000000110110011;
ROM[9331] <= 32'b01111001000000100000000011101111;
ROM[9332] <= 32'b11111111110000010000000100010011;
ROM[9333] <= 32'b00000000000000010010001110000011;
ROM[9334] <= 32'b00000010011100011010010000100011;
ROM[9335] <= 32'b00000010100000011010001110000011;
ROM[9336] <= 32'b00000000011100010010000000100011;
ROM[9337] <= 32'b00000000010000010000000100010011;
ROM[9338] <= 32'b00000010110000011010001110000011;
ROM[9339] <= 32'b00000000011100010010000000100011;
ROM[9340] <= 32'b00000000010000010000000100010011;
ROM[9341] <= 32'b11111111110000010000000100010011;
ROM[9342] <= 32'b00000000000000010010001110000011;
ROM[9343] <= 32'b11111111110000010000000100010011;
ROM[9344] <= 32'b00000000000000010010010000000011;
ROM[9345] <= 32'b00000000011101000010010010110011;
ROM[9346] <= 32'b00000000100000111010010100110011;
ROM[9347] <= 32'b00000000101001001000001110110011;
ROM[9348] <= 32'b00000000000100111000001110010011;
ROM[9349] <= 32'b00000000000100111111001110010011;
ROM[9350] <= 32'b00000000011100010010000000100011;
ROM[9351] <= 32'b00000000010000010000000100010011;
ROM[9352] <= 32'b11111111110000010000000100010011;
ROM[9353] <= 32'b00000000000000010010001110000011;
ROM[9354] <= 32'b00000000000000111000101001100011;
ROM[9355] <= 32'b00000000000000001001001110110111;
ROM[9356] <= 32'b00100100000000111000001110010011;
ROM[9357] <= 32'b00000000111000111000001110110011;
ROM[9358] <= 32'b00000000000000111000000011100111;
ROM[9359] <= 32'b00000001110000000000000011101111;
ROM[9360] <= 32'b00000000000100000000001110010011;
ROM[9361] <= 32'b00000000011100010010000000100011;
ROM[9362] <= 32'b00000000010000010000000100010011;
ROM[9363] <= 32'b11111111110000010000000100010011;
ROM[9364] <= 32'b00000000000000010010001110000011;
ROM[9365] <= 32'b00000010011100011010101000100011;
ROM[9366] <= 32'b00000000110000011010001110000011;
ROM[9367] <= 32'b00000000011100010010000000100011;
ROM[9368] <= 32'b00000000010000010000000100010011;
ROM[9369] <= 32'b00000000000100000000001110010011;
ROM[9370] <= 32'b00000000011100010010000000100011;
ROM[9371] <= 32'b00000000010000010000000100010011;
ROM[9372] <= 32'b11111111110000010000000100010011;
ROM[9373] <= 32'b00000000000000010010001110000011;
ROM[9374] <= 32'b11111111110000010000000100010011;
ROM[9375] <= 32'b00000000000000010010010000000011;
ROM[9376] <= 32'b00000000011101000000001110110011;
ROM[9377] <= 32'b00000000011100010010000000100011;
ROM[9378] <= 32'b00000000010000010000000100010011;
ROM[9379] <= 32'b11111111110000010000000100010011;
ROM[9380] <= 32'b00000000000000010010001110000011;
ROM[9381] <= 32'b00000000011100011010011000100011;
ROM[9382] <= 32'b11100001010111111111000011101111;
ROM[9383] <= 32'b00000011010000011010001110000011;
ROM[9384] <= 32'b00000000011100010010000000100011;
ROM[9385] <= 32'b00000000010000010000000100010011;
ROM[9386] <= 32'b00000000000000000000001110010011;
ROM[9387] <= 32'b00000000011100010010000000100011;
ROM[9388] <= 32'b00000000010000010000000100010011;
ROM[9389] <= 32'b11111111110000010000000100010011;
ROM[9390] <= 32'b00000000000000010010001110000011;
ROM[9391] <= 32'b11111111110000010000000100010011;
ROM[9392] <= 32'b00000000000000010010010000000011;
ROM[9393] <= 32'b00000000011101000010010010110011;
ROM[9394] <= 32'b00000000100000111010010100110011;
ROM[9395] <= 32'b00000000101001001000001110110011;
ROM[9396] <= 32'b00000000000100111000001110010011;
ROM[9397] <= 32'b00000000000100111111001110010011;
ROM[9398] <= 32'b00000000011100010010000000100011;
ROM[9399] <= 32'b00000000010000010000000100010011;
ROM[9400] <= 32'b11111111110000010000000100010011;
ROM[9401] <= 32'b00000000000000010010001110000011;
ROM[9402] <= 32'b00000000000000111000101001100011;
ROM[9403] <= 32'b00000000000000001001001110110111;
ROM[9404] <= 32'b00110000000000111000001110010011;
ROM[9405] <= 32'b00000000111000111000001110110011;
ROM[9406] <= 32'b00000000000000111000000011100111;
ROM[9407] <= 32'b00111100000000000001000011101111;
ROM[9408] <= 32'b00000000000100000000001110010011;
ROM[9409] <= 32'b00000000011100010010000000100011;
ROM[9410] <= 32'b00000000010000010000000100010011;
ROM[9411] <= 32'b11111111110000010000000100010011;
ROM[9412] <= 32'b00000000000000010010001110000011;
ROM[9413] <= 32'b00000010011100011010000000100011;
ROM[9414] <= 32'b00000010011000000000001110010011;
ROM[9415] <= 32'b00000000011100010010000000100011;
ROM[9416] <= 32'b00000000010000010000000100010011;
ROM[9417] <= 32'b00000000000000001001001110110111;
ROM[9418] <= 32'b00110111000000111000001110010011;
ROM[9419] <= 32'b00000000111000111000001110110011;
ROM[9420] <= 32'b00000000011100010010000000100011;
ROM[9421] <= 32'b00000000010000010000000100010011;
ROM[9422] <= 32'b00000000001100010010000000100011;
ROM[9423] <= 32'b00000000010000010000000100010011;
ROM[9424] <= 32'b00000000010000010010000000100011;
ROM[9425] <= 32'b00000000010000010000000100010011;
ROM[9426] <= 32'b00000000010100010010000000100011;
ROM[9427] <= 32'b00000000010000010000000100010011;
ROM[9428] <= 32'b00000000011000010010000000100011;
ROM[9429] <= 32'b00000000010000010000000100010011;
ROM[9430] <= 32'b00000001010000000000001110010011;
ROM[9431] <= 32'b00000000010000111000001110010011;
ROM[9432] <= 32'b01000000011100010000001110110011;
ROM[9433] <= 32'b00000000011100000000001000110011;
ROM[9434] <= 32'b00000000001000000000000110110011;
ROM[9435] <= 32'b00111101000000100000000011101111;
ROM[9436] <= 32'b00000110001100000000001110010011;
ROM[9437] <= 32'b00000000011100010010000000100011;
ROM[9438] <= 32'b00000000010000010000000100010011;
ROM[9439] <= 32'b00000000000000001001001110110111;
ROM[9440] <= 32'b00111100100000111000001110010011;
ROM[9441] <= 32'b00000000111000111000001110110011;
ROM[9442] <= 32'b00000000011100010010000000100011;
ROM[9443] <= 32'b00000000010000010000000100010011;
ROM[9444] <= 32'b00000000001100010010000000100011;
ROM[9445] <= 32'b00000000010000010000000100010011;
ROM[9446] <= 32'b00000000010000010010000000100011;
ROM[9447] <= 32'b00000000010000010000000100010011;
ROM[9448] <= 32'b00000000010100010010000000100011;
ROM[9449] <= 32'b00000000010000010000000100010011;
ROM[9450] <= 32'b00000000011000010010000000100011;
ROM[9451] <= 32'b00000000010000010000000100010011;
ROM[9452] <= 32'b00000001010000000000001110010011;
ROM[9453] <= 32'b00000000100000111000001110010011;
ROM[9454] <= 32'b01000000011100010000001110110011;
ROM[9455] <= 32'b00000000011100000000001000110011;
ROM[9456] <= 32'b00000000001000000000000110110011;
ROM[9457] <= 32'b01111110100000100000000011101111;
ROM[9458] <= 32'b00000110111100000000001110010011;
ROM[9459] <= 32'b00000000011100010010000000100011;
ROM[9460] <= 32'b00000000010000010000000100010011;
ROM[9461] <= 32'b00000000000000001001001110110111;
ROM[9462] <= 32'b01000010000000111000001110010011;
ROM[9463] <= 32'b00000000111000111000001110110011;
ROM[9464] <= 32'b00000000011100010010000000100011;
ROM[9465] <= 32'b00000000010000010000000100010011;
ROM[9466] <= 32'b00000000001100010010000000100011;
ROM[9467] <= 32'b00000000010000010000000100010011;
ROM[9468] <= 32'b00000000010000010010000000100011;
ROM[9469] <= 32'b00000000010000010000000100010011;
ROM[9470] <= 32'b00000000010100010010000000100011;
ROM[9471] <= 32'b00000000010000010000000100010011;
ROM[9472] <= 32'b00000000011000010010000000100011;
ROM[9473] <= 32'b00000000010000010000000100010011;
ROM[9474] <= 32'b00000001010000000000001110010011;
ROM[9475] <= 32'b00000000100000111000001110010011;
ROM[9476] <= 32'b01000000011100010000001110110011;
ROM[9477] <= 32'b00000000011100000000001000110011;
ROM[9478] <= 32'b00000000001000000000000110110011;
ROM[9479] <= 32'b01111001000000100000000011101111;
ROM[9480] <= 32'b00000110111000000000001110010011;
ROM[9481] <= 32'b00000000011100010010000000100011;
ROM[9482] <= 32'b00000000010000010000000100010011;
ROM[9483] <= 32'b00000000000000001001001110110111;
ROM[9484] <= 32'b01000111100000111000001110010011;
ROM[9485] <= 32'b00000000111000111000001110110011;
ROM[9486] <= 32'b00000000011100010010000000100011;
ROM[9487] <= 32'b00000000010000010000000100010011;
ROM[9488] <= 32'b00000000001100010010000000100011;
ROM[9489] <= 32'b00000000010000010000000100010011;
ROM[9490] <= 32'b00000000010000010010000000100011;
ROM[9491] <= 32'b00000000010000010000000100010011;
ROM[9492] <= 32'b00000000010100010010000000100011;
ROM[9493] <= 32'b00000000010000010000000100010011;
ROM[9494] <= 32'b00000000011000010010000000100011;
ROM[9495] <= 32'b00000000010000010000000100010011;
ROM[9496] <= 32'b00000001010000000000001110010011;
ROM[9497] <= 32'b00000000100000111000001110010011;
ROM[9498] <= 32'b01000000011100010000001110110011;
ROM[9499] <= 32'b00000000011100000000001000110011;
ROM[9500] <= 32'b00000000001000000000000110110011;
ROM[9501] <= 32'b01110011100000100000000011101111;
ROM[9502] <= 32'b00000110011100000000001110010011;
ROM[9503] <= 32'b00000000011100010010000000100011;
ROM[9504] <= 32'b00000000010000010000000100010011;
ROM[9505] <= 32'b00000000000000001001001110110111;
ROM[9506] <= 32'b01001101000000111000001110010011;
ROM[9507] <= 32'b00000000111000111000001110110011;
ROM[9508] <= 32'b00000000011100010010000000100011;
ROM[9509] <= 32'b00000000010000010000000100010011;
ROM[9510] <= 32'b00000000001100010010000000100011;
ROM[9511] <= 32'b00000000010000010000000100010011;
ROM[9512] <= 32'b00000000010000010010000000100011;
ROM[9513] <= 32'b00000000010000010000000100010011;
ROM[9514] <= 32'b00000000010100010010000000100011;
ROM[9515] <= 32'b00000000010000010000000100010011;
ROM[9516] <= 32'b00000000011000010010000000100011;
ROM[9517] <= 32'b00000000010000010000000100010011;
ROM[9518] <= 32'b00000001010000000000001110010011;
ROM[9519] <= 32'b00000000100000111000001110010011;
ROM[9520] <= 32'b01000000011100010000001110110011;
ROM[9521] <= 32'b00000000011100000000001000110011;
ROM[9522] <= 32'b00000000001000000000000110110011;
ROM[9523] <= 32'b01101110000000100000000011101111;
ROM[9524] <= 32'b00000111001000000000001110010011;
ROM[9525] <= 32'b00000000011100010010000000100011;
ROM[9526] <= 32'b00000000010000010000000100010011;
ROM[9527] <= 32'b00000000000000001001001110110111;
ROM[9528] <= 32'b01010010100000111000001110010011;
ROM[9529] <= 32'b00000000111000111000001110110011;
ROM[9530] <= 32'b00000000011100010010000000100011;
ROM[9531] <= 32'b00000000010000010000000100010011;
ROM[9532] <= 32'b00000000001100010010000000100011;
ROM[9533] <= 32'b00000000010000010000000100010011;
ROM[9534] <= 32'b00000000010000010010000000100011;
ROM[9535] <= 32'b00000000010000010000000100010011;
ROM[9536] <= 32'b00000000010100010010000000100011;
ROM[9537] <= 32'b00000000010000010000000100010011;
ROM[9538] <= 32'b00000000011000010010000000100011;
ROM[9539] <= 32'b00000000010000010000000100010011;
ROM[9540] <= 32'b00000001010000000000001110010011;
ROM[9541] <= 32'b00000000100000111000001110010011;
ROM[9542] <= 32'b01000000011100010000001110110011;
ROM[9543] <= 32'b00000000011100000000001000110011;
ROM[9544] <= 32'b00000000001000000000000110110011;
ROM[9545] <= 32'b01101000100000100000000011101111;
ROM[9546] <= 32'b00000110000100000000001110010011;
ROM[9547] <= 32'b00000000011100010010000000100011;
ROM[9548] <= 32'b00000000010000010000000100010011;
ROM[9549] <= 32'b00000000000000001001001110110111;
ROM[9550] <= 32'b01011000000000111000001110010011;
ROM[9551] <= 32'b00000000111000111000001110110011;
ROM[9552] <= 32'b00000000011100010010000000100011;
ROM[9553] <= 32'b00000000010000010000000100010011;
ROM[9554] <= 32'b00000000001100010010000000100011;
ROM[9555] <= 32'b00000000010000010000000100010011;
ROM[9556] <= 32'b00000000010000010010000000100011;
ROM[9557] <= 32'b00000000010000010000000100010011;
ROM[9558] <= 32'b00000000010100010010000000100011;
ROM[9559] <= 32'b00000000010000010000000100010011;
ROM[9560] <= 32'b00000000011000010010000000100011;
ROM[9561] <= 32'b00000000010000010000000100010011;
ROM[9562] <= 32'b00000001010000000000001110010011;
ROM[9563] <= 32'b00000000100000111000001110010011;
ROM[9564] <= 32'b01000000011100010000001110110011;
ROM[9565] <= 32'b00000000011100000000001000110011;
ROM[9566] <= 32'b00000000001000000000000110110011;
ROM[9567] <= 32'b01100011000000100000000011101111;
ROM[9568] <= 32'b00000111010000000000001110010011;
ROM[9569] <= 32'b00000000011100010010000000100011;
ROM[9570] <= 32'b00000000010000010000000100010011;
ROM[9571] <= 32'b00000000000000001001001110110111;
ROM[9572] <= 32'b01011101100000111000001110010011;
ROM[9573] <= 32'b00000000111000111000001110110011;
ROM[9574] <= 32'b00000000011100010010000000100011;
ROM[9575] <= 32'b00000000010000010000000100010011;
ROM[9576] <= 32'b00000000001100010010000000100011;
ROM[9577] <= 32'b00000000010000010000000100010011;
ROM[9578] <= 32'b00000000010000010010000000100011;
ROM[9579] <= 32'b00000000010000010000000100010011;
ROM[9580] <= 32'b00000000010100010010000000100011;
ROM[9581] <= 32'b00000000010000010000000100010011;
ROM[9582] <= 32'b00000000011000010010000000100011;
ROM[9583] <= 32'b00000000010000010000000100010011;
ROM[9584] <= 32'b00000001010000000000001110010011;
ROM[9585] <= 32'b00000000100000111000001110010011;
ROM[9586] <= 32'b01000000011100010000001110110011;
ROM[9587] <= 32'b00000000011100000000001000110011;
ROM[9588] <= 32'b00000000001000000000000110110011;
ROM[9589] <= 32'b01011101100000100000000011101111;
ROM[9590] <= 32'b00000111010100000000001110010011;
ROM[9591] <= 32'b00000000011100010010000000100011;
ROM[9592] <= 32'b00000000010000010000000100010011;
ROM[9593] <= 32'b00000000000000001001001110110111;
ROM[9594] <= 32'b01100011000000111000001110010011;
ROM[9595] <= 32'b00000000111000111000001110110011;
ROM[9596] <= 32'b00000000011100010010000000100011;
ROM[9597] <= 32'b00000000010000010000000100010011;
ROM[9598] <= 32'b00000000001100010010000000100011;
ROM[9599] <= 32'b00000000010000010000000100010011;
ROM[9600] <= 32'b00000000010000010010000000100011;
ROM[9601] <= 32'b00000000010000010000000100010011;
ROM[9602] <= 32'b00000000010100010010000000100011;
ROM[9603] <= 32'b00000000010000010000000100010011;
ROM[9604] <= 32'b00000000011000010010000000100011;
ROM[9605] <= 32'b00000000010000010000000100010011;
ROM[9606] <= 32'b00000001010000000000001110010011;
ROM[9607] <= 32'b00000000100000111000001110010011;
ROM[9608] <= 32'b01000000011100010000001110110011;
ROM[9609] <= 32'b00000000011100000000001000110011;
ROM[9610] <= 32'b00000000001000000000000110110011;
ROM[9611] <= 32'b01011000000000100000000011101111;
ROM[9612] <= 32'b00000110110000000000001110010011;
ROM[9613] <= 32'b00000000011100010010000000100011;
ROM[9614] <= 32'b00000000010000010000000100010011;
ROM[9615] <= 32'b00000000000000001001001110110111;
ROM[9616] <= 32'b01101000100000111000001110010011;
ROM[9617] <= 32'b00000000111000111000001110110011;
ROM[9618] <= 32'b00000000011100010010000000100011;
ROM[9619] <= 32'b00000000010000010000000100010011;
ROM[9620] <= 32'b00000000001100010010000000100011;
ROM[9621] <= 32'b00000000010000010000000100010011;
ROM[9622] <= 32'b00000000010000010010000000100011;
ROM[9623] <= 32'b00000000010000010000000100010011;
ROM[9624] <= 32'b00000000010100010010000000100011;
ROM[9625] <= 32'b00000000010000010000000100010011;
ROM[9626] <= 32'b00000000011000010010000000100011;
ROM[9627] <= 32'b00000000010000010000000100010011;
ROM[9628] <= 32'b00000001010000000000001110010011;
ROM[9629] <= 32'b00000000100000111000001110010011;
ROM[9630] <= 32'b01000000011100010000001110110011;
ROM[9631] <= 32'b00000000011100000000001000110011;
ROM[9632] <= 32'b00000000001000000000000110110011;
ROM[9633] <= 32'b01010010100000100000000011101111;
ROM[9634] <= 32'b00000110000100000000001110010011;
ROM[9635] <= 32'b00000000011100010010000000100011;
ROM[9636] <= 32'b00000000010000010000000100010011;
ROM[9637] <= 32'b00000000000000001001001110110111;
ROM[9638] <= 32'b01101110000000111000001110010011;
ROM[9639] <= 32'b00000000111000111000001110110011;
ROM[9640] <= 32'b00000000011100010010000000100011;
ROM[9641] <= 32'b00000000010000010000000100010011;
ROM[9642] <= 32'b00000000001100010010000000100011;
ROM[9643] <= 32'b00000000010000010000000100010011;
ROM[9644] <= 32'b00000000010000010010000000100011;
ROM[9645] <= 32'b00000000010000010000000100010011;
ROM[9646] <= 32'b00000000010100010010000000100011;
ROM[9647] <= 32'b00000000010000010000000100010011;
ROM[9648] <= 32'b00000000011000010010000000100011;
ROM[9649] <= 32'b00000000010000010000000100010011;
ROM[9650] <= 32'b00000001010000000000001110010011;
ROM[9651] <= 32'b00000000100000111000001110010011;
ROM[9652] <= 32'b01000000011100010000001110110011;
ROM[9653] <= 32'b00000000011100000000001000110011;
ROM[9654] <= 32'b00000000001000000000000110110011;
ROM[9655] <= 32'b01001101000000100000000011101111;
ROM[9656] <= 32'b00000111010000000000001110010011;
ROM[9657] <= 32'b00000000011100010010000000100011;
ROM[9658] <= 32'b00000000010000010000000100010011;
ROM[9659] <= 32'b00000000000000001001001110110111;
ROM[9660] <= 32'b01110011100000111000001110010011;
ROM[9661] <= 32'b00000000111000111000001110110011;
ROM[9662] <= 32'b00000000011100010010000000100011;
ROM[9663] <= 32'b00000000010000010000000100010011;
ROM[9664] <= 32'b00000000001100010010000000100011;
ROM[9665] <= 32'b00000000010000010000000100010011;
ROM[9666] <= 32'b00000000010000010010000000100011;
ROM[9667] <= 32'b00000000010000010000000100010011;
ROM[9668] <= 32'b00000000010100010010000000100011;
ROM[9669] <= 32'b00000000010000010000000100010011;
ROM[9670] <= 32'b00000000011000010010000000100011;
ROM[9671] <= 32'b00000000010000010000000100010011;
ROM[9672] <= 32'b00000001010000000000001110010011;
ROM[9673] <= 32'b00000000100000111000001110010011;
ROM[9674] <= 32'b01000000011100010000001110110011;
ROM[9675] <= 32'b00000000011100000000001000110011;
ROM[9676] <= 32'b00000000001000000000000110110011;
ROM[9677] <= 32'b01000111100000100000000011101111;
ROM[9678] <= 32'b00000110100100000000001110010011;
ROM[9679] <= 32'b00000000011100010010000000100011;
ROM[9680] <= 32'b00000000010000010000000100010011;
ROM[9681] <= 32'b00000000000000001001001110110111;
ROM[9682] <= 32'b01111001000000111000001110010011;
ROM[9683] <= 32'b00000000111000111000001110110011;
ROM[9684] <= 32'b00000000011100010010000000100011;
ROM[9685] <= 32'b00000000010000010000000100010011;
ROM[9686] <= 32'b00000000001100010010000000100011;
ROM[9687] <= 32'b00000000010000010000000100010011;
ROM[9688] <= 32'b00000000010000010010000000100011;
ROM[9689] <= 32'b00000000010000010000000100010011;
ROM[9690] <= 32'b00000000010100010010000000100011;
ROM[9691] <= 32'b00000000010000010000000100010011;
ROM[9692] <= 32'b00000000011000010010000000100011;
ROM[9693] <= 32'b00000000010000010000000100010011;
ROM[9694] <= 32'b00000001010000000000001110010011;
ROM[9695] <= 32'b00000000100000111000001110010011;
ROM[9696] <= 32'b01000000011100010000001110110011;
ROM[9697] <= 32'b00000000011100000000001000110011;
ROM[9698] <= 32'b00000000001000000000000110110011;
ROM[9699] <= 32'b01000010000000100000000011101111;
ROM[9700] <= 32'b00000110111100000000001110010011;
ROM[9701] <= 32'b00000000011100010010000000100011;
ROM[9702] <= 32'b00000000010000010000000100010011;
ROM[9703] <= 32'b00000000000000001001001110110111;
ROM[9704] <= 32'b01111110100000111000001110010011;
ROM[9705] <= 32'b00000000111000111000001110110011;
ROM[9706] <= 32'b00000000011100010010000000100011;
ROM[9707] <= 32'b00000000010000010000000100010011;
ROM[9708] <= 32'b00000000001100010010000000100011;
ROM[9709] <= 32'b00000000010000010000000100010011;
ROM[9710] <= 32'b00000000010000010010000000100011;
ROM[9711] <= 32'b00000000010000010000000100010011;
ROM[9712] <= 32'b00000000010100010010000000100011;
ROM[9713] <= 32'b00000000010000010000000100010011;
ROM[9714] <= 32'b00000000011000010010000000100011;
ROM[9715] <= 32'b00000000010000010000000100010011;
ROM[9716] <= 32'b00000001010000000000001110010011;
ROM[9717] <= 32'b00000000100000111000001110010011;
ROM[9718] <= 32'b01000000011100010000001110110011;
ROM[9719] <= 32'b00000000011100000000001000110011;
ROM[9720] <= 32'b00000000001000000000000110110011;
ROM[9721] <= 32'b00111100100000100000000011101111;
ROM[9722] <= 32'b00000110111000000000001110010011;
ROM[9723] <= 32'b00000000011100010010000000100011;
ROM[9724] <= 32'b00000000010000010000000100010011;
ROM[9725] <= 32'b00000000000000001010001110110111;
ROM[9726] <= 32'b10000100000000111000001110010011;
ROM[9727] <= 32'b00000000111000111000001110110011;
ROM[9728] <= 32'b00000000011100010010000000100011;
ROM[9729] <= 32'b00000000010000010000000100010011;
ROM[9730] <= 32'b00000000001100010010000000100011;
ROM[9731] <= 32'b00000000010000010000000100010011;
ROM[9732] <= 32'b00000000010000010010000000100011;
ROM[9733] <= 32'b00000000010000010000000100010011;
ROM[9734] <= 32'b00000000010100010010000000100011;
ROM[9735] <= 32'b00000000010000010000000100010011;
ROM[9736] <= 32'b00000000011000010010000000100011;
ROM[9737] <= 32'b00000000010000010000000100010011;
ROM[9738] <= 32'b00000001010000000000001110010011;
ROM[9739] <= 32'b00000000100000111000001110010011;
ROM[9740] <= 32'b01000000011100010000001110110011;
ROM[9741] <= 32'b00000000011100000000001000110011;
ROM[9742] <= 32'b00000000001000000000000110110011;
ROM[9743] <= 32'b00110111000000100000000011101111;
ROM[9744] <= 32'b00000111001100000000001110010011;
ROM[9745] <= 32'b00000000011100010010000000100011;
ROM[9746] <= 32'b00000000010000010000000100010011;
ROM[9747] <= 32'b00000000000000001010001110110111;
ROM[9748] <= 32'b10001001100000111000001110010011;
ROM[9749] <= 32'b00000000111000111000001110110011;
ROM[9750] <= 32'b00000000011100010010000000100011;
ROM[9751] <= 32'b00000000010000010000000100010011;
ROM[9752] <= 32'b00000000001100010010000000100011;
ROM[9753] <= 32'b00000000010000010000000100010011;
ROM[9754] <= 32'b00000000010000010010000000100011;
ROM[9755] <= 32'b00000000010000010000000100010011;
ROM[9756] <= 32'b00000000010100010010000000100011;
ROM[9757] <= 32'b00000000010000010000000100010011;
ROM[9758] <= 32'b00000000011000010010000000100011;
ROM[9759] <= 32'b00000000010000010000000100010011;
ROM[9760] <= 32'b00000001010000000000001110010011;
ROM[9761] <= 32'b00000000100000111000001110010011;
ROM[9762] <= 32'b01000000011100010000001110110011;
ROM[9763] <= 32'b00000000011100000000001000110011;
ROM[9764] <= 32'b00000000001000000000000110110011;
ROM[9765] <= 32'b00110001100000100000000011101111;
ROM[9766] <= 32'b00000010000000000000001110010011;
ROM[9767] <= 32'b00000000011100010010000000100011;
ROM[9768] <= 32'b00000000010000010000000100010011;
ROM[9769] <= 32'b00000000000000001010001110110111;
ROM[9770] <= 32'b10001111000000111000001110010011;
ROM[9771] <= 32'b00000000111000111000001110110011;
ROM[9772] <= 32'b00000000011100010010000000100011;
ROM[9773] <= 32'b00000000010000010000000100010011;
ROM[9774] <= 32'b00000000001100010010000000100011;
ROM[9775] <= 32'b00000000010000010000000100010011;
ROM[9776] <= 32'b00000000010000010010000000100011;
ROM[9777] <= 32'b00000000010000010000000100010011;
ROM[9778] <= 32'b00000000010100010010000000100011;
ROM[9779] <= 32'b00000000010000010000000100010011;
ROM[9780] <= 32'b00000000011000010010000000100011;
ROM[9781] <= 32'b00000000010000010000000100010011;
ROM[9782] <= 32'b00000001010000000000001110010011;
ROM[9783] <= 32'b00000000100000111000001110010011;
ROM[9784] <= 32'b01000000011100010000001110110011;
ROM[9785] <= 32'b00000000011100000000001000110011;
ROM[9786] <= 32'b00000000001000000000000110110011;
ROM[9787] <= 32'b00101100000000100000000011101111;
ROM[9788] <= 32'b00000111100100000000001110010011;
ROM[9789] <= 32'b00000000011100010010000000100011;
ROM[9790] <= 32'b00000000010000010000000100010011;
ROM[9791] <= 32'b00000000000000001010001110110111;
ROM[9792] <= 32'b10010100100000111000001110010011;
ROM[9793] <= 32'b00000000111000111000001110110011;
ROM[9794] <= 32'b00000000011100010010000000100011;
ROM[9795] <= 32'b00000000010000010000000100010011;
ROM[9796] <= 32'b00000000001100010010000000100011;
ROM[9797] <= 32'b00000000010000010000000100010011;
ROM[9798] <= 32'b00000000010000010010000000100011;
ROM[9799] <= 32'b00000000010000010000000100010011;
ROM[9800] <= 32'b00000000010100010010000000100011;
ROM[9801] <= 32'b00000000010000010000000100010011;
ROM[9802] <= 32'b00000000011000010010000000100011;
ROM[9803] <= 32'b00000000010000010000000100010011;
ROM[9804] <= 32'b00000001010000000000001110010011;
ROM[9805] <= 32'b00000000100000111000001110010011;
ROM[9806] <= 32'b01000000011100010000001110110011;
ROM[9807] <= 32'b00000000011100000000001000110011;
ROM[9808] <= 32'b00000000001000000000000110110011;
ROM[9809] <= 32'b00100110100000100000000011101111;
ROM[9810] <= 32'b00000110111100000000001110010011;
ROM[9811] <= 32'b00000000011100010010000000100011;
ROM[9812] <= 32'b00000000010000010000000100010011;
ROM[9813] <= 32'b00000000000000001010001110110111;
ROM[9814] <= 32'b10011010000000111000001110010011;
ROM[9815] <= 32'b00000000111000111000001110110011;
ROM[9816] <= 32'b00000000011100010010000000100011;
ROM[9817] <= 32'b00000000010000010000000100010011;
ROM[9818] <= 32'b00000000001100010010000000100011;
ROM[9819] <= 32'b00000000010000010000000100010011;
ROM[9820] <= 32'b00000000010000010010000000100011;
ROM[9821] <= 32'b00000000010000010000000100010011;
ROM[9822] <= 32'b00000000010100010010000000100011;
ROM[9823] <= 32'b00000000010000010000000100010011;
ROM[9824] <= 32'b00000000011000010010000000100011;
ROM[9825] <= 32'b00000000010000010000000100010011;
ROM[9826] <= 32'b00000001010000000000001110010011;
ROM[9827] <= 32'b00000000100000111000001110010011;
ROM[9828] <= 32'b01000000011100010000001110110011;
ROM[9829] <= 32'b00000000011100000000001000110011;
ROM[9830] <= 32'b00000000001000000000000110110011;
ROM[9831] <= 32'b00100001000000100000000011101111;
ROM[9832] <= 32'b00000111010100000000001110010011;
ROM[9833] <= 32'b00000000011100010010000000100011;
ROM[9834] <= 32'b00000000010000010000000100010011;
ROM[9835] <= 32'b00000000000000001010001110110111;
ROM[9836] <= 32'b10011111100000111000001110010011;
ROM[9837] <= 32'b00000000111000111000001110110011;
ROM[9838] <= 32'b00000000011100010010000000100011;
ROM[9839] <= 32'b00000000010000010000000100010011;
ROM[9840] <= 32'b00000000001100010010000000100011;
ROM[9841] <= 32'b00000000010000010000000100010011;
ROM[9842] <= 32'b00000000010000010010000000100011;
ROM[9843] <= 32'b00000000010000010000000100010011;
ROM[9844] <= 32'b00000000010100010010000000100011;
ROM[9845] <= 32'b00000000010000010000000100010011;
ROM[9846] <= 32'b00000000011000010010000000100011;
ROM[9847] <= 32'b00000000010000010000000100010011;
ROM[9848] <= 32'b00000001010000000000001110010011;
ROM[9849] <= 32'b00000000100000111000001110010011;
ROM[9850] <= 32'b01000000011100010000001110110011;
ROM[9851] <= 32'b00000000011100000000001000110011;
ROM[9852] <= 32'b00000000001000000000000110110011;
ROM[9853] <= 32'b00011011100000100000000011101111;
ROM[9854] <= 32'b00000010000000000000001110010011;
ROM[9855] <= 32'b00000000011100010010000000100011;
ROM[9856] <= 32'b00000000010000010000000100010011;
ROM[9857] <= 32'b00000000000000001010001110110111;
ROM[9858] <= 32'b10100101000000111000001110010011;
ROM[9859] <= 32'b00000000111000111000001110110011;
ROM[9860] <= 32'b00000000011100010010000000100011;
ROM[9861] <= 32'b00000000010000010000000100010011;
ROM[9862] <= 32'b00000000001100010010000000100011;
ROM[9863] <= 32'b00000000010000010000000100010011;
ROM[9864] <= 32'b00000000010000010010000000100011;
ROM[9865] <= 32'b00000000010000010000000100010011;
ROM[9866] <= 32'b00000000010100010010000000100011;
ROM[9867] <= 32'b00000000010000010000000100010011;
ROM[9868] <= 32'b00000000011000010010000000100011;
ROM[9869] <= 32'b00000000010000010000000100010011;
ROM[9870] <= 32'b00000001010000000000001110010011;
ROM[9871] <= 32'b00000000100000111000001110010011;
ROM[9872] <= 32'b01000000011100010000001110110011;
ROM[9873] <= 32'b00000000011100000000001000110011;
ROM[9874] <= 32'b00000000001000000000000110110011;
ROM[9875] <= 32'b00010110000000100000000011101111;
ROM[9876] <= 32'b00000110100000000000001110010011;
ROM[9877] <= 32'b00000000011100010010000000100011;
ROM[9878] <= 32'b00000000010000010000000100010011;
ROM[9879] <= 32'b00000000000000001010001110110111;
ROM[9880] <= 32'b10101010100000111000001110010011;
ROM[9881] <= 32'b00000000111000111000001110110011;
ROM[9882] <= 32'b00000000011100010010000000100011;
ROM[9883] <= 32'b00000000010000010000000100010011;
ROM[9884] <= 32'b00000000001100010010000000100011;
ROM[9885] <= 32'b00000000010000010000000100010011;
ROM[9886] <= 32'b00000000010000010010000000100011;
ROM[9887] <= 32'b00000000010000010000000100010011;
ROM[9888] <= 32'b00000000010100010010000000100011;
ROM[9889] <= 32'b00000000010000010000000100010011;
ROM[9890] <= 32'b00000000011000010010000000100011;
ROM[9891] <= 32'b00000000010000010000000100010011;
ROM[9892] <= 32'b00000001010000000000001110010011;
ROM[9893] <= 32'b00000000100000111000001110010011;
ROM[9894] <= 32'b01000000011100010000001110110011;
ROM[9895] <= 32'b00000000011100000000001000110011;
ROM[9896] <= 32'b00000000001000000000000110110011;
ROM[9897] <= 32'b00010000100000100000000011101111;
ROM[9898] <= 32'b00000110000100000000001110010011;
ROM[9899] <= 32'b00000000011100010010000000100011;
ROM[9900] <= 32'b00000000010000010000000100010011;
ROM[9901] <= 32'b00000000000000001010001110110111;
ROM[9902] <= 32'b10110000000000111000001110010011;
ROM[9903] <= 32'b00000000111000111000001110110011;
ROM[9904] <= 32'b00000000011100010010000000100011;
ROM[9905] <= 32'b00000000010000010000000100010011;
ROM[9906] <= 32'b00000000001100010010000000100011;
ROM[9907] <= 32'b00000000010000010000000100010011;
ROM[9908] <= 32'b00000000010000010010000000100011;
ROM[9909] <= 32'b00000000010000010000000100010011;
ROM[9910] <= 32'b00000000010100010010000000100011;
ROM[9911] <= 32'b00000000010000010000000100010011;
ROM[9912] <= 32'b00000000011000010010000000100011;
ROM[9913] <= 32'b00000000010000010000000100010011;
ROM[9914] <= 32'b00000001010000000000001110010011;
ROM[9915] <= 32'b00000000100000111000001110010011;
ROM[9916] <= 32'b01000000011100010000001110110011;
ROM[9917] <= 32'b00000000011100000000001000110011;
ROM[9918] <= 32'b00000000001000000000000110110011;
ROM[9919] <= 32'b00001011000000100000000011101111;
ROM[9920] <= 32'b00000111011000000000001110010011;
ROM[9921] <= 32'b00000000011100010010000000100011;
ROM[9922] <= 32'b00000000010000010000000100010011;
ROM[9923] <= 32'b00000000000000001010001110110111;
ROM[9924] <= 32'b10110101100000111000001110010011;
ROM[9925] <= 32'b00000000111000111000001110110011;
ROM[9926] <= 32'b00000000011100010010000000100011;
ROM[9927] <= 32'b00000000010000010000000100010011;
ROM[9928] <= 32'b00000000001100010010000000100011;
ROM[9929] <= 32'b00000000010000010000000100010011;
ROM[9930] <= 32'b00000000010000010010000000100011;
ROM[9931] <= 32'b00000000010000010000000100010011;
ROM[9932] <= 32'b00000000010100010010000000100011;
ROM[9933] <= 32'b00000000010000010000000100010011;
ROM[9934] <= 32'b00000000011000010010000000100011;
ROM[9935] <= 32'b00000000010000010000000100010011;
ROM[9936] <= 32'b00000001010000000000001110010011;
ROM[9937] <= 32'b00000000100000111000001110010011;
ROM[9938] <= 32'b01000000011100010000001110110011;
ROM[9939] <= 32'b00000000011100000000001000110011;
ROM[9940] <= 32'b00000000001000000000000110110011;
ROM[9941] <= 32'b00000101100000100000000011101111;
ROM[9942] <= 32'b00000110010100000000001110010011;
ROM[9943] <= 32'b00000000011100010010000000100011;
ROM[9944] <= 32'b00000000010000010000000100010011;
ROM[9945] <= 32'b00000000000000001010001110110111;
ROM[9946] <= 32'b10111011000000111000001110010011;
ROM[9947] <= 32'b00000000111000111000001110110011;
ROM[9948] <= 32'b00000000011100010010000000100011;
ROM[9949] <= 32'b00000000010000010000000100010011;
ROM[9950] <= 32'b00000000001100010010000000100011;
ROM[9951] <= 32'b00000000010000010000000100010011;
ROM[9952] <= 32'b00000000010000010010000000100011;
ROM[9953] <= 32'b00000000010000010000000100010011;
ROM[9954] <= 32'b00000000010100010010000000100011;
ROM[9955] <= 32'b00000000010000010000000100010011;
ROM[9956] <= 32'b00000000011000010010000000100011;
ROM[9957] <= 32'b00000000010000010000000100010011;
ROM[9958] <= 32'b00000001010000000000001110010011;
ROM[9959] <= 32'b00000000100000111000001110010011;
ROM[9960] <= 32'b01000000011100010000001110110011;
ROM[9961] <= 32'b00000000011100000000001000110011;
ROM[9962] <= 32'b00000000001000000000000110110011;
ROM[9963] <= 32'b00000000000000100000000011101111;
ROM[9964] <= 32'b00000010000000000000001110010011;
ROM[9965] <= 32'b00000000011100010010000000100011;
ROM[9966] <= 32'b00000000010000010000000100010011;
ROM[9967] <= 32'b00000000000000001010001110110111;
ROM[9968] <= 32'b11000000100000111000001110010011;
ROM[9969] <= 32'b00000000111000111000001110110011;
ROM[9970] <= 32'b00000000011100010010000000100011;
ROM[9971] <= 32'b00000000010000010000000100010011;
ROM[9972] <= 32'b00000000001100010010000000100011;
ROM[9973] <= 32'b00000000010000010000000100010011;
ROM[9974] <= 32'b00000000010000010010000000100011;
ROM[9975] <= 32'b00000000010000010000000100010011;
ROM[9976] <= 32'b00000000010100010010000000100011;
ROM[9977] <= 32'b00000000010000010000000100010011;
ROM[9978] <= 32'b00000000011000010010000000100011;
ROM[9979] <= 32'b00000000010000010000000100010011;
ROM[9980] <= 32'b00000001010000000000001110010011;
ROM[9981] <= 32'b00000000100000111000001110010011;
ROM[9982] <= 32'b01000000011100010000001110110011;
ROM[9983] <= 32'b00000000011100000000001000110011;
ROM[9984] <= 32'b00000000001000000000000110110011;
ROM[9985] <= 32'b01111010100100011111000011101111;
ROM[9986] <= 32'b00000111011100000000001110010011;
ROM[9987] <= 32'b00000000011100010010000000100011;
ROM[9988] <= 32'b00000000010000010000000100010011;
ROM[9989] <= 32'b00000000000000001010001110110111;
ROM[9990] <= 32'b11000110000000111000001110010011;
ROM[9991] <= 32'b00000000111000111000001110110011;
ROM[9992] <= 32'b00000000011100010010000000100011;
ROM[9993] <= 32'b00000000010000010000000100010011;
ROM[9994] <= 32'b00000000001100010010000000100011;
ROM[9995] <= 32'b00000000010000010000000100010011;
ROM[9996] <= 32'b00000000010000010010000000100011;
ROM[9997] <= 32'b00000000010000010000000100010011;
ROM[9998] <= 32'b00000000010100010010000000100011;
ROM[9999] <= 32'b00000000010000010000000100010011;
ROM[10000] <= 32'b00000000011000010010000000100011;
ROM[10001] <= 32'b00000000010000010000000100010011;
ROM[10002] <= 32'b00000001010000000000001110010011;
ROM[10003] <= 32'b00000000100000111000001110010011;
ROM[10004] <= 32'b01000000011100010000001110110011;
ROM[10005] <= 32'b00000000011100000000001000110011;
ROM[10006] <= 32'b00000000001000000000000110110011;
ROM[10007] <= 32'b01110101000100011111000011101111;
ROM[10008] <= 32'b00000110111100000000001110010011;
ROM[10009] <= 32'b00000000011100010010000000100011;
ROM[10010] <= 32'b00000000010000010000000100010011;
ROM[10011] <= 32'b00000000000000001010001110110111;
ROM[10012] <= 32'b11001011100000111000001110010011;
ROM[10013] <= 32'b00000000111000111000001110110011;
ROM[10014] <= 32'b00000000011100010010000000100011;
ROM[10015] <= 32'b00000000010000010000000100010011;
ROM[10016] <= 32'b00000000001100010010000000100011;
ROM[10017] <= 32'b00000000010000010000000100010011;
ROM[10018] <= 32'b00000000010000010010000000100011;
ROM[10019] <= 32'b00000000010000010000000100010011;
ROM[10020] <= 32'b00000000010100010010000000100011;
ROM[10021] <= 32'b00000000010000010000000100010011;
ROM[10022] <= 32'b00000000011000010010000000100011;
ROM[10023] <= 32'b00000000010000010000000100010011;
ROM[10024] <= 32'b00000001010000000000001110010011;
ROM[10025] <= 32'b00000000100000111000001110010011;
ROM[10026] <= 32'b01000000011100010000001110110011;
ROM[10027] <= 32'b00000000011100000000001000110011;
ROM[10028] <= 32'b00000000001000000000000110110011;
ROM[10029] <= 32'b01101111100100011111000011101111;
ROM[10030] <= 32'b00000110111000000000001110010011;
ROM[10031] <= 32'b00000000011100010010000000100011;
ROM[10032] <= 32'b00000000010000010000000100010011;
ROM[10033] <= 32'b00000000000000001010001110110111;
ROM[10034] <= 32'b11010001000000111000001110010011;
ROM[10035] <= 32'b00000000111000111000001110110011;
ROM[10036] <= 32'b00000000011100010010000000100011;
ROM[10037] <= 32'b00000000010000010000000100010011;
ROM[10038] <= 32'b00000000001100010010000000100011;
ROM[10039] <= 32'b00000000010000010000000100010011;
ROM[10040] <= 32'b00000000010000010010000000100011;
ROM[10041] <= 32'b00000000010000010000000100010011;
ROM[10042] <= 32'b00000000010100010010000000100011;
ROM[10043] <= 32'b00000000010000010000000100010011;
ROM[10044] <= 32'b00000000011000010010000000100011;
ROM[10045] <= 32'b00000000010000010000000100010011;
ROM[10046] <= 32'b00000001010000000000001110010011;
ROM[10047] <= 32'b00000000100000111000001110010011;
ROM[10048] <= 32'b01000000011100010000001110110011;
ROM[10049] <= 32'b00000000011100000000001000110011;
ROM[10050] <= 32'b00000000001000000000000110110011;
ROM[10051] <= 32'b01101010000100011111000011101111;
ROM[10052] <= 32'b00000010000000000000001110010011;
ROM[10053] <= 32'b00000000011100010010000000100011;
ROM[10054] <= 32'b00000000010000010000000100010011;
ROM[10055] <= 32'b00000000000000001010001110110111;
ROM[10056] <= 32'b11010110100000111000001110010011;
ROM[10057] <= 32'b00000000111000111000001110110011;
ROM[10058] <= 32'b00000000011100010010000000100011;
ROM[10059] <= 32'b00000000010000010000000100010011;
ROM[10060] <= 32'b00000000001100010010000000100011;
ROM[10061] <= 32'b00000000010000010000000100010011;
ROM[10062] <= 32'b00000000010000010010000000100011;
ROM[10063] <= 32'b00000000010000010000000100010011;
ROM[10064] <= 32'b00000000010100010010000000100011;
ROM[10065] <= 32'b00000000010000010000000100010011;
ROM[10066] <= 32'b00000000011000010010000000100011;
ROM[10067] <= 32'b00000000010000010000000100010011;
ROM[10068] <= 32'b00000001010000000000001110010011;
ROM[10069] <= 32'b00000000100000111000001110010011;
ROM[10070] <= 32'b01000000011100010000001110110011;
ROM[10071] <= 32'b00000000011100000000001000110011;
ROM[10072] <= 32'b00000000001000000000000110110011;
ROM[10073] <= 32'b01100100100100011111000011101111;
ROM[10074] <= 32'b00000111010000000000001110010011;
ROM[10075] <= 32'b00000000011100010010000000100011;
ROM[10076] <= 32'b00000000010000010000000100010011;
ROM[10077] <= 32'b00000000000000001010001110110111;
ROM[10078] <= 32'b11011100000000111000001110010011;
ROM[10079] <= 32'b00000000111000111000001110110011;
ROM[10080] <= 32'b00000000011100010010000000100011;
ROM[10081] <= 32'b00000000010000010000000100010011;
ROM[10082] <= 32'b00000000001100010010000000100011;
ROM[10083] <= 32'b00000000010000010000000100010011;
ROM[10084] <= 32'b00000000010000010010000000100011;
ROM[10085] <= 32'b00000000010000010000000100010011;
ROM[10086] <= 32'b00000000010100010010000000100011;
ROM[10087] <= 32'b00000000010000010000000100010011;
ROM[10088] <= 32'b00000000011000010010000000100011;
ROM[10089] <= 32'b00000000010000010000000100010011;
ROM[10090] <= 32'b00000001010000000000001110010011;
ROM[10091] <= 32'b00000000100000111000001110010011;
ROM[10092] <= 32'b01000000011100010000001110110011;
ROM[10093] <= 32'b00000000011100000000001000110011;
ROM[10094] <= 32'b00000000001000000000000110110011;
ROM[10095] <= 32'b01011111000100011111000011101111;
ROM[10096] <= 32'b00000110100000000000001110010011;
ROM[10097] <= 32'b00000000011100010010000000100011;
ROM[10098] <= 32'b00000000010000010000000100010011;
ROM[10099] <= 32'b00000000000000001010001110110111;
ROM[10100] <= 32'b11100001100000111000001110010011;
ROM[10101] <= 32'b00000000111000111000001110110011;
ROM[10102] <= 32'b00000000011100010010000000100011;
ROM[10103] <= 32'b00000000010000010000000100010011;
ROM[10104] <= 32'b00000000001100010010000000100011;
ROM[10105] <= 32'b00000000010000010000000100010011;
ROM[10106] <= 32'b00000000010000010010000000100011;
ROM[10107] <= 32'b00000000010000010000000100010011;
ROM[10108] <= 32'b00000000010100010010000000100011;
ROM[10109] <= 32'b00000000010000010000000100010011;
ROM[10110] <= 32'b00000000011000010010000000100011;
ROM[10111] <= 32'b00000000010000010000000100010011;
ROM[10112] <= 32'b00000001010000000000001110010011;
ROM[10113] <= 32'b00000000100000111000001110010011;
ROM[10114] <= 32'b01000000011100010000001110110011;
ROM[10115] <= 32'b00000000011100000000001000110011;
ROM[10116] <= 32'b00000000001000000000000110110011;
ROM[10117] <= 32'b01011001100100011111000011101111;
ROM[10118] <= 32'b00000110010100000000001110010011;
ROM[10119] <= 32'b00000000011100010010000000100011;
ROM[10120] <= 32'b00000000010000010000000100010011;
ROM[10121] <= 32'b00000000000000001010001110110111;
ROM[10122] <= 32'b11100111000000111000001110010011;
ROM[10123] <= 32'b00000000111000111000001110110011;
ROM[10124] <= 32'b00000000011100010010000000100011;
ROM[10125] <= 32'b00000000010000010000000100010011;
ROM[10126] <= 32'b00000000001100010010000000100011;
ROM[10127] <= 32'b00000000010000010000000100010011;
ROM[10128] <= 32'b00000000010000010010000000100011;
ROM[10129] <= 32'b00000000010000010000000100010011;
ROM[10130] <= 32'b00000000010100010010000000100011;
ROM[10131] <= 32'b00000000010000010000000100010011;
ROM[10132] <= 32'b00000000011000010010000000100011;
ROM[10133] <= 32'b00000000010000010000000100010011;
ROM[10134] <= 32'b00000001010000000000001110010011;
ROM[10135] <= 32'b00000000100000111000001110010011;
ROM[10136] <= 32'b01000000011100010000001110110011;
ROM[10137] <= 32'b00000000011100000000001000110011;
ROM[10138] <= 32'b00000000001000000000000110110011;
ROM[10139] <= 32'b01010100000100011111000011101111;
ROM[10140] <= 32'b00000010000000000000001110010011;
ROM[10141] <= 32'b00000000011100010010000000100011;
ROM[10142] <= 32'b00000000010000010000000100010011;
ROM[10143] <= 32'b00000000000000001010001110110111;
ROM[10144] <= 32'b11101100100000111000001110010011;
ROM[10145] <= 32'b00000000111000111000001110110011;
ROM[10146] <= 32'b00000000011100010010000000100011;
ROM[10147] <= 32'b00000000010000010000000100010011;
ROM[10148] <= 32'b00000000001100010010000000100011;
ROM[10149] <= 32'b00000000010000010000000100010011;
ROM[10150] <= 32'b00000000010000010010000000100011;
ROM[10151] <= 32'b00000000010000010000000100010011;
ROM[10152] <= 32'b00000000010100010010000000100011;
ROM[10153] <= 32'b00000000010000010000000100010011;
ROM[10154] <= 32'b00000000011000010010000000100011;
ROM[10155] <= 32'b00000000010000010000000100010011;
ROM[10156] <= 32'b00000001010000000000001110010011;
ROM[10157] <= 32'b00000000100000111000001110010011;
ROM[10158] <= 32'b01000000011100010000001110110011;
ROM[10159] <= 32'b00000000011100000000001000110011;
ROM[10160] <= 32'b00000000001000000000000110110011;
ROM[10161] <= 32'b01001110100100011111000011101111;
ROM[10162] <= 32'b00000110011100000000001110010011;
ROM[10163] <= 32'b00000000011100010010000000100011;
ROM[10164] <= 32'b00000000010000010000000100010011;
ROM[10165] <= 32'b00000000000000001010001110110111;
ROM[10166] <= 32'b11110010000000111000001110010011;
ROM[10167] <= 32'b00000000111000111000001110110011;
ROM[10168] <= 32'b00000000011100010010000000100011;
ROM[10169] <= 32'b00000000010000010000000100010011;
ROM[10170] <= 32'b00000000001100010010000000100011;
ROM[10171] <= 32'b00000000010000010000000100010011;
ROM[10172] <= 32'b00000000010000010010000000100011;
ROM[10173] <= 32'b00000000010000010000000100010011;
ROM[10174] <= 32'b00000000010100010010000000100011;
ROM[10175] <= 32'b00000000010000010000000100010011;
ROM[10176] <= 32'b00000000011000010010000000100011;
ROM[10177] <= 32'b00000000010000010000000100010011;
ROM[10178] <= 32'b00000001010000000000001110010011;
ROM[10179] <= 32'b00000000100000111000001110010011;
ROM[10180] <= 32'b01000000011100010000001110110011;
ROM[10181] <= 32'b00000000011100000000001000110011;
ROM[10182] <= 32'b00000000001000000000000110110011;
ROM[10183] <= 32'b01001001000100011111000011101111;
ROM[10184] <= 32'b00000110000100000000001110010011;
ROM[10185] <= 32'b00000000011100010010000000100011;
ROM[10186] <= 32'b00000000010000010000000100010011;
ROM[10187] <= 32'b00000000000000001010001110110111;
ROM[10188] <= 32'b11110111100000111000001110010011;
ROM[10189] <= 32'b00000000111000111000001110110011;
ROM[10190] <= 32'b00000000011100010010000000100011;
ROM[10191] <= 32'b00000000010000010000000100010011;
ROM[10192] <= 32'b00000000001100010010000000100011;
ROM[10193] <= 32'b00000000010000010000000100010011;
ROM[10194] <= 32'b00000000010000010010000000100011;
ROM[10195] <= 32'b00000000010000010000000100010011;
ROM[10196] <= 32'b00000000010100010010000000100011;
ROM[10197] <= 32'b00000000010000010000000100010011;
ROM[10198] <= 32'b00000000011000010010000000100011;
ROM[10199] <= 32'b00000000010000010000000100010011;
ROM[10200] <= 32'b00000001010000000000001110010011;
ROM[10201] <= 32'b00000000100000111000001110010011;
ROM[10202] <= 32'b01000000011100010000001110110011;
ROM[10203] <= 32'b00000000011100000000001000110011;
ROM[10204] <= 32'b00000000001000000000000110110011;
ROM[10205] <= 32'b01000011100100011111000011101111;
ROM[10206] <= 32'b00000110110100000000001110010011;
ROM[10207] <= 32'b00000000011100010010000000100011;
ROM[10208] <= 32'b00000000010000010000000100010011;
ROM[10209] <= 32'b00000000000000001010001110110111;
ROM[10210] <= 32'b11111101000000111000001110010011;
ROM[10211] <= 32'b00000000111000111000001110110011;
ROM[10212] <= 32'b00000000011100010010000000100011;
ROM[10213] <= 32'b00000000010000010000000100010011;
ROM[10214] <= 32'b00000000001100010010000000100011;
ROM[10215] <= 32'b00000000010000010000000100010011;
ROM[10216] <= 32'b00000000010000010010000000100011;
ROM[10217] <= 32'b00000000010000010000000100010011;
ROM[10218] <= 32'b00000000010100010010000000100011;
ROM[10219] <= 32'b00000000010000010000000100010011;
ROM[10220] <= 32'b00000000011000010010000000100011;
ROM[10221] <= 32'b00000000010000010000000100010011;
ROM[10222] <= 32'b00000001010000000000001110010011;
ROM[10223] <= 32'b00000000100000111000001110010011;
ROM[10224] <= 32'b01000000011100010000001110110011;
ROM[10225] <= 32'b00000000011100000000001000110011;
ROM[10226] <= 32'b00000000001000000000000110110011;
ROM[10227] <= 32'b00111110000100011111000011101111;
ROM[10228] <= 32'b00000110010100000000001110010011;
ROM[10229] <= 32'b00000000011100010010000000100011;
ROM[10230] <= 32'b00000000010000010000000100010011;
ROM[10231] <= 32'b00000000000000001010001110110111;
ROM[10232] <= 32'b00000010100000111000001110010011;
ROM[10233] <= 32'b00000000111000111000001110110011;
ROM[10234] <= 32'b00000000011100010010000000100011;
ROM[10235] <= 32'b00000000010000010000000100010011;
ROM[10236] <= 32'b00000000001100010010000000100011;
ROM[10237] <= 32'b00000000010000010000000100010011;
ROM[10238] <= 32'b00000000010000010010000000100011;
ROM[10239] <= 32'b00000000010000010000000100010011;
ROM[10240] <= 32'b00000000010100010010000000100011;
ROM[10241] <= 32'b00000000010000010000000100010011;
ROM[10242] <= 32'b00000000011000010010000000100011;
ROM[10243] <= 32'b00000000010000010000000100010011;
ROM[10244] <= 32'b00000001010000000000001110010011;
ROM[10245] <= 32'b00000000100000111000001110010011;
ROM[10246] <= 32'b01000000011100010000001110110011;
ROM[10247] <= 32'b00000000011100000000001000110011;
ROM[10248] <= 32'b00000000001000000000000110110011;
ROM[10249] <= 32'b00111000100100011111000011101111;
ROM[10250] <= 32'b00000010000100000000001110010011;
ROM[10251] <= 32'b00000000011100010010000000100011;
ROM[10252] <= 32'b00000000010000010000000100010011;
ROM[10253] <= 32'b00000000000000001010001110110111;
ROM[10254] <= 32'b00001000000000111000001110010011;
ROM[10255] <= 32'b00000000111000111000001110110011;
ROM[10256] <= 32'b00000000011100010010000000100011;
ROM[10257] <= 32'b00000000010000010000000100010011;
ROM[10258] <= 32'b00000000001100010010000000100011;
ROM[10259] <= 32'b00000000010000010000000100010011;
ROM[10260] <= 32'b00000000010000010010000000100011;
ROM[10261] <= 32'b00000000010000010000000100010011;
ROM[10262] <= 32'b00000000010100010010000000100011;
ROM[10263] <= 32'b00000000010000010000000100010011;
ROM[10264] <= 32'b00000000011000010010000000100011;
ROM[10265] <= 32'b00000000010000010000000100010011;
ROM[10266] <= 32'b00000001010000000000001110010011;
ROM[10267] <= 32'b00000000100000111000001110010011;
ROM[10268] <= 32'b01000000011100010000001110110011;
ROM[10269] <= 32'b00000000011100000000001000110011;
ROM[10270] <= 32'b00000000001000000000000110110011;
ROM[10271] <= 32'b00110011000100011111000011101111;
ROM[10272] <= 32'b00000000000000001010001110110111;
ROM[10273] <= 32'b00001100110000111000001110010011;
ROM[10274] <= 32'b00000000111000111000001110110011;
ROM[10275] <= 32'b00000000011100010010000000100011;
ROM[10276] <= 32'b00000000010000010000000100010011;
ROM[10277] <= 32'b00000000001100010010000000100011;
ROM[10278] <= 32'b00000000010000010000000100010011;
ROM[10279] <= 32'b00000000010000010010000000100011;
ROM[10280] <= 32'b00000000010000010000000100010011;
ROM[10281] <= 32'b00000000010100010010000000100011;
ROM[10282] <= 32'b00000000010000010000000100010011;
ROM[10283] <= 32'b00000000011000010010000000100011;
ROM[10284] <= 32'b00000000010000010000000100010011;
ROM[10285] <= 32'b00000001010000000000001110010011;
ROM[10286] <= 32'b00000000010000111000001110010011;
ROM[10287] <= 32'b01000000011100010000001110110011;
ROM[10288] <= 32'b00000000011100000000001000110011;
ROM[10289] <= 32'b00000000001000000000000110110011;
ROM[10290] <= 32'b01101010000100001100000011101111;
ROM[10291] <= 32'b11111111110000010000000100010011;
ROM[10292] <= 32'b00000000000000010010001110000011;
ROM[10293] <= 32'b00000000011101100010000000100011;
ROM[10294] <= 32'b00000000000000001010001110110111;
ROM[10295] <= 32'b00010010010000111000001110010011;
ROM[10296] <= 32'b00000000111000111000001110110011;
ROM[10297] <= 32'b00000000011100010010000000100011;
ROM[10298] <= 32'b00000000010000010000000100010011;
ROM[10299] <= 32'b00000000001100010010000000100011;
ROM[10300] <= 32'b00000000010000010000000100010011;
ROM[10301] <= 32'b00000000010000010010000000100011;
ROM[10302] <= 32'b00000000010000010000000100010011;
ROM[10303] <= 32'b00000000010100010010000000100011;
ROM[10304] <= 32'b00000000010000010000000100010011;
ROM[10305] <= 32'b00000000011000010010000000100011;
ROM[10306] <= 32'b00000000010000010000000100010011;
ROM[10307] <= 32'b00000001010000000000001110010011;
ROM[10308] <= 32'b00000000000000111000001110010011;
ROM[10309] <= 32'b01000000011100010000001110110011;
ROM[10310] <= 32'b00000000011100000000001000110011;
ROM[10311] <= 32'b00000000001000000000000110110011;
ROM[10312] <= 32'b00100100100000001101000011101111;
ROM[10313] <= 32'b11111111110000010000000100010011;
ROM[10314] <= 32'b00000000000000010010001110000011;
ROM[10315] <= 32'b00000000011101100010000000100011;
ROM[10316] <= 32'b00000000110000000000001110010011;
ROM[10317] <= 32'b00000000011100010010000000100011;
ROM[10318] <= 32'b00000000010000010000000100010011;
ROM[10319] <= 32'b00000000000000001010001110110111;
ROM[10320] <= 32'b00011000100000111000001110010011;
ROM[10321] <= 32'b00000000111000111000001110110011;
ROM[10322] <= 32'b00000000011100010010000000100011;
ROM[10323] <= 32'b00000000010000010000000100010011;
ROM[10324] <= 32'b00000000001100010010000000100011;
ROM[10325] <= 32'b00000000010000010000000100010011;
ROM[10326] <= 32'b00000000010000010010000000100011;
ROM[10327] <= 32'b00000000010000010000000100010011;
ROM[10328] <= 32'b00000000010100010010000000100011;
ROM[10329] <= 32'b00000000010000010000000100010011;
ROM[10330] <= 32'b00000000011000010010000000100011;
ROM[10331] <= 32'b00000000010000010000000100010011;
ROM[10332] <= 32'b00000001010000000000001110010011;
ROM[10333] <= 32'b00000000010000111000001110010011;
ROM[10334] <= 32'b01000000011100010000001110110011;
ROM[10335] <= 32'b00000000011100000000001000110011;
ROM[10336] <= 32'b00000000001000000000000110110011;
ROM[10337] <= 32'b01011011100000011111000011101111;
ROM[10338] <= 32'b00000101010000000000001110010011;
ROM[10339] <= 32'b00000000011100010010000000100011;
ROM[10340] <= 32'b00000000010000010000000100010011;
ROM[10341] <= 32'b00000000000000001010001110110111;
ROM[10342] <= 32'b00011110000000111000001110010011;
ROM[10343] <= 32'b00000000111000111000001110110011;
ROM[10344] <= 32'b00000000011100010010000000100011;
ROM[10345] <= 32'b00000000010000010000000100010011;
ROM[10346] <= 32'b00000000001100010010000000100011;
ROM[10347] <= 32'b00000000010000010000000100010011;
ROM[10348] <= 32'b00000000010000010010000000100011;
ROM[10349] <= 32'b00000000010000010000000100010011;
ROM[10350] <= 32'b00000000010100010010000000100011;
ROM[10351] <= 32'b00000000010000010000000100010011;
ROM[10352] <= 32'b00000000011000010010000000100011;
ROM[10353] <= 32'b00000000010000010000000100010011;
ROM[10354] <= 32'b00000001010000000000001110010011;
ROM[10355] <= 32'b00000000100000111000001110010011;
ROM[10356] <= 32'b01000000011100010000001110110011;
ROM[10357] <= 32'b00000000011100000000001000110011;
ROM[10358] <= 32'b00000000001000000000000110110011;
ROM[10359] <= 32'b00011101000100011111000011101111;
ROM[10360] <= 32'b00000110100000000000001110010011;
ROM[10361] <= 32'b00000000011100010010000000100011;
ROM[10362] <= 32'b00000000010000010000000100010011;
ROM[10363] <= 32'b00000000000000001010001110110111;
ROM[10364] <= 32'b00100011100000111000001110010011;
ROM[10365] <= 32'b00000000111000111000001110110011;
ROM[10366] <= 32'b00000000011100010010000000100011;
ROM[10367] <= 32'b00000000010000010000000100010011;
ROM[10368] <= 32'b00000000001100010010000000100011;
ROM[10369] <= 32'b00000000010000010000000100010011;
ROM[10370] <= 32'b00000000010000010010000000100011;
ROM[10371] <= 32'b00000000010000010000000100010011;
ROM[10372] <= 32'b00000000010100010010000000100011;
ROM[10373] <= 32'b00000000010000010000000100010011;
ROM[10374] <= 32'b00000000011000010010000000100011;
ROM[10375] <= 32'b00000000010000010000000100010011;
ROM[10376] <= 32'b00000001010000000000001110010011;
ROM[10377] <= 32'b00000000100000111000001110010011;
ROM[10378] <= 32'b01000000011100010000001110110011;
ROM[10379] <= 32'b00000000011100000000001000110011;
ROM[10380] <= 32'b00000000001000000000000110110011;
ROM[10381] <= 32'b00010111100100011111000011101111;
ROM[10382] <= 32'b00000110010100000000001110010011;
ROM[10383] <= 32'b00000000011100010010000000100011;
ROM[10384] <= 32'b00000000010000010000000100010011;
ROM[10385] <= 32'b00000000000000001010001110110111;
ROM[10386] <= 32'b00101001000000111000001110010011;
ROM[10387] <= 32'b00000000111000111000001110110011;
ROM[10388] <= 32'b00000000011100010010000000100011;
ROM[10389] <= 32'b00000000010000010000000100010011;
ROM[10390] <= 32'b00000000001100010010000000100011;
ROM[10391] <= 32'b00000000010000010000000100010011;
ROM[10392] <= 32'b00000000010000010010000000100011;
ROM[10393] <= 32'b00000000010000010000000100010011;
ROM[10394] <= 32'b00000000010100010010000000100011;
ROM[10395] <= 32'b00000000010000010000000100010011;
ROM[10396] <= 32'b00000000011000010010000000100011;
ROM[10397] <= 32'b00000000010000010000000100010011;
ROM[10398] <= 32'b00000001010000000000001110010011;
ROM[10399] <= 32'b00000000100000111000001110010011;
ROM[10400] <= 32'b01000000011100010000001110110011;
ROM[10401] <= 32'b00000000011100000000001000110011;
ROM[10402] <= 32'b00000000001000000000000110110011;
ROM[10403] <= 32'b00010010000100011111000011101111;
ROM[10404] <= 32'b00000010000000000000001110010011;
ROM[10405] <= 32'b00000000011100010010000000100011;
ROM[10406] <= 32'b00000000010000010000000100010011;
ROM[10407] <= 32'b00000000000000001010001110110111;
ROM[10408] <= 32'b00101110100000111000001110010011;
ROM[10409] <= 32'b00000000111000111000001110110011;
ROM[10410] <= 32'b00000000011100010010000000100011;
ROM[10411] <= 32'b00000000010000010000000100010011;
ROM[10412] <= 32'b00000000001100010010000000100011;
ROM[10413] <= 32'b00000000010000010000000100010011;
ROM[10414] <= 32'b00000000010000010010000000100011;
ROM[10415] <= 32'b00000000010000010000000100010011;
ROM[10416] <= 32'b00000000010100010010000000100011;
ROM[10417] <= 32'b00000000010000010000000100010011;
ROM[10418] <= 32'b00000000011000010010000000100011;
ROM[10419] <= 32'b00000000010000010000000100010011;
ROM[10420] <= 32'b00000001010000000000001110010011;
ROM[10421] <= 32'b00000000100000111000001110010011;
ROM[10422] <= 32'b01000000011100010000001110110011;
ROM[10423] <= 32'b00000000011100000000001000110011;
ROM[10424] <= 32'b00000000001000000000000110110011;
ROM[10425] <= 32'b00001100100100011111000011101111;
ROM[10426] <= 32'b00000111011100000000001110010011;
ROM[10427] <= 32'b00000000011100010010000000100011;
ROM[10428] <= 32'b00000000010000010000000100010011;
ROM[10429] <= 32'b00000000000000001010001110110111;
ROM[10430] <= 32'b00110100000000111000001110010011;
ROM[10431] <= 32'b00000000111000111000001110110011;
ROM[10432] <= 32'b00000000011100010010000000100011;
ROM[10433] <= 32'b00000000010000010000000100010011;
ROM[10434] <= 32'b00000000001100010010000000100011;
ROM[10435] <= 32'b00000000010000010000000100010011;
ROM[10436] <= 32'b00000000010000010010000000100011;
ROM[10437] <= 32'b00000000010000010000000100010011;
ROM[10438] <= 32'b00000000010100010010000000100011;
ROM[10439] <= 32'b00000000010000010000000100010011;
ROM[10440] <= 32'b00000000011000010010000000100011;
ROM[10441] <= 32'b00000000010000010000000100010011;
ROM[10442] <= 32'b00000001010000000000001110010011;
ROM[10443] <= 32'b00000000100000111000001110010011;
ROM[10444] <= 32'b01000000011100010000001110110011;
ROM[10445] <= 32'b00000000011100000000001000110011;
ROM[10446] <= 32'b00000000001000000000000110110011;
ROM[10447] <= 32'b00000111000100011111000011101111;
ROM[10448] <= 32'b00000110111100000000001110010011;
ROM[10449] <= 32'b00000000011100010010000000100011;
ROM[10450] <= 32'b00000000010000010000000100010011;
ROM[10451] <= 32'b00000000000000001010001110110111;
ROM[10452] <= 32'b00111001100000111000001110010011;
ROM[10453] <= 32'b00000000111000111000001110110011;
ROM[10454] <= 32'b00000000011100010010000000100011;
ROM[10455] <= 32'b00000000010000010000000100010011;
ROM[10456] <= 32'b00000000001100010010000000100011;
ROM[10457] <= 32'b00000000010000010000000100010011;
ROM[10458] <= 32'b00000000010000010010000000100011;
ROM[10459] <= 32'b00000000010000010000000100010011;
ROM[10460] <= 32'b00000000010100010010000000100011;
ROM[10461] <= 32'b00000000010000010000000100010011;
ROM[10462] <= 32'b00000000011000010010000000100011;
ROM[10463] <= 32'b00000000010000010000000100010011;
ROM[10464] <= 32'b00000001010000000000001110010011;
ROM[10465] <= 32'b00000000100000111000001110010011;
ROM[10466] <= 32'b01000000011100010000001110110011;
ROM[10467] <= 32'b00000000011100000000001000110011;
ROM[10468] <= 32'b00000000001000000000000110110011;
ROM[10469] <= 32'b00000001100100011111000011101111;
ROM[10470] <= 32'b00000111001000000000001110010011;
ROM[10471] <= 32'b00000000011100010010000000100011;
ROM[10472] <= 32'b00000000010000010000000100010011;
ROM[10473] <= 32'b00000000000000001010001110110111;
ROM[10474] <= 32'b00111111000000111000001110010011;
ROM[10475] <= 32'b00000000111000111000001110110011;
ROM[10476] <= 32'b00000000011100010010000000100011;
ROM[10477] <= 32'b00000000010000010000000100010011;
ROM[10478] <= 32'b00000000001100010010000000100011;
ROM[10479] <= 32'b00000000010000010000000100010011;
ROM[10480] <= 32'b00000000010000010010000000100011;
ROM[10481] <= 32'b00000000010000010000000100010011;
ROM[10482] <= 32'b00000000010100010010000000100011;
ROM[10483] <= 32'b00000000010000010000000100010011;
ROM[10484] <= 32'b00000000011000010010000000100011;
ROM[10485] <= 32'b00000000010000010000000100010011;
ROM[10486] <= 32'b00000001010000000000001110010011;
ROM[10487] <= 32'b00000000100000111000001110010011;
ROM[10488] <= 32'b01000000011100010000001110110011;
ROM[10489] <= 32'b00000000011100000000001000110011;
ROM[10490] <= 32'b00000000001000000000000110110011;
ROM[10491] <= 32'b01111100000000011111000011101111;
ROM[10492] <= 32'b00000110010000000000001110010011;
ROM[10493] <= 32'b00000000011100010010000000100011;
ROM[10494] <= 32'b00000000010000010000000100010011;
ROM[10495] <= 32'b00000000000000001010001110110111;
ROM[10496] <= 32'b01000100100000111000001110010011;
ROM[10497] <= 32'b00000000111000111000001110110011;
ROM[10498] <= 32'b00000000011100010010000000100011;
ROM[10499] <= 32'b00000000010000010000000100010011;
ROM[10500] <= 32'b00000000001100010010000000100011;
ROM[10501] <= 32'b00000000010000010000000100010011;
ROM[10502] <= 32'b00000000010000010010000000100011;
ROM[10503] <= 32'b00000000010000010000000100010011;
ROM[10504] <= 32'b00000000010100010010000000100011;
ROM[10505] <= 32'b00000000010000010000000100010011;
ROM[10506] <= 32'b00000000011000010010000000100011;
ROM[10507] <= 32'b00000000010000010000000100010011;
ROM[10508] <= 32'b00000001010000000000001110010011;
ROM[10509] <= 32'b00000000100000111000001110010011;
ROM[10510] <= 32'b01000000011100010000001110110011;
ROM[10511] <= 32'b00000000011100000000001000110011;
ROM[10512] <= 32'b00000000001000000000000110110011;
ROM[10513] <= 32'b01110110100000011111000011101111;
ROM[10514] <= 32'b00000010000000000000001110010011;
ROM[10515] <= 32'b00000000011100010010000000100011;
ROM[10516] <= 32'b00000000010000010000000100010011;
ROM[10517] <= 32'b00000000000000001010001110110111;
ROM[10518] <= 32'b01001010000000111000001110010011;
ROM[10519] <= 32'b00000000111000111000001110110011;
ROM[10520] <= 32'b00000000011100010010000000100011;
ROM[10521] <= 32'b00000000010000010000000100010011;
ROM[10522] <= 32'b00000000001100010010000000100011;
ROM[10523] <= 32'b00000000010000010000000100010011;
ROM[10524] <= 32'b00000000010000010010000000100011;
ROM[10525] <= 32'b00000000010000010000000100010011;
ROM[10526] <= 32'b00000000010100010010000000100011;
ROM[10527] <= 32'b00000000010000010000000100010011;
ROM[10528] <= 32'b00000000011000010010000000100011;
ROM[10529] <= 32'b00000000010000010000000100010011;
ROM[10530] <= 32'b00000001010000000000001110010011;
ROM[10531] <= 32'b00000000100000111000001110010011;
ROM[10532] <= 32'b01000000011100010000001110110011;
ROM[10533] <= 32'b00000000011100000000001000110011;
ROM[10534] <= 32'b00000000001000000000000110110011;
ROM[10535] <= 32'b01110001000000011111000011101111;
ROM[10536] <= 32'b00000110100100000000001110010011;
ROM[10537] <= 32'b00000000011100010010000000100011;
ROM[10538] <= 32'b00000000010000010000000100010011;
ROM[10539] <= 32'b00000000000000001010001110110111;
ROM[10540] <= 32'b01001111100000111000001110010011;
ROM[10541] <= 32'b00000000111000111000001110110011;
ROM[10542] <= 32'b00000000011100010010000000100011;
ROM[10543] <= 32'b00000000010000010000000100010011;
ROM[10544] <= 32'b00000000001100010010000000100011;
ROM[10545] <= 32'b00000000010000010000000100010011;
ROM[10546] <= 32'b00000000010000010010000000100011;
ROM[10547] <= 32'b00000000010000010000000100010011;
ROM[10548] <= 32'b00000000010100010010000000100011;
ROM[10549] <= 32'b00000000010000010000000100010011;
ROM[10550] <= 32'b00000000011000010010000000100011;
ROM[10551] <= 32'b00000000010000010000000100010011;
ROM[10552] <= 32'b00000001010000000000001110010011;
ROM[10553] <= 32'b00000000100000111000001110010011;
ROM[10554] <= 32'b01000000011100010000001110110011;
ROM[10555] <= 32'b00000000011100000000001000110011;
ROM[10556] <= 32'b00000000001000000000000110110011;
ROM[10557] <= 32'b01101011100000011111000011101111;
ROM[10558] <= 32'b00000111001100000000001110010011;
ROM[10559] <= 32'b00000000011100010010000000100011;
ROM[10560] <= 32'b00000000010000010000000100010011;
ROM[10561] <= 32'b00000000000000001010001110110111;
ROM[10562] <= 32'b01010101000000111000001110010011;
ROM[10563] <= 32'b00000000111000111000001110110011;
ROM[10564] <= 32'b00000000011100010010000000100011;
ROM[10565] <= 32'b00000000010000010000000100010011;
ROM[10566] <= 32'b00000000001100010010000000100011;
ROM[10567] <= 32'b00000000010000010000000100010011;
ROM[10568] <= 32'b00000000010000010010000000100011;
ROM[10569] <= 32'b00000000010000010000000100010011;
ROM[10570] <= 32'b00000000010100010010000000100011;
ROM[10571] <= 32'b00000000010000010000000100010011;
ROM[10572] <= 32'b00000000011000010010000000100011;
ROM[10573] <= 32'b00000000010000010000000100010011;
ROM[10574] <= 32'b00000001010000000000001110010011;
ROM[10575] <= 32'b00000000100000111000001110010011;
ROM[10576] <= 32'b01000000011100010000001110110011;
ROM[10577] <= 32'b00000000011100000000001000110011;
ROM[10578] <= 32'b00000000001000000000000110110011;
ROM[10579] <= 32'b01100110000000011111000011101111;
ROM[10580] <= 32'b00000010000000000000001110010011;
ROM[10581] <= 32'b00000000011100010010000000100011;
ROM[10582] <= 32'b00000000010000010000000100010011;
ROM[10583] <= 32'b00000000000000001010001110110111;
ROM[10584] <= 32'b01011010100000111000001110010011;
ROM[10585] <= 32'b00000000111000111000001110110011;
ROM[10586] <= 32'b00000000011100010010000000100011;
ROM[10587] <= 32'b00000000010000010000000100010011;
ROM[10588] <= 32'b00000000001100010010000000100011;
ROM[10589] <= 32'b00000000010000010000000100010011;
ROM[10590] <= 32'b00000000010000010010000000100011;
ROM[10591] <= 32'b00000000010000010000000100010011;
ROM[10592] <= 32'b00000000010100010010000000100011;
ROM[10593] <= 32'b00000000010000010000000100010011;
ROM[10594] <= 32'b00000000011000010010000000100011;
ROM[10595] <= 32'b00000000010000010000000100010011;
ROM[10596] <= 32'b00000001010000000000001110010011;
ROM[10597] <= 32'b00000000100000111000001110010011;
ROM[10598] <= 32'b01000000011100010000001110110011;
ROM[10599] <= 32'b00000000011100000000001000110011;
ROM[10600] <= 32'b00000000001000000000000110110011;
ROM[10601] <= 32'b01100000100000011111000011101111;
ROM[10602] <= 32'b00000000000000001010001110110111;
ROM[10603] <= 32'b01011111010000111000001110010011;
ROM[10604] <= 32'b00000000111000111000001110110011;
ROM[10605] <= 32'b00000000011100010010000000100011;
ROM[10606] <= 32'b00000000010000010000000100010011;
ROM[10607] <= 32'b00000000001100010010000000100011;
ROM[10608] <= 32'b00000000010000010000000100010011;
ROM[10609] <= 32'b00000000010000010010000000100011;
ROM[10610] <= 32'b00000000010000010000000100010011;
ROM[10611] <= 32'b00000000010100010010000000100011;
ROM[10612] <= 32'b00000000010000010000000100010011;
ROM[10613] <= 32'b00000000011000010010000000100011;
ROM[10614] <= 32'b00000000010000010000000100010011;
ROM[10615] <= 32'b00000001010000000000001110010011;
ROM[10616] <= 32'b00000000010000111000001110010011;
ROM[10617] <= 32'b01000000011100010000001110110011;
ROM[10618] <= 32'b00000000011100000000001000110011;
ROM[10619] <= 32'b00000000001000000000000110110011;
ROM[10620] <= 32'b00010111100100001100000011101111;
ROM[10621] <= 32'b11111111110000010000000100010011;
ROM[10622] <= 32'b00000000000000010010001110000011;
ROM[10623] <= 32'b00000000011101100010000000100011;
ROM[10624] <= 32'b00000001100000011010001110000011;
ROM[10625] <= 32'b00000000011100010010000000100011;
ROM[10626] <= 32'b00000000010000010000000100010011;
ROM[10627] <= 32'b00000000000000001010001110110111;
ROM[10628] <= 32'b01100101100000111000001110010011;
ROM[10629] <= 32'b00000000111000111000001110110011;
ROM[10630] <= 32'b00000000011100010010000000100011;
ROM[10631] <= 32'b00000000010000010000000100010011;
ROM[10632] <= 32'b00000000001100010010000000100011;
ROM[10633] <= 32'b00000000010000010000000100010011;
ROM[10634] <= 32'b00000000010000010010000000100011;
ROM[10635] <= 32'b00000000010000010000000100010011;
ROM[10636] <= 32'b00000000010100010010000000100011;
ROM[10637] <= 32'b00000000010000010000000100010011;
ROM[10638] <= 32'b00000000011000010010000000100011;
ROM[10639] <= 32'b00000000010000010000000100010011;
ROM[10640] <= 32'b00000001010000000000001110010011;
ROM[10641] <= 32'b00000000010000111000001110010011;
ROM[10642] <= 32'b01000000011100010000001110110011;
ROM[10643] <= 32'b00000000011100000000001000110011;
ROM[10644] <= 32'b00000000001000000000000110110011;
ROM[10645] <= 32'b00010001010100001100000011101111;
ROM[10646] <= 32'b11111111110000010000000100010011;
ROM[10647] <= 32'b00000000000000010010001110000011;
ROM[10648] <= 32'b00000000011101100010000000100011;
ROM[10649] <= 32'b00000000000000001010001110110111;
ROM[10650] <= 32'b01101011000000111000001110010011;
ROM[10651] <= 32'b00000000111000111000001110110011;
ROM[10652] <= 32'b00000000011100010010000000100011;
ROM[10653] <= 32'b00000000010000010000000100010011;
ROM[10654] <= 32'b00000000001100010010000000100011;
ROM[10655] <= 32'b00000000010000010000000100010011;
ROM[10656] <= 32'b00000000010000010010000000100011;
ROM[10657] <= 32'b00000000010000010000000100010011;
ROM[10658] <= 32'b00000000010100010010000000100011;
ROM[10659] <= 32'b00000000010000010000000100010011;
ROM[10660] <= 32'b00000000011000010010000000100011;
ROM[10661] <= 32'b00000000010000010000000100010011;
ROM[10662] <= 32'b00000001010000000000001110010011;
ROM[10663] <= 32'b00000000000000111000001110010011;
ROM[10664] <= 32'b01000000011100010000001110110011;
ROM[10665] <= 32'b00000000011100000000001000110011;
ROM[10666] <= 32'b00000000001000000000000110110011;
ROM[10667] <= 32'b01001011110100001100000011101111;
ROM[10668] <= 32'b11111111110000010000000100010011;
ROM[10669] <= 32'b00000000000000010010001110000011;
ROM[10670] <= 32'b00000000011101100010000000100011;
ROM[10671] <= 32'b01111001110100000001000011101111;
ROM[10672] <= 32'b00000001010000011010001110000011;
ROM[10673] <= 32'b00000000011100010010000000100011;
ROM[10674] <= 32'b00000000010000010000000100010011;
ROM[10675] <= 32'b00000000000100000000001110010011;
ROM[10676] <= 32'b00000000011100010010000000100011;
ROM[10677] <= 32'b00000000010000010000000100010011;
ROM[10678] <= 32'b11111111110000010000000100010011;
ROM[10679] <= 32'b00000000000000010010001110000011;
ROM[10680] <= 32'b11111111110000010000000100010011;
ROM[10681] <= 32'b00000000000000010010010000000011;
ROM[10682] <= 32'b00000000011101000010010010110011;
ROM[10683] <= 32'b00000000100000111010010100110011;
ROM[10684] <= 32'b00000000101001001000001110110011;
ROM[10685] <= 32'b00000000000100111000001110010011;
ROM[10686] <= 32'b00000000000100111111001110010011;
ROM[10687] <= 32'b00000000011100010010000000100011;
ROM[10688] <= 32'b00000000010000010000000100010011;
ROM[10689] <= 32'b11111111110000010000000100010011;
ROM[10690] <= 32'b00000000000000010010001110000011;
ROM[10691] <= 32'b00000000000000111000101001100011;
ROM[10692] <= 32'b00000000000000001011001110110111;
ROM[10693] <= 32'b01110101100000111000001110010011;
ROM[10694] <= 32'b00000000111000111000001110110011;
ROM[10695] <= 32'b00000000000000111000000011100111;
ROM[10696] <= 32'b00000001011000000000001110010011;
ROM[10697] <= 32'b00000000011100010010000000100011;
ROM[10698] <= 32'b00000000010000010000000100010011;
ROM[10699] <= 32'b00000000000000001010001110110111;
ROM[10700] <= 32'b01110111100000111000001110010011;
ROM[10701] <= 32'b00000000111000111000001110110011;
ROM[10702] <= 32'b00000000011100010010000000100011;
ROM[10703] <= 32'b00000000010000010000000100010011;
ROM[10704] <= 32'b00000000001100010010000000100011;
ROM[10705] <= 32'b00000000010000010000000100010011;
ROM[10706] <= 32'b00000000010000010010000000100011;
ROM[10707] <= 32'b00000000010000010000000100010011;
ROM[10708] <= 32'b00000000010100010010000000100011;
ROM[10709] <= 32'b00000000010000010000000100010011;
ROM[10710] <= 32'b00000000011000010010000000100011;
ROM[10711] <= 32'b00000000010000010000000100010011;
ROM[10712] <= 32'b00000001010000000000001110010011;
ROM[10713] <= 32'b00000000010000111000001110010011;
ROM[10714] <= 32'b01000000011100010000001110110011;
ROM[10715] <= 32'b00000000011100000000001000110011;
ROM[10716] <= 32'b00000000001000000000000110110011;
ROM[10717] <= 32'b01111100100100011110000011101111;
ROM[10718] <= 32'b00000101011100000000001110010011;
ROM[10719] <= 32'b00000000011100010010000000100011;
ROM[10720] <= 32'b00000000010000010000000100010011;
ROM[10721] <= 32'b00000000000000001010001110110111;
ROM[10722] <= 32'b01111101000000111000001110010011;
ROM[10723] <= 32'b00000000111000111000001110110011;
ROM[10724] <= 32'b00000000011100010010000000100011;
ROM[10725] <= 32'b00000000010000010000000100010011;
ROM[10726] <= 32'b00000000001100010010000000100011;
ROM[10727] <= 32'b00000000010000010000000100010011;
ROM[10728] <= 32'b00000000010000010010000000100011;
ROM[10729] <= 32'b00000000010000010000000100010011;
ROM[10730] <= 32'b00000000010100010010000000100011;
ROM[10731] <= 32'b00000000010000010000000100010011;
ROM[10732] <= 32'b00000000011000010010000000100011;
ROM[10733] <= 32'b00000000010000010000000100010011;
ROM[10734] <= 32'b00000001010000000000001110010011;
ROM[10735] <= 32'b00000000100000111000001110010011;
ROM[10736] <= 32'b01000000011100010000001110110011;
ROM[10737] <= 32'b00000000011100000000001000110011;
ROM[10738] <= 32'b00000000001000000000000110110011;
ROM[10739] <= 32'b00111110000000011111000011101111;
ROM[10740] <= 32'b00000111001000000000001110010011;
ROM[10741] <= 32'b00000000011100010010000000100011;
ROM[10742] <= 32'b00000000010000010000000100010011;
ROM[10743] <= 32'b00000000000000001011001110110111;
ROM[10744] <= 32'b10000010100000111000001110010011;
ROM[10745] <= 32'b00000000111000111000001110110011;
ROM[10746] <= 32'b00000000011100010010000000100011;
ROM[10747] <= 32'b00000000010000010000000100010011;
ROM[10748] <= 32'b00000000001100010010000000100011;
ROM[10749] <= 32'b00000000010000010000000100010011;
ROM[10750] <= 32'b00000000010000010010000000100011;
ROM[10751] <= 32'b00000000010000010000000100010011;
ROM[10752] <= 32'b00000000010100010010000000100011;
ROM[10753] <= 32'b00000000010000010000000100010011;
ROM[10754] <= 32'b00000000011000010010000000100011;
ROM[10755] <= 32'b00000000010000010000000100010011;
ROM[10756] <= 32'b00000001010000000000001110010011;
ROM[10757] <= 32'b00000000100000111000001110010011;
ROM[10758] <= 32'b01000000011100010000001110110011;
ROM[10759] <= 32'b00000000011100000000001000110011;
ROM[10760] <= 32'b00000000001000000000000110110011;
ROM[10761] <= 32'b00111000100000011111000011101111;
ROM[10762] <= 32'b00000110111100000000001110010011;
ROM[10763] <= 32'b00000000011100010010000000100011;
ROM[10764] <= 32'b00000000010000010000000100010011;
ROM[10765] <= 32'b00000000000000001011001110110111;
ROM[10766] <= 32'b10001000000000111000001110010011;
ROM[10767] <= 32'b00000000111000111000001110110011;
ROM[10768] <= 32'b00000000011100010010000000100011;
ROM[10769] <= 32'b00000000010000010000000100010011;
ROM[10770] <= 32'b00000000001100010010000000100011;
ROM[10771] <= 32'b00000000010000010000000100010011;
ROM[10772] <= 32'b00000000010000010010000000100011;
ROM[10773] <= 32'b00000000010000010000000100010011;
ROM[10774] <= 32'b00000000010100010010000000100011;
ROM[10775] <= 32'b00000000010000010000000100010011;
ROM[10776] <= 32'b00000000011000010010000000100011;
ROM[10777] <= 32'b00000000010000010000000100010011;
ROM[10778] <= 32'b00000001010000000000001110010011;
ROM[10779] <= 32'b00000000100000111000001110010011;
ROM[10780] <= 32'b01000000011100010000001110110011;
ROM[10781] <= 32'b00000000011100000000001000110011;
ROM[10782] <= 32'b00000000001000000000000110110011;
ROM[10783] <= 32'b00110011000000011111000011101111;
ROM[10784] <= 32'b00000110111000000000001110010011;
ROM[10785] <= 32'b00000000011100010010000000100011;
ROM[10786] <= 32'b00000000010000010000000100010011;
ROM[10787] <= 32'b00000000000000001011001110110111;
ROM[10788] <= 32'b10001101100000111000001110010011;
ROM[10789] <= 32'b00000000111000111000001110110011;
ROM[10790] <= 32'b00000000011100010010000000100011;
ROM[10791] <= 32'b00000000010000010000000100010011;
ROM[10792] <= 32'b00000000001100010010000000100011;
ROM[10793] <= 32'b00000000010000010000000100010011;
ROM[10794] <= 32'b00000000010000010010000000100011;
ROM[10795] <= 32'b00000000010000010000000100010011;
ROM[10796] <= 32'b00000000010100010010000000100011;
ROM[10797] <= 32'b00000000010000010000000100010011;
ROM[10798] <= 32'b00000000011000010010000000100011;
ROM[10799] <= 32'b00000000010000010000000100010011;
ROM[10800] <= 32'b00000001010000000000001110010011;
ROM[10801] <= 32'b00000000100000111000001110010011;
ROM[10802] <= 32'b01000000011100010000001110110011;
ROM[10803] <= 32'b00000000011100000000001000110011;
ROM[10804] <= 32'b00000000001000000000000110110011;
ROM[10805] <= 32'b00101101100000011111000011101111;
ROM[10806] <= 32'b00000110011100000000001110010011;
ROM[10807] <= 32'b00000000011100010010000000100011;
ROM[10808] <= 32'b00000000010000010000000100010011;
ROM[10809] <= 32'b00000000000000001011001110110111;
ROM[10810] <= 32'b10010011000000111000001110010011;
ROM[10811] <= 32'b00000000111000111000001110110011;
ROM[10812] <= 32'b00000000011100010010000000100011;
ROM[10813] <= 32'b00000000010000010000000100010011;
ROM[10814] <= 32'b00000000001100010010000000100011;
ROM[10815] <= 32'b00000000010000010000000100010011;
ROM[10816] <= 32'b00000000010000010010000000100011;
ROM[10817] <= 32'b00000000010000010000000100010011;
ROM[10818] <= 32'b00000000010100010010000000100011;
ROM[10819] <= 32'b00000000010000010000000100010011;
ROM[10820] <= 32'b00000000011000010010000000100011;
ROM[10821] <= 32'b00000000010000010000000100010011;
ROM[10822] <= 32'b00000001010000000000001110010011;
ROM[10823] <= 32'b00000000100000111000001110010011;
ROM[10824] <= 32'b01000000011100010000001110110011;
ROM[10825] <= 32'b00000000011100000000001000110011;
ROM[10826] <= 32'b00000000001000000000000110110011;
ROM[10827] <= 32'b00101000000000011111000011101111;
ROM[10828] <= 32'b00000010000000000000001110010011;
ROM[10829] <= 32'b00000000011100010010000000100011;
ROM[10830] <= 32'b00000000010000010000000100010011;
ROM[10831] <= 32'b00000000000000001011001110110111;
ROM[10832] <= 32'b10011000100000111000001110010011;
ROM[10833] <= 32'b00000000111000111000001110110011;
ROM[10834] <= 32'b00000000011100010010000000100011;
ROM[10835] <= 32'b00000000010000010000000100010011;
ROM[10836] <= 32'b00000000001100010010000000100011;
ROM[10837] <= 32'b00000000010000010000000100010011;
ROM[10838] <= 32'b00000000010000010010000000100011;
ROM[10839] <= 32'b00000000010000010000000100010011;
ROM[10840] <= 32'b00000000010100010010000000100011;
ROM[10841] <= 32'b00000000010000010000000100010011;
ROM[10842] <= 32'b00000000011000010010000000100011;
ROM[10843] <= 32'b00000000010000010000000100010011;
ROM[10844] <= 32'b00000001010000000000001110010011;
ROM[10845] <= 32'b00000000100000111000001110010011;
ROM[10846] <= 32'b01000000011100010000001110110011;
ROM[10847] <= 32'b00000000011100000000001000110011;
ROM[10848] <= 32'b00000000001000000000000110110011;
ROM[10849] <= 32'b00100010100000011111000011101111;
ROM[10850] <= 32'b00000110011100000000001110010011;
ROM[10851] <= 32'b00000000011100010010000000100011;
ROM[10852] <= 32'b00000000010000010000000100010011;
ROM[10853] <= 32'b00000000000000001011001110110111;
ROM[10854] <= 32'b10011110000000111000001110010011;
ROM[10855] <= 32'b00000000111000111000001110110011;
ROM[10856] <= 32'b00000000011100010010000000100011;
ROM[10857] <= 32'b00000000010000010000000100010011;
ROM[10858] <= 32'b00000000001100010010000000100011;
ROM[10859] <= 32'b00000000010000010000000100010011;
ROM[10860] <= 32'b00000000010000010010000000100011;
ROM[10861] <= 32'b00000000010000010000000100010011;
ROM[10862] <= 32'b00000000010100010010000000100011;
ROM[10863] <= 32'b00000000010000010000000100010011;
ROM[10864] <= 32'b00000000011000010010000000100011;
ROM[10865] <= 32'b00000000010000010000000100010011;
ROM[10866] <= 32'b00000001010000000000001110010011;
ROM[10867] <= 32'b00000000100000111000001110010011;
ROM[10868] <= 32'b01000000011100010000001110110011;
ROM[10869] <= 32'b00000000011100000000001000110011;
ROM[10870] <= 32'b00000000001000000000000110110011;
ROM[10871] <= 32'b00011101000000011111000011101111;
ROM[10872] <= 32'b00000111010100000000001110010011;
ROM[10873] <= 32'b00000000011100010010000000100011;
ROM[10874] <= 32'b00000000010000010000000100010011;
ROM[10875] <= 32'b00000000000000001011001110110111;
ROM[10876] <= 32'b10100011100000111000001110010011;
ROM[10877] <= 32'b00000000111000111000001110110011;
ROM[10878] <= 32'b00000000011100010010000000100011;
ROM[10879] <= 32'b00000000010000010000000100010011;
ROM[10880] <= 32'b00000000001100010010000000100011;
ROM[10881] <= 32'b00000000010000010000000100010011;
ROM[10882] <= 32'b00000000010000010010000000100011;
ROM[10883] <= 32'b00000000010000010000000100010011;
ROM[10884] <= 32'b00000000010100010010000000100011;
ROM[10885] <= 32'b00000000010000010000000100010011;
ROM[10886] <= 32'b00000000011000010010000000100011;
ROM[10887] <= 32'b00000000010000010000000100010011;
ROM[10888] <= 32'b00000001010000000000001110010011;
ROM[10889] <= 32'b00000000100000111000001110010011;
ROM[10890] <= 32'b01000000011100010000001110110011;
ROM[10891] <= 32'b00000000011100000000001000110011;
ROM[10892] <= 32'b00000000001000000000000110110011;
ROM[10893] <= 32'b00010111100000011111000011101111;
ROM[10894] <= 32'b00000110010100000000001110010011;
ROM[10895] <= 32'b00000000011100010010000000100011;
ROM[10896] <= 32'b00000000010000010000000100010011;
ROM[10897] <= 32'b00000000000000001011001110110111;
ROM[10898] <= 32'b10101001000000111000001110010011;
ROM[10899] <= 32'b00000000111000111000001110110011;
ROM[10900] <= 32'b00000000011100010010000000100011;
ROM[10901] <= 32'b00000000010000010000000100010011;
ROM[10902] <= 32'b00000000001100010010000000100011;
ROM[10903] <= 32'b00000000010000010000000100010011;
ROM[10904] <= 32'b00000000010000010010000000100011;
ROM[10905] <= 32'b00000000010000010000000100010011;
ROM[10906] <= 32'b00000000010100010010000000100011;
ROM[10907] <= 32'b00000000010000010000000100010011;
ROM[10908] <= 32'b00000000011000010010000000100011;
ROM[10909] <= 32'b00000000010000010000000100010011;
ROM[10910] <= 32'b00000001010000000000001110010011;
ROM[10911] <= 32'b00000000100000111000001110010011;
ROM[10912] <= 32'b01000000011100010000001110110011;
ROM[10913] <= 32'b00000000011100000000001000110011;
ROM[10914] <= 32'b00000000001000000000000110110011;
ROM[10915] <= 32'b00010010000000011111000011101111;
ROM[10916] <= 32'b00000111001100000000001110010011;
ROM[10917] <= 32'b00000000011100010010000000100011;
ROM[10918] <= 32'b00000000010000010000000100010011;
ROM[10919] <= 32'b00000000000000001011001110110111;
ROM[10920] <= 32'b10101110100000111000001110010011;
ROM[10921] <= 32'b00000000111000111000001110110011;
ROM[10922] <= 32'b00000000011100010010000000100011;
ROM[10923] <= 32'b00000000010000010000000100010011;
ROM[10924] <= 32'b00000000001100010010000000100011;
ROM[10925] <= 32'b00000000010000010000000100010011;
ROM[10926] <= 32'b00000000010000010010000000100011;
ROM[10927] <= 32'b00000000010000010000000100010011;
ROM[10928] <= 32'b00000000010100010010000000100011;
ROM[10929] <= 32'b00000000010000010000000100010011;
ROM[10930] <= 32'b00000000011000010010000000100011;
ROM[10931] <= 32'b00000000010000010000000100010011;
ROM[10932] <= 32'b00000001010000000000001110010011;
ROM[10933] <= 32'b00000000100000111000001110010011;
ROM[10934] <= 32'b01000000011100010000001110110011;
ROM[10935] <= 32'b00000000011100000000001000110011;
ROM[10936] <= 32'b00000000001000000000000110110011;
ROM[10937] <= 32'b00001100100000011111000011101111;
ROM[10938] <= 32'b00000111001100000000001110010011;
ROM[10939] <= 32'b00000000011100010010000000100011;
ROM[10940] <= 32'b00000000010000010000000100010011;
ROM[10941] <= 32'b00000000000000001011001110110111;
ROM[10942] <= 32'b10110100000000111000001110010011;
ROM[10943] <= 32'b00000000111000111000001110110011;
ROM[10944] <= 32'b00000000011100010010000000100011;
ROM[10945] <= 32'b00000000010000010000000100010011;
ROM[10946] <= 32'b00000000001100010010000000100011;
ROM[10947] <= 32'b00000000010000010000000100010011;
ROM[10948] <= 32'b00000000010000010010000000100011;
ROM[10949] <= 32'b00000000010000010000000100010011;
ROM[10950] <= 32'b00000000010100010010000000100011;
ROM[10951] <= 32'b00000000010000010000000100010011;
ROM[10952] <= 32'b00000000011000010010000000100011;
ROM[10953] <= 32'b00000000010000010000000100010011;
ROM[10954] <= 32'b00000001010000000000001110010011;
ROM[10955] <= 32'b00000000100000111000001110010011;
ROM[10956] <= 32'b01000000011100010000001110110011;
ROM[10957] <= 32'b00000000011100000000001000110011;
ROM[10958] <= 32'b00000000001000000000000110110011;
ROM[10959] <= 32'b00000111000000011111000011101111;
ROM[10960] <= 32'b00000010110000000000001110010011;
ROM[10961] <= 32'b00000000011100010010000000100011;
ROM[10962] <= 32'b00000000010000010000000100010011;
ROM[10963] <= 32'b00000000000000001011001110110111;
ROM[10964] <= 32'b10111001100000111000001110010011;
ROM[10965] <= 32'b00000000111000111000001110110011;
ROM[10966] <= 32'b00000000011100010010000000100011;
ROM[10967] <= 32'b00000000010000010000000100010011;
ROM[10968] <= 32'b00000000001100010010000000100011;
ROM[10969] <= 32'b00000000010000010000000100010011;
ROM[10970] <= 32'b00000000010000010010000000100011;
ROM[10971] <= 32'b00000000010000010000000100010011;
ROM[10972] <= 32'b00000000010100010010000000100011;
ROM[10973] <= 32'b00000000010000010000000100010011;
ROM[10974] <= 32'b00000000011000010010000000100011;
ROM[10975] <= 32'b00000000010000010000000100010011;
ROM[10976] <= 32'b00000001010000000000001110010011;
ROM[10977] <= 32'b00000000100000111000001110010011;
ROM[10978] <= 32'b01000000011100010000001110110011;
ROM[10979] <= 32'b00000000011100000000001000110011;
ROM[10980] <= 32'b00000000001000000000000110110011;
ROM[10981] <= 32'b00000001100000011111000011101111;
ROM[10982] <= 32'b00000010000000000000001110010011;
ROM[10983] <= 32'b00000000011100010010000000100011;
ROM[10984] <= 32'b00000000010000010000000100010011;
ROM[10985] <= 32'b00000000000000001011001110110111;
ROM[10986] <= 32'b10111111000000111000001110010011;
ROM[10987] <= 32'b00000000111000111000001110110011;
ROM[10988] <= 32'b00000000011100010010000000100011;
ROM[10989] <= 32'b00000000010000010000000100010011;
ROM[10990] <= 32'b00000000001100010010000000100011;
ROM[10991] <= 32'b00000000010000010000000100010011;
ROM[10992] <= 32'b00000000010000010010000000100011;
ROM[10993] <= 32'b00000000010000010000000100010011;
ROM[10994] <= 32'b00000000010100010010000000100011;
ROM[10995] <= 32'b00000000010000010000000100010011;
ROM[10996] <= 32'b00000000011000010010000000100011;
ROM[10997] <= 32'b00000000010000010000000100010011;
ROM[10998] <= 32'b00000001010000000000001110010011;
ROM[10999] <= 32'b00000000100000111000001110010011;
ROM[11000] <= 32'b01000000011100010000001110110011;
ROM[11001] <= 32'b00000000011100000000001000110011;
ROM[11002] <= 32'b00000000001000000000000110110011;
ROM[11003] <= 32'b01111100000100011110000011101111;
ROM[11004] <= 32'b00000111100100000000001110010011;
ROM[11005] <= 32'b00000000011100010010000000100011;
ROM[11006] <= 32'b00000000010000010000000100010011;
ROM[11007] <= 32'b00000000000000001011001110110111;
ROM[11008] <= 32'b11000100100000111000001110010011;
ROM[11009] <= 32'b00000000111000111000001110110011;
ROM[11010] <= 32'b00000000011100010010000000100011;
ROM[11011] <= 32'b00000000010000010000000100010011;
ROM[11012] <= 32'b00000000001100010010000000100011;
ROM[11013] <= 32'b00000000010000010000000100010011;
ROM[11014] <= 32'b00000000010000010010000000100011;
ROM[11015] <= 32'b00000000010000010000000100010011;
ROM[11016] <= 32'b00000000010100010010000000100011;
ROM[11017] <= 32'b00000000010000010000000100010011;
ROM[11018] <= 32'b00000000011000010010000000100011;
ROM[11019] <= 32'b00000000010000010000000100010011;
ROM[11020] <= 32'b00000001010000000000001110010011;
ROM[11021] <= 32'b00000000100000111000001110010011;
ROM[11022] <= 32'b01000000011100010000001110110011;
ROM[11023] <= 32'b00000000011100000000001000110011;
ROM[11024] <= 32'b00000000001000000000000110110011;
ROM[11025] <= 32'b01110110100100011110000011101111;
ROM[11026] <= 32'b00000110111100000000001110010011;
ROM[11027] <= 32'b00000000011100010010000000100011;
ROM[11028] <= 32'b00000000010000010000000100010011;
ROM[11029] <= 32'b00000000000000001011001110110111;
ROM[11030] <= 32'b11001010000000111000001110010011;
ROM[11031] <= 32'b00000000111000111000001110110011;
ROM[11032] <= 32'b00000000011100010010000000100011;
ROM[11033] <= 32'b00000000010000010000000100010011;
ROM[11034] <= 32'b00000000001100010010000000100011;
ROM[11035] <= 32'b00000000010000010000000100010011;
ROM[11036] <= 32'b00000000010000010010000000100011;
ROM[11037] <= 32'b00000000010000010000000100010011;
ROM[11038] <= 32'b00000000010100010010000000100011;
ROM[11039] <= 32'b00000000010000010000000100010011;
ROM[11040] <= 32'b00000000011000010010000000100011;
ROM[11041] <= 32'b00000000010000010000000100010011;
ROM[11042] <= 32'b00000001010000000000001110010011;
ROM[11043] <= 32'b00000000100000111000001110010011;
ROM[11044] <= 32'b01000000011100010000001110110011;
ROM[11045] <= 32'b00000000011100000000001000110011;
ROM[11046] <= 32'b00000000001000000000000110110011;
ROM[11047] <= 32'b01110001000100011110000011101111;
ROM[11048] <= 32'b00000111010100000000001110010011;
ROM[11049] <= 32'b00000000011100010010000000100011;
ROM[11050] <= 32'b00000000010000010000000100010011;
ROM[11051] <= 32'b00000000000000001011001110110111;
ROM[11052] <= 32'b11001111100000111000001110010011;
ROM[11053] <= 32'b00000000111000111000001110110011;
ROM[11054] <= 32'b00000000011100010010000000100011;
ROM[11055] <= 32'b00000000010000010000000100010011;
ROM[11056] <= 32'b00000000001100010010000000100011;
ROM[11057] <= 32'b00000000010000010000000100010011;
ROM[11058] <= 32'b00000000010000010010000000100011;
ROM[11059] <= 32'b00000000010000010000000100010011;
ROM[11060] <= 32'b00000000010100010010000000100011;
ROM[11061] <= 32'b00000000010000010000000100010011;
ROM[11062] <= 32'b00000000011000010010000000100011;
ROM[11063] <= 32'b00000000010000010000000100010011;
ROM[11064] <= 32'b00000001010000000000001110010011;
ROM[11065] <= 32'b00000000100000111000001110010011;
ROM[11066] <= 32'b01000000011100010000001110110011;
ROM[11067] <= 32'b00000000011100000000001000110011;
ROM[11068] <= 32'b00000000001000000000000110110011;
ROM[11069] <= 32'b01101011100100011110000011101111;
ROM[11070] <= 32'b00000010000000000000001110010011;
ROM[11071] <= 32'b00000000011100010010000000100011;
ROM[11072] <= 32'b00000000010000010000000100010011;
ROM[11073] <= 32'b00000000000000001011001110110111;
ROM[11074] <= 32'b11010101000000111000001110010011;
ROM[11075] <= 32'b00000000111000111000001110110011;
ROM[11076] <= 32'b00000000011100010010000000100011;
ROM[11077] <= 32'b00000000010000010000000100010011;
ROM[11078] <= 32'b00000000001100010010000000100011;
ROM[11079] <= 32'b00000000010000010000000100010011;
ROM[11080] <= 32'b00000000010000010010000000100011;
ROM[11081] <= 32'b00000000010000010000000100010011;
ROM[11082] <= 32'b00000000010100010010000000100011;
ROM[11083] <= 32'b00000000010000010000000100010011;
ROM[11084] <= 32'b00000000011000010010000000100011;
ROM[11085] <= 32'b00000000010000010000000100010011;
ROM[11086] <= 32'b00000001010000000000001110010011;
ROM[11087] <= 32'b00000000100000111000001110010011;
ROM[11088] <= 32'b01000000011100010000001110110011;
ROM[11089] <= 32'b00000000011100000000001000110011;
ROM[11090] <= 32'b00000000001000000000000110110011;
ROM[11091] <= 32'b01100110000100011110000011101111;
ROM[11092] <= 32'b00000110100000000000001110010011;
ROM[11093] <= 32'b00000000011100010010000000100011;
ROM[11094] <= 32'b00000000010000010000000100010011;
ROM[11095] <= 32'b00000000000000001011001110110111;
ROM[11096] <= 32'b11011010100000111000001110010011;
ROM[11097] <= 32'b00000000111000111000001110110011;
ROM[11098] <= 32'b00000000011100010010000000100011;
ROM[11099] <= 32'b00000000010000010000000100010011;
ROM[11100] <= 32'b00000000001100010010000000100011;
ROM[11101] <= 32'b00000000010000010000000100010011;
ROM[11102] <= 32'b00000000010000010010000000100011;
ROM[11103] <= 32'b00000000010000010000000100010011;
ROM[11104] <= 32'b00000000010100010010000000100011;
ROM[11105] <= 32'b00000000010000010000000100010011;
ROM[11106] <= 32'b00000000011000010010000000100011;
ROM[11107] <= 32'b00000000010000010000000100010011;
ROM[11108] <= 32'b00000001010000000000001110010011;
ROM[11109] <= 32'b00000000100000111000001110010011;
ROM[11110] <= 32'b01000000011100010000001110110011;
ROM[11111] <= 32'b00000000011100000000001000110011;
ROM[11112] <= 32'b00000000001000000000000110110011;
ROM[11113] <= 32'b01100000100100011110000011101111;
ROM[11114] <= 32'b00000110000100000000001110010011;
ROM[11115] <= 32'b00000000011100010010000000100011;
ROM[11116] <= 32'b00000000010000010000000100010011;
ROM[11117] <= 32'b00000000000000001011001110110111;
ROM[11118] <= 32'b11100000000000111000001110010011;
ROM[11119] <= 32'b00000000111000111000001110110011;
ROM[11120] <= 32'b00000000011100010010000000100011;
ROM[11121] <= 32'b00000000010000010000000100010011;
ROM[11122] <= 32'b00000000001100010010000000100011;
ROM[11123] <= 32'b00000000010000010000000100010011;
ROM[11124] <= 32'b00000000010000010010000000100011;
ROM[11125] <= 32'b00000000010000010000000100010011;
ROM[11126] <= 32'b00000000010100010010000000100011;
ROM[11127] <= 32'b00000000010000010000000100010011;
ROM[11128] <= 32'b00000000011000010010000000100011;
ROM[11129] <= 32'b00000000010000010000000100010011;
ROM[11130] <= 32'b00000001010000000000001110010011;
ROM[11131] <= 32'b00000000100000111000001110010011;
ROM[11132] <= 32'b01000000011100010000001110110011;
ROM[11133] <= 32'b00000000011100000000001000110011;
ROM[11134] <= 32'b00000000001000000000000110110011;
ROM[11135] <= 32'b01011011000100011110000011101111;
ROM[11136] <= 32'b00000111011000000000001110010011;
ROM[11137] <= 32'b00000000011100010010000000100011;
ROM[11138] <= 32'b00000000010000010000000100010011;
ROM[11139] <= 32'b00000000000000001011001110110111;
ROM[11140] <= 32'b11100101100000111000001110010011;
ROM[11141] <= 32'b00000000111000111000001110110011;
ROM[11142] <= 32'b00000000011100010010000000100011;
ROM[11143] <= 32'b00000000010000010000000100010011;
ROM[11144] <= 32'b00000000001100010010000000100011;
ROM[11145] <= 32'b00000000010000010000000100010011;
ROM[11146] <= 32'b00000000010000010010000000100011;
ROM[11147] <= 32'b00000000010000010000000100010011;
ROM[11148] <= 32'b00000000010100010010000000100011;
ROM[11149] <= 32'b00000000010000010000000100010011;
ROM[11150] <= 32'b00000000011000010010000000100011;
ROM[11151] <= 32'b00000000010000010000000100010011;
ROM[11152] <= 32'b00000001010000000000001110010011;
ROM[11153] <= 32'b00000000100000111000001110010011;
ROM[11154] <= 32'b01000000011100010000001110110011;
ROM[11155] <= 32'b00000000011100000000001000110011;
ROM[11156] <= 32'b00000000001000000000000110110011;
ROM[11157] <= 32'b01010101100100011110000011101111;
ROM[11158] <= 32'b00000110010100000000001110010011;
ROM[11159] <= 32'b00000000011100010010000000100011;
ROM[11160] <= 32'b00000000010000010000000100010011;
ROM[11161] <= 32'b00000000000000001011001110110111;
ROM[11162] <= 32'b11101011000000111000001110010011;
ROM[11163] <= 32'b00000000111000111000001110110011;
ROM[11164] <= 32'b00000000011100010010000000100011;
ROM[11165] <= 32'b00000000010000010000000100010011;
ROM[11166] <= 32'b00000000001100010010000000100011;
ROM[11167] <= 32'b00000000010000010000000100010011;
ROM[11168] <= 32'b00000000010000010010000000100011;
ROM[11169] <= 32'b00000000010000010000000100010011;
ROM[11170] <= 32'b00000000010100010010000000100011;
ROM[11171] <= 32'b00000000010000010000000100010011;
ROM[11172] <= 32'b00000000011000010010000000100011;
ROM[11173] <= 32'b00000000010000010000000100010011;
ROM[11174] <= 32'b00000001010000000000001110010011;
ROM[11175] <= 32'b00000000100000111000001110010011;
ROM[11176] <= 32'b01000000011100010000001110110011;
ROM[11177] <= 32'b00000000011100000000001000110011;
ROM[11178] <= 32'b00000000001000000000000110110011;
ROM[11179] <= 32'b01010000000100011110000011101111;
ROM[11180] <= 32'b00000010000000000000001110010011;
ROM[11181] <= 32'b00000000011100010010000000100011;
ROM[11182] <= 32'b00000000010000010000000100010011;
ROM[11183] <= 32'b00000000000000001011001110110111;
ROM[11184] <= 32'b11110000100000111000001110010011;
ROM[11185] <= 32'b00000000111000111000001110110011;
ROM[11186] <= 32'b00000000011100010010000000100011;
ROM[11187] <= 32'b00000000010000010000000100010011;
ROM[11188] <= 32'b00000000001100010010000000100011;
ROM[11189] <= 32'b00000000010000010000000100010011;
ROM[11190] <= 32'b00000000010000010010000000100011;
ROM[11191] <= 32'b00000000010000010000000100010011;
ROM[11192] <= 32'b00000000010100010010000000100011;
ROM[11193] <= 32'b00000000010000010000000100010011;
ROM[11194] <= 32'b00000000011000010010000000100011;
ROM[11195] <= 32'b00000000010000010000000100010011;
ROM[11196] <= 32'b00000001010000000000001110010011;
ROM[11197] <= 32'b00000000100000111000001110010011;
ROM[11198] <= 32'b01000000011100010000001110110011;
ROM[11199] <= 32'b00000000011100000000001000110011;
ROM[11200] <= 32'b00000000001000000000000110110011;
ROM[11201] <= 32'b01001010100100011110000011101111;
ROM[11202] <= 32'b00000000000000001011001110110111;
ROM[11203] <= 32'b11110101010000111000001110010011;
ROM[11204] <= 32'b00000000111000111000001110110011;
ROM[11205] <= 32'b00000000011100010010000000100011;
ROM[11206] <= 32'b00000000010000010000000100010011;
ROM[11207] <= 32'b00000000001100010010000000100011;
ROM[11208] <= 32'b00000000010000010000000100010011;
ROM[11209] <= 32'b00000000010000010010000000100011;
ROM[11210] <= 32'b00000000010000010000000100010011;
ROM[11211] <= 32'b00000000010100010010000000100011;
ROM[11212] <= 32'b00000000010000010000000100010011;
ROM[11213] <= 32'b00000000011000010010000000100011;
ROM[11214] <= 32'b00000000010000010000000100010011;
ROM[11215] <= 32'b00000001010000000000001110010011;
ROM[11216] <= 32'b00000000010000111000001110010011;
ROM[11217] <= 32'b01000000011100010000001110110011;
ROM[11218] <= 32'b00000000011100000000001000110011;
ROM[11219] <= 32'b00000000001000000000000110110011;
ROM[11220] <= 32'b00000001100000001100000011101111;
ROM[11221] <= 32'b11111111110000010000000100010011;
ROM[11222] <= 32'b00000000000000010010001110000011;
ROM[11223] <= 32'b00000000011101100010000000100011;
ROM[11224] <= 32'b00000001010000011010001110000011;
ROM[11225] <= 32'b00000000011100010010000000100011;
ROM[11226] <= 32'b00000000010000010000000100010011;
ROM[11227] <= 32'b00000000000000001011001110110111;
ROM[11228] <= 32'b11111011100000111000001110010011;
ROM[11229] <= 32'b00000000111000111000001110110011;
ROM[11230] <= 32'b00000000011100010010000000100011;
ROM[11231] <= 32'b00000000010000010000000100010011;
ROM[11232] <= 32'b00000000001100010010000000100011;
ROM[11233] <= 32'b00000000010000010000000100010011;
ROM[11234] <= 32'b00000000010000010010000000100011;
ROM[11235] <= 32'b00000000010000010000000100010011;
ROM[11236] <= 32'b00000000010100010010000000100011;
ROM[11237] <= 32'b00000000010000010000000100010011;
ROM[11238] <= 32'b00000000011000010010000000100011;
ROM[11239] <= 32'b00000000010000010000000100010011;
ROM[11240] <= 32'b00000001010000000000001110010011;
ROM[11241] <= 32'b00000000010000111000001110010011;
ROM[11242] <= 32'b01000000011100010000001110110011;
ROM[11243] <= 32'b00000000011100000000001000110011;
ROM[11244] <= 32'b00000000001000000000000110110011;
ROM[11245] <= 32'b00011100110000001100000011101111;
ROM[11246] <= 32'b11111111110000010000000100010011;
ROM[11247] <= 32'b00000000000000010010001110000011;
ROM[11248] <= 32'b00000000011101100010000000100011;
ROM[11249] <= 32'b00000001001100000000001110010011;
ROM[11250] <= 32'b00000000011100010010000000100011;
ROM[11251] <= 32'b00000000010000010000000100010011;
ROM[11252] <= 32'b00000000000000001011001110110111;
ROM[11253] <= 32'b00000001110000111000001110010011;
ROM[11254] <= 32'b00000000111000111000001110110011;
ROM[11255] <= 32'b00000000011100010010000000100011;
ROM[11256] <= 32'b00000000010000010000000100010011;
ROM[11257] <= 32'b00000000001100010010000000100011;
ROM[11258] <= 32'b00000000010000010000000100010011;
ROM[11259] <= 32'b00000000010000010010000000100011;
ROM[11260] <= 32'b00000000010000010000000100010011;
ROM[11261] <= 32'b00000000010100010010000000100011;
ROM[11262] <= 32'b00000000010000010000000100010011;
ROM[11263] <= 32'b00000000011000010010000000100011;
ROM[11264] <= 32'b00000000010000010000000100010011;
ROM[11265] <= 32'b00000001010000000000001110010011;
ROM[11266] <= 32'b00000000010000111000001110010011;
ROM[11267] <= 32'b01000000011100010000001110110011;
ROM[11268] <= 32'b00000000011100000000001000110011;
ROM[11269] <= 32'b00000000001000000000000110110011;
ROM[11270] <= 32'b01110010010000011110000011101111;
ROM[11271] <= 32'b00000010000000000000001110010011;
ROM[11272] <= 32'b00000000011100010010000000100011;
ROM[11273] <= 32'b00000000010000010000000100010011;
ROM[11274] <= 32'b00000000000000001011001110110111;
ROM[11275] <= 32'b00000111010000111000001110010011;
ROM[11276] <= 32'b00000000111000111000001110110011;
ROM[11277] <= 32'b00000000011100010010000000100011;
ROM[11278] <= 32'b00000000010000010000000100010011;
ROM[11279] <= 32'b00000000001100010010000000100011;
ROM[11280] <= 32'b00000000010000010000000100010011;
ROM[11281] <= 32'b00000000010000010010000000100011;
ROM[11282] <= 32'b00000000010000010000000100010011;
ROM[11283] <= 32'b00000000010100010010000000100011;
ROM[11284] <= 32'b00000000010000010000000100010011;
ROM[11285] <= 32'b00000000011000010010000000100011;
ROM[11286] <= 32'b00000000010000010000000100010011;
ROM[11287] <= 32'b00000001010000000000001110010011;
ROM[11288] <= 32'b00000000100000111000001110010011;
ROM[11289] <= 32'b01000000011100010000001110110011;
ROM[11290] <= 32'b00000000011100000000001000110011;
ROM[11291] <= 32'b00000000001000000000000110110011;
ROM[11292] <= 32'b00110011110100011110000011101111;
ROM[11293] <= 32'b00000110000100000000001110010011;
ROM[11294] <= 32'b00000000011100010010000000100011;
ROM[11295] <= 32'b00000000010000010000000100010011;
ROM[11296] <= 32'b00000000000000001011001110110111;
ROM[11297] <= 32'b00001100110000111000001110010011;
ROM[11298] <= 32'b00000000111000111000001110110011;
ROM[11299] <= 32'b00000000011100010010000000100011;
ROM[11300] <= 32'b00000000010000010000000100010011;
ROM[11301] <= 32'b00000000001100010010000000100011;
ROM[11302] <= 32'b00000000010000010000000100010011;
ROM[11303] <= 32'b00000000010000010010000000100011;
ROM[11304] <= 32'b00000000010000010000000100010011;
ROM[11305] <= 32'b00000000010100010010000000100011;
ROM[11306] <= 32'b00000000010000010000000100010011;
ROM[11307] <= 32'b00000000011000010010000000100011;
ROM[11308] <= 32'b00000000010000010000000100010011;
ROM[11309] <= 32'b00000001010000000000001110010011;
ROM[11310] <= 32'b00000000100000111000001110010011;
ROM[11311] <= 32'b01000000011100010000001110110011;
ROM[11312] <= 32'b00000000011100000000001000110011;
ROM[11313] <= 32'b00000000001000000000000110110011;
ROM[11314] <= 32'b00101110010100011110000011101111;
ROM[11315] <= 32'b00000111010000000000001110010011;
ROM[11316] <= 32'b00000000011100010010000000100011;
ROM[11317] <= 32'b00000000010000010000000100010011;
ROM[11318] <= 32'b00000000000000001011001110110111;
ROM[11319] <= 32'b00010010010000111000001110010011;
ROM[11320] <= 32'b00000000111000111000001110110011;
ROM[11321] <= 32'b00000000011100010010000000100011;
ROM[11322] <= 32'b00000000010000010000000100010011;
ROM[11323] <= 32'b00000000001100010010000000100011;
ROM[11324] <= 32'b00000000010000010000000100010011;
ROM[11325] <= 32'b00000000010000010010000000100011;
ROM[11326] <= 32'b00000000010000010000000100010011;
ROM[11327] <= 32'b00000000010100010010000000100011;
ROM[11328] <= 32'b00000000010000010000000100010011;
ROM[11329] <= 32'b00000000011000010010000000100011;
ROM[11330] <= 32'b00000000010000010000000100010011;
ROM[11331] <= 32'b00000001010000000000001110010011;
ROM[11332] <= 32'b00000000100000111000001110010011;
ROM[11333] <= 32'b01000000011100010000001110110011;
ROM[11334] <= 32'b00000000011100000000001000110011;
ROM[11335] <= 32'b00000000001000000000000110110011;
ROM[11336] <= 32'b00101000110100011110000011101111;
ROM[11337] <= 32'b00000111010000000000001110010011;
ROM[11338] <= 32'b00000000011100010010000000100011;
ROM[11339] <= 32'b00000000010000010000000100010011;
ROM[11340] <= 32'b00000000000000001011001110110111;
ROM[11341] <= 32'b00010111110000111000001110010011;
ROM[11342] <= 32'b00000000111000111000001110110011;
ROM[11343] <= 32'b00000000011100010010000000100011;
ROM[11344] <= 32'b00000000010000010000000100010011;
ROM[11345] <= 32'b00000000001100010010000000100011;
ROM[11346] <= 32'b00000000010000010000000100010011;
ROM[11347] <= 32'b00000000010000010010000000100011;
ROM[11348] <= 32'b00000000010000010000000100010011;
ROM[11349] <= 32'b00000000010100010010000000100011;
ROM[11350] <= 32'b00000000010000010000000100010011;
ROM[11351] <= 32'b00000000011000010010000000100011;
ROM[11352] <= 32'b00000000010000010000000100010011;
ROM[11353] <= 32'b00000001010000000000001110010011;
ROM[11354] <= 32'b00000000100000111000001110010011;
ROM[11355] <= 32'b01000000011100010000001110110011;
ROM[11356] <= 32'b00000000011100000000001000110011;
ROM[11357] <= 32'b00000000001000000000000110110011;
ROM[11358] <= 32'b00100011010100011110000011101111;
ROM[11359] <= 32'b00000110010100000000001110010011;
ROM[11360] <= 32'b00000000011100010010000000100011;
ROM[11361] <= 32'b00000000010000010000000100010011;
ROM[11362] <= 32'b00000000000000001011001110110111;
ROM[11363] <= 32'b00011101010000111000001110010011;
ROM[11364] <= 32'b00000000111000111000001110110011;
ROM[11365] <= 32'b00000000011100010010000000100011;
ROM[11366] <= 32'b00000000010000010000000100010011;
ROM[11367] <= 32'b00000000001100010010000000100011;
ROM[11368] <= 32'b00000000010000010000000100010011;
ROM[11369] <= 32'b00000000010000010010000000100011;
ROM[11370] <= 32'b00000000010000010000000100010011;
ROM[11371] <= 32'b00000000010100010010000000100011;
ROM[11372] <= 32'b00000000010000010000000100010011;
ROM[11373] <= 32'b00000000011000010010000000100011;
ROM[11374] <= 32'b00000000010000010000000100010011;
ROM[11375] <= 32'b00000001010000000000001110010011;
ROM[11376] <= 32'b00000000100000111000001110010011;
ROM[11377] <= 32'b01000000011100010000001110110011;
ROM[11378] <= 32'b00000000011100000000001000110011;
ROM[11379] <= 32'b00000000001000000000000110110011;
ROM[11380] <= 32'b00011101110100011110000011101111;
ROM[11381] <= 32'b00000110110100000000001110010011;
ROM[11382] <= 32'b00000000011100010010000000100011;
ROM[11383] <= 32'b00000000010000010000000100010011;
ROM[11384] <= 32'b00000000000000001011001110110111;
ROM[11385] <= 32'b00100010110000111000001110010011;
ROM[11386] <= 32'b00000000111000111000001110110011;
ROM[11387] <= 32'b00000000011100010010000000100011;
ROM[11388] <= 32'b00000000010000010000000100010011;
ROM[11389] <= 32'b00000000001100010010000000100011;
ROM[11390] <= 32'b00000000010000010000000100010011;
ROM[11391] <= 32'b00000000010000010010000000100011;
ROM[11392] <= 32'b00000000010000010000000100010011;
ROM[11393] <= 32'b00000000010100010010000000100011;
ROM[11394] <= 32'b00000000010000010000000100010011;
ROM[11395] <= 32'b00000000011000010010000000100011;
ROM[11396] <= 32'b00000000010000010000000100010011;
ROM[11397] <= 32'b00000001010000000000001110010011;
ROM[11398] <= 32'b00000000100000111000001110010011;
ROM[11399] <= 32'b01000000011100010000001110110011;
ROM[11400] <= 32'b00000000011100000000001000110011;
ROM[11401] <= 32'b00000000001000000000000110110011;
ROM[11402] <= 32'b00011000010100011110000011101111;
ROM[11403] <= 32'b00000111000000000000001110010011;
ROM[11404] <= 32'b00000000011100010010000000100011;
ROM[11405] <= 32'b00000000010000010000000100010011;
ROM[11406] <= 32'b00000000000000001011001110110111;
ROM[11407] <= 32'b00101000010000111000001110010011;
ROM[11408] <= 32'b00000000111000111000001110110011;
ROM[11409] <= 32'b00000000011100010010000000100011;
ROM[11410] <= 32'b00000000010000010000000100010011;
ROM[11411] <= 32'b00000000001100010010000000100011;
ROM[11412] <= 32'b00000000010000010000000100010011;
ROM[11413] <= 32'b00000000010000010010000000100011;
ROM[11414] <= 32'b00000000010000010000000100010011;
ROM[11415] <= 32'b00000000010100010010000000100011;
ROM[11416] <= 32'b00000000010000010000000100010011;
ROM[11417] <= 32'b00000000011000010010000000100011;
ROM[11418] <= 32'b00000000010000010000000100010011;
ROM[11419] <= 32'b00000001010000000000001110010011;
ROM[11420] <= 32'b00000000100000111000001110010011;
ROM[11421] <= 32'b01000000011100010000001110110011;
ROM[11422] <= 32'b00000000011100000000001000110011;
ROM[11423] <= 32'b00000000001000000000000110110011;
ROM[11424] <= 32'b00010010110100011110000011101111;
ROM[11425] <= 32'b00000111010000000000001110010011;
ROM[11426] <= 32'b00000000011100010010000000100011;
ROM[11427] <= 32'b00000000010000010000000100010011;
ROM[11428] <= 32'b00000000000000001011001110110111;
ROM[11429] <= 32'b00101101110000111000001110010011;
ROM[11430] <= 32'b00000000111000111000001110110011;
ROM[11431] <= 32'b00000000011100010010000000100011;
ROM[11432] <= 32'b00000000010000010000000100010011;
ROM[11433] <= 32'b00000000001100010010000000100011;
ROM[11434] <= 32'b00000000010000010000000100010011;
ROM[11435] <= 32'b00000000010000010010000000100011;
ROM[11436] <= 32'b00000000010000010000000100010011;
ROM[11437] <= 32'b00000000010100010010000000100011;
ROM[11438] <= 32'b00000000010000010000000100010011;
ROM[11439] <= 32'b00000000011000010010000000100011;
ROM[11440] <= 32'b00000000010000010000000100010011;
ROM[11441] <= 32'b00000001010000000000001110010011;
ROM[11442] <= 32'b00000000100000111000001110010011;
ROM[11443] <= 32'b01000000011100010000001110110011;
ROM[11444] <= 32'b00000000011100000000001000110011;
ROM[11445] <= 32'b00000000001000000000000110110011;
ROM[11446] <= 32'b00001101010100011110000011101111;
ROM[11447] <= 32'b00000111001100000000001110010011;
ROM[11448] <= 32'b00000000011100010010000000100011;
ROM[11449] <= 32'b00000000010000010000000100010011;
ROM[11450] <= 32'b00000000000000001011001110110111;
ROM[11451] <= 32'b00110011010000111000001110010011;
ROM[11452] <= 32'b00000000111000111000001110110011;
ROM[11453] <= 32'b00000000011100010010000000100011;
ROM[11454] <= 32'b00000000010000010000000100010011;
ROM[11455] <= 32'b00000000001100010010000000100011;
ROM[11456] <= 32'b00000000010000010000000100010011;
ROM[11457] <= 32'b00000000010000010010000000100011;
ROM[11458] <= 32'b00000000010000010000000100010011;
ROM[11459] <= 32'b00000000010100010010000000100011;
ROM[11460] <= 32'b00000000010000010000000100010011;
ROM[11461] <= 32'b00000000011000010010000000100011;
ROM[11462] <= 32'b00000000010000010000000100010011;
ROM[11463] <= 32'b00000001010000000000001110010011;
ROM[11464] <= 32'b00000000100000111000001110010011;
ROM[11465] <= 32'b01000000011100010000001110110011;
ROM[11466] <= 32'b00000000011100000000001000110011;
ROM[11467] <= 32'b00000000001000000000000110110011;
ROM[11468] <= 32'b00000111110100011110000011101111;
ROM[11469] <= 32'b00000010000000000000001110010011;
ROM[11470] <= 32'b00000000011100010010000000100011;
ROM[11471] <= 32'b00000000010000010000000100010011;
ROM[11472] <= 32'b00000000000000001011001110110111;
ROM[11473] <= 32'b00111000110000111000001110010011;
ROM[11474] <= 32'b00000000111000111000001110110011;
ROM[11475] <= 32'b00000000011100010010000000100011;
ROM[11476] <= 32'b00000000010000010000000100010011;
ROM[11477] <= 32'b00000000001100010010000000100011;
ROM[11478] <= 32'b00000000010000010000000100010011;
ROM[11479] <= 32'b00000000010000010010000000100011;
ROM[11480] <= 32'b00000000010000010000000100010011;
ROM[11481] <= 32'b00000000010100010010000000100011;
ROM[11482] <= 32'b00000000010000010000000100010011;
ROM[11483] <= 32'b00000000011000010010000000100011;
ROM[11484] <= 32'b00000000010000010000000100010011;
ROM[11485] <= 32'b00000001010000000000001110010011;
ROM[11486] <= 32'b00000000100000111000001110010011;
ROM[11487] <= 32'b01000000011100010000001110110011;
ROM[11488] <= 32'b00000000011100000000001000110011;
ROM[11489] <= 32'b00000000001000000000000110110011;
ROM[11490] <= 32'b00000010010100011110000011101111;
ROM[11491] <= 32'b00000111001000000000001110010011;
ROM[11492] <= 32'b00000000011100010010000000100011;
ROM[11493] <= 32'b00000000010000010000000100010011;
ROM[11494] <= 32'b00000000000000001011001110110111;
ROM[11495] <= 32'b00111110010000111000001110010011;
ROM[11496] <= 32'b00000000111000111000001110110011;
ROM[11497] <= 32'b00000000011100010010000000100011;
ROM[11498] <= 32'b00000000010000010000000100010011;
ROM[11499] <= 32'b00000000001100010010000000100011;
ROM[11500] <= 32'b00000000010000010000000100010011;
ROM[11501] <= 32'b00000000010000010010000000100011;
ROM[11502] <= 32'b00000000010000010000000100010011;
ROM[11503] <= 32'b00000000010100010010000000100011;
ROM[11504] <= 32'b00000000010000010000000100010011;
ROM[11505] <= 32'b00000000011000010010000000100011;
ROM[11506] <= 32'b00000000010000010000000100010011;
ROM[11507] <= 32'b00000001010000000000001110010011;
ROM[11508] <= 32'b00000000100000111000001110010011;
ROM[11509] <= 32'b01000000011100010000001110110011;
ROM[11510] <= 32'b00000000011100000000001000110011;
ROM[11511] <= 32'b00000000001000000000000110110011;
ROM[11512] <= 32'b01111100110000011110000011101111;
ROM[11513] <= 32'b00000110010100000000001110010011;
ROM[11514] <= 32'b00000000011100010010000000100011;
ROM[11515] <= 32'b00000000010000010000000100010011;
ROM[11516] <= 32'b00000000000000001011001110110111;
ROM[11517] <= 32'b01000011110000111000001110010011;
ROM[11518] <= 32'b00000000111000111000001110110011;
ROM[11519] <= 32'b00000000011100010010000000100011;
ROM[11520] <= 32'b00000000010000010000000100010011;
ROM[11521] <= 32'b00000000001100010010000000100011;
ROM[11522] <= 32'b00000000010000010000000100010011;
ROM[11523] <= 32'b00000000010000010010000000100011;
ROM[11524] <= 32'b00000000010000010000000100010011;
ROM[11525] <= 32'b00000000010100010010000000100011;
ROM[11526] <= 32'b00000000010000010000000100010011;
ROM[11527] <= 32'b00000000011000010010000000100011;
ROM[11528] <= 32'b00000000010000010000000100010011;
ROM[11529] <= 32'b00000001010000000000001110010011;
ROM[11530] <= 32'b00000000100000111000001110010011;
ROM[11531] <= 32'b01000000011100010000001110110011;
ROM[11532] <= 32'b00000000011100000000001000110011;
ROM[11533] <= 32'b00000000001000000000000110110011;
ROM[11534] <= 32'b01110111010000011110000011101111;
ROM[11535] <= 32'b00000110110100000000001110010011;
ROM[11536] <= 32'b00000000011100010010000000100011;
ROM[11537] <= 32'b00000000010000010000000100010011;
ROM[11538] <= 32'b00000000000000001011001110110111;
ROM[11539] <= 32'b01001001010000111000001110010011;
ROM[11540] <= 32'b00000000111000111000001110110011;
ROM[11541] <= 32'b00000000011100010010000000100011;
ROM[11542] <= 32'b00000000010000010000000100010011;
ROM[11543] <= 32'b00000000001100010010000000100011;
ROM[11544] <= 32'b00000000010000010000000100010011;
ROM[11545] <= 32'b00000000010000010010000000100011;
ROM[11546] <= 32'b00000000010000010000000100010011;
ROM[11547] <= 32'b00000000010100010010000000100011;
ROM[11548] <= 32'b00000000010000010000000100010011;
ROM[11549] <= 32'b00000000011000010010000000100011;
ROM[11550] <= 32'b00000000010000010000000100010011;
ROM[11551] <= 32'b00000001010000000000001110010011;
ROM[11552] <= 32'b00000000100000111000001110010011;
ROM[11553] <= 32'b01000000011100010000001110110011;
ROM[11554] <= 32'b00000000011100000000001000110011;
ROM[11555] <= 32'b00000000001000000000000110110011;
ROM[11556] <= 32'b01110001110000011110000011101111;
ROM[11557] <= 32'b00000110000100000000001110010011;
ROM[11558] <= 32'b00000000011100010010000000100011;
ROM[11559] <= 32'b00000000010000010000000100010011;
ROM[11560] <= 32'b00000000000000001011001110110111;
ROM[11561] <= 32'b01001110110000111000001110010011;
ROM[11562] <= 32'b00000000111000111000001110110011;
ROM[11563] <= 32'b00000000011100010010000000100011;
ROM[11564] <= 32'b00000000010000010000000100010011;
ROM[11565] <= 32'b00000000001100010010000000100011;
ROM[11566] <= 32'b00000000010000010000000100010011;
ROM[11567] <= 32'b00000000010000010010000000100011;
ROM[11568] <= 32'b00000000010000010000000100010011;
ROM[11569] <= 32'b00000000010100010010000000100011;
ROM[11570] <= 32'b00000000010000010000000100010011;
ROM[11571] <= 32'b00000000011000010010000000100011;
ROM[11572] <= 32'b00000000010000010000000100010011;
ROM[11573] <= 32'b00000001010000000000001110010011;
ROM[11574] <= 32'b00000000100000111000001110010011;
ROM[11575] <= 32'b01000000011100010000001110110011;
ROM[11576] <= 32'b00000000011100000000001000110011;
ROM[11577] <= 32'b00000000001000000000000110110011;
ROM[11578] <= 32'b01101100010000011110000011101111;
ROM[11579] <= 32'b00000110100100000000001110010011;
ROM[11580] <= 32'b00000000011100010010000000100011;
ROM[11581] <= 32'b00000000010000010000000100010011;
ROM[11582] <= 32'b00000000000000001011001110110111;
ROM[11583] <= 32'b01010100010000111000001110010011;
ROM[11584] <= 32'b00000000111000111000001110110011;
ROM[11585] <= 32'b00000000011100010010000000100011;
ROM[11586] <= 32'b00000000010000010000000100010011;
ROM[11587] <= 32'b00000000001100010010000000100011;
ROM[11588] <= 32'b00000000010000010000000100010011;
ROM[11589] <= 32'b00000000010000010010000000100011;
ROM[11590] <= 32'b00000000010000010000000100010011;
ROM[11591] <= 32'b00000000010100010010000000100011;
ROM[11592] <= 32'b00000000010000010000000100010011;
ROM[11593] <= 32'b00000000011000010010000000100011;
ROM[11594] <= 32'b00000000010000010000000100010011;
ROM[11595] <= 32'b00000001010000000000001110010011;
ROM[11596] <= 32'b00000000100000111000001110010011;
ROM[11597] <= 32'b01000000011100010000001110110011;
ROM[11598] <= 32'b00000000011100000000001000110011;
ROM[11599] <= 32'b00000000001000000000000110110011;
ROM[11600] <= 32'b01100110110000011110000011101111;
ROM[11601] <= 32'b00000110111000000000001110010011;
ROM[11602] <= 32'b00000000011100010010000000100011;
ROM[11603] <= 32'b00000000010000010000000100010011;
ROM[11604] <= 32'b00000000000000001011001110110111;
ROM[11605] <= 32'b01011001110000111000001110010011;
ROM[11606] <= 32'b00000000111000111000001110110011;
ROM[11607] <= 32'b00000000011100010010000000100011;
ROM[11608] <= 32'b00000000010000010000000100010011;
ROM[11609] <= 32'b00000000001100010010000000100011;
ROM[11610] <= 32'b00000000010000010000000100010011;
ROM[11611] <= 32'b00000000010000010010000000100011;
ROM[11612] <= 32'b00000000010000010000000100010011;
ROM[11613] <= 32'b00000000010100010010000000100011;
ROM[11614] <= 32'b00000000010000010000000100010011;
ROM[11615] <= 32'b00000000011000010010000000100011;
ROM[11616] <= 32'b00000000010000010000000100010011;
ROM[11617] <= 32'b00000001010000000000001110010011;
ROM[11618] <= 32'b00000000100000111000001110010011;
ROM[11619] <= 32'b01000000011100010000001110110011;
ROM[11620] <= 32'b00000000011100000000001000110011;
ROM[11621] <= 32'b00000000001000000000000110110011;
ROM[11622] <= 32'b01100001010000011110000011101111;
ROM[11623] <= 32'b00000110100100000000001110010011;
ROM[11624] <= 32'b00000000011100010010000000100011;
ROM[11625] <= 32'b00000000010000010000000100010011;
ROM[11626] <= 32'b00000000000000001011001110110111;
ROM[11627] <= 32'b01011111010000111000001110010011;
ROM[11628] <= 32'b00000000111000111000001110110011;
ROM[11629] <= 32'b00000000011100010010000000100011;
ROM[11630] <= 32'b00000000010000010000000100010011;
ROM[11631] <= 32'b00000000001100010010000000100011;
ROM[11632] <= 32'b00000000010000010000000100010011;
ROM[11633] <= 32'b00000000010000010010000000100011;
ROM[11634] <= 32'b00000000010000010000000100010011;
ROM[11635] <= 32'b00000000010100010010000000100011;
ROM[11636] <= 32'b00000000010000010000000100010011;
ROM[11637] <= 32'b00000000011000010010000000100011;
ROM[11638] <= 32'b00000000010000010000000100010011;
ROM[11639] <= 32'b00000001010000000000001110010011;
ROM[11640] <= 32'b00000000100000111000001110010011;
ROM[11641] <= 32'b01000000011100010000001110110011;
ROM[11642] <= 32'b00000000011100000000001000110011;
ROM[11643] <= 32'b00000000001000000000000110110011;
ROM[11644] <= 32'b01011011110000011110000011101111;
ROM[11645] <= 32'b00000110111000000000001110010011;
ROM[11646] <= 32'b00000000011100010010000000100011;
ROM[11647] <= 32'b00000000010000010000000100010011;
ROM[11648] <= 32'b00000000000000001011001110110111;
ROM[11649] <= 32'b01100100110000111000001110010011;
ROM[11650] <= 32'b00000000111000111000001110110011;
ROM[11651] <= 32'b00000000011100010010000000100011;
ROM[11652] <= 32'b00000000010000010000000100010011;
ROM[11653] <= 32'b00000000001100010010000000100011;
ROM[11654] <= 32'b00000000010000010000000100010011;
ROM[11655] <= 32'b00000000010000010010000000100011;
ROM[11656] <= 32'b00000000010000010000000100010011;
ROM[11657] <= 32'b00000000010100010010000000100011;
ROM[11658] <= 32'b00000000010000010000000100010011;
ROM[11659] <= 32'b00000000011000010010000000100011;
ROM[11660] <= 32'b00000000010000010000000100010011;
ROM[11661] <= 32'b00000001010000000000001110010011;
ROM[11662] <= 32'b00000000100000111000001110010011;
ROM[11663] <= 32'b01000000011100010000001110110011;
ROM[11664] <= 32'b00000000011100000000001000110011;
ROM[11665] <= 32'b00000000001000000000000110110011;
ROM[11666] <= 32'b01010110010000011110000011101111;
ROM[11667] <= 32'b00000110011100000000001110010011;
ROM[11668] <= 32'b00000000011100010010000000100011;
ROM[11669] <= 32'b00000000010000010000000100010011;
ROM[11670] <= 32'b00000000000000001011001110110111;
ROM[11671] <= 32'b01101010010000111000001110010011;
ROM[11672] <= 32'b00000000111000111000001110110011;
ROM[11673] <= 32'b00000000011100010010000000100011;
ROM[11674] <= 32'b00000000010000010000000100010011;
ROM[11675] <= 32'b00000000001100010010000000100011;
ROM[11676] <= 32'b00000000010000010000000100010011;
ROM[11677] <= 32'b00000000010000010010000000100011;
ROM[11678] <= 32'b00000000010000010000000100010011;
ROM[11679] <= 32'b00000000010100010010000000100011;
ROM[11680] <= 32'b00000000010000010000000100010011;
ROM[11681] <= 32'b00000000011000010010000000100011;
ROM[11682] <= 32'b00000000010000010000000100010011;
ROM[11683] <= 32'b00000001010000000000001110010011;
ROM[11684] <= 32'b00000000100000111000001110010011;
ROM[11685] <= 32'b01000000011100010000001110110011;
ROM[11686] <= 32'b00000000011100000000001000110011;
ROM[11687] <= 32'b00000000001000000000000110110011;
ROM[11688] <= 32'b01010000110000011110000011101111;
ROM[11689] <= 32'b00000000000000001011001110110111;
ROM[11690] <= 32'b01101111000000111000001110010011;
ROM[11691] <= 32'b00000000111000111000001110110011;
ROM[11692] <= 32'b00000000011100010010000000100011;
ROM[11693] <= 32'b00000000010000010000000100010011;
ROM[11694] <= 32'b00000000001100010010000000100011;
ROM[11695] <= 32'b00000000010000010000000100010011;
ROM[11696] <= 32'b00000000010000010010000000100011;
ROM[11697] <= 32'b00000000010000010000000100010011;
ROM[11698] <= 32'b00000000010100010010000000100011;
ROM[11699] <= 32'b00000000010000010000000100010011;
ROM[11700] <= 32'b00000000011000010010000000100011;
ROM[11701] <= 32'b00000000010000010000000100010011;
ROM[11702] <= 32'b00000001010000000000001110010011;
ROM[11703] <= 32'b00000000010000111000001110010011;
ROM[11704] <= 32'b01000000011100010000001110110011;
ROM[11705] <= 32'b00000000011100000000001000110011;
ROM[11706] <= 32'b00000000001000000000000110110011;
ROM[11707] <= 32'b00000111110100001011000011101111;
ROM[11708] <= 32'b11111111110000010000000100010011;
ROM[11709] <= 32'b00000000000000010010001110000011;
ROM[11710] <= 32'b00000000011101100010000000100011;
ROM[11711] <= 32'b00000000000000001011001110110111;
ROM[11712] <= 32'b01110100100000111000001110010011;
ROM[11713] <= 32'b00000000111000111000001110110011;
ROM[11714] <= 32'b00000000011100010010000000100011;
ROM[11715] <= 32'b00000000010000010000000100010011;
ROM[11716] <= 32'b00000000001100010010000000100011;
ROM[11717] <= 32'b00000000010000010000000100010011;
ROM[11718] <= 32'b00000000010000010010000000100011;
ROM[11719] <= 32'b00000000010000010000000100010011;
ROM[11720] <= 32'b00000000010100010010000000100011;
ROM[11721] <= 32'b00000000010000010000000100010011;
ROM[11722] <= 32'b00000000011000010010000000100011;
ROM[11723] <= 32'b00000000010000010000000100010011;
ROM[11724] <= 32'b00000001010000000000001110010011;
ROM[11725] <= 32'b00000000000000111000001110010011;
ROM[11726] <= 32'b01000000011100010000001110110011;
ROM[11727] <= 32'b00000000011100000000001000110011;
ROM[11728] <= 32'b00000000001000000000000110110011;
ROM[11729] <= 32'b01000010010100001011000011101111;
ROM[11730] <= 32'b11111111110000010000000100010011;
ROM[11731] <= 32'b00000000000000010010001110000011;
ROM[11732] <= 32'b00000000011101100010000000100011;
ROM[11733] <= 32'b01101100010100000000000011101111;
ROM[11734] <= 32'b00000001011100000000001110010011;
ROM[11735] <= 32'b00000000011100010010000000100011;
ROM[11736] <= 32'b00000000010000010000000100010011;
ROM[11737] <= 32'b00000000000000001011001110110111;
ROM[11738] <= 32'b01111011000000111000001110010011;
ROM[11739] <= 32'b00000000111000111000001110110011;
ROM[11740] <= 32'b00000000011100010010000000100011;
ROM[11741] <= 32'b00000000010000010000000100010011;
ROM[11742] <= 32'b00000000001100010010000000100011;
ROM[11743] <= 32'b00000000010000010000000100010011;
ROM[11744] <= 32'b00000000010000010010000000100011;
ROM[11745] <= 32'b00000000010000010000000100010011;
ROM[11746] <= 32'b00000000010100010010000000100011;
ROM[11747] <= 32'b00000000010000010000000100010011;
ROM[11748] <= 32'b00000000011000010010000000100011;
ROM[11749] <= 32'b00000000010000010000000100010011;
ROM[11750] <= 32'b00000001010000000000001110010011;
ROM[11751] <= 32'b00000000010000111000001110010011;
ROM[11752] <= 32'b01000000011100010000001110110011;
ROM[11753] <= 32'b00000000011100000000001000110011;
ROM[11754] <= 32'b00000000001000000000000110110011;
ROM[11755] <= 32'b01111001000100011101000011101111;
ROM[11756] <= 32'b00000101011100000000001110010011;
ROM[11757] <= 32'b00000000011100010010000000100011;
ROM[11758] <= 32'b00000000010000010000000100010011;
ROM[11759] <= 32'b00000000000000001100001110110111;
ROM[11760] <= 32'b10000000100000111000001110010011;
ROM[11761] <= 32'b00000000111000111000001110110011;
ROM[11762] <= 32'b00000000011100010010000000100011;
ROM[11763] <= 32'b00000000010000010000000100010011;
ROM[11764] <= 32'b00000000001100010010000000100011;
ROM[11765] <= 32'b00000000010000010000000100010011;
ROM[11766] <= 32'b00000000010000010010000000100011;
ROM[11767] <= 32'b00000000010000010000000100010011;
ROM[11768] <= 32'b00000000010100010010000000100011;
ROM[11769] <= 32'b00000000010000010000000100010011;
ROM[11770] <= 32'b00000000011000010010000000100011;
ROM[11771] <= 32'b00000000010000010000000100010011;
ROM[11772] <= 32'b00000001010000000000001110010011;
ROM[11773] <= 32'b00000000100000111000001110010011;
ROM[11774] <= 32'b01000000011100010000001110110011;
ROM[11775] <= 32'b00000000011100000000001000110011;
ROM[11776] <= 32'b00000000001000000000000110110011;
ROM[11777] <= 32'b00111010100000011110000011101111;
ROM[11778] <= 32'b00000111001000000000001110010011;
ROM[11779] <= 32'b00000000011100010010000000100011;
ROM[11780] <= 32'b00000000010000010000000100010011;
ROM[11781] <= 32'b00000000000000001100001110110111;
ROM[11782] <= 32'b10000110000000111000001110010011;
ROM[11783] <= 32'b00000000111000111000001110110011;
ROM[11784] <= 32'b00000000011100010010000000100011;
ROM[11785] <= 32'b00000000010000010000000100010011;
ROM[11786] <= 32'b00000000001100010010000000100011;
ROM[11787] <= 32'b00000000010000010000000100010011;
ROM[11788] <= 32'b00000000010000010010000000100011;
ROM[11789] <= 32'b00000000010000010000000100010011;
ROM[11790] <= 32'b00000000010100010010000000100011;
ROM[11791] <= 32'b00000000010000010000000100010011;
ROM[11792] <= 32'b00000000011000010010000000100011;
ROM[11793] <= 32'b00000000010000010000000100010011;
ROM[11794] <= 32'b00000001010000000000001110010011;
ROM[11795] <= 32'b00000000100000111000001110010011;
ROM[11796] <= 32'b01000000011100010000001110110011;
ROM[11797] <= 32'b00000000011100000000001000110011;
ROM[11798] <= 32'b00000000001000000000000110110011;
ROM[11799] <= 32'b00110101000000011110000011101111;
ROM[11800] <= 32'b00000110111100000000001110010011;
ROM[11801] <= 32'b00000000011100010010000000100011;
ROM[11802] <= 32'b00000000010000010000000100010011;
ROM[11803] <= 32'b00000000000000001100001110110111;
ROM[11804] <= 32'b10001011100000111000001110010011;
ROM[11805] <= 32'b00000000111000111000001110110011;
ROM[11806] <= 32'b00000000011100010010000000100011;
ROM[11807] <= 32'b00000000010000010000000100010011;
ROM[11808] <= 32'b00000000001100010010000000100011;
ROM[11809] <= 32'b00000000010000010000000100010011;
ROM[11810] <= 32'b00000000010000010010000000100011;
ROM[11811] <= 32'b00000000010000010000000100010011;
ROM[11812] <= 32'b00000000010100010010000000100011;
ROM[11813] <= 32'b00000000010000010000000100010011;
ROM[11814] <= 32'b00000000011000010010000000100011;
ROM[11815] <= 32'b00000000010000010000000100010011;
ROM[11816] <= 32'b00000001010000000000001110010011;
ROM[11817] <= 32'b00000000100000111000001110010011;
ROM[11818] <= 32'b01000000011100010000001110110011;
ROM[11819] <= 32'b00000000011100000000001000110011;
ROM[11820] <= 32'b00000000001000000000000110110011;
ROM[11821] <= 32'b00101111100000011110000011101111;
ROM[11822] <= 32'b00000110111000000000001110010011;
ROM[11823] <= 32'b00000000011100010010000000100011;
ROM[11824] <= 32'b00000000010000010000000100010011;
ROM[11825] <= 32'b00000000000000001100001110110111;
ROM[11826] <= 32'b10010001000000111000001110010011;
ROM[11827] <= 32'b00000000111000111000001110110011;
ROM[11828] <= 32'b00000000011100010010000000100011;
ROM[11829] <= 32'b00000000010000010000000100010011;
ROM[11830] <= 32'b00000000001100010010000000100011;
ROM[11831] <= 32'b00000000010000010000000100010011;
ROM[11832] <= 32'b00000000010000010010000000100011;
ROM[11833] <= 32'b00000000010000010000000100010011;
ROM[11834] <= 32'b00000000010100010010000000100011;
ROM[11835] <= 32'b00000000010000010000000100010011;
ROM[11836] <= 32'b00000000011000010010000000100011;
ROM[11837] <= 32'b00000000010000010000000100010011;
ROM[11838] <= 32'b00000001010000000000001110010011;
ROM[11839] <= 32'b00000000100000111000001110010011;
ROM[11840] <= 32'b01000000011100010000001110110011;
ROM[11841] <= 32'b00000000011100000000001000110011;
ROM[11842] <= 32'b00000000001000000000000110110011;
ROM[11843] <= 32'b00101010000000011110000011101111;
ROM[11844] <= 32'b00000110011100000000001110010011;
ROM[11845] <= 32'b00000000011100010010000000100011;
ROM[11846] <= 32'b00000000010000010000000100010011;
ROM[11847] <= 32'b00000000000000001100001110110111;
ROM[11848] <= 32'b10010110100000111000001110010011;
ROM[11849] <= 32'b00000000111000111000001110110011;
ROM[11850] <= 32'b00000000011100010010000000100011;
ROM[11851] <= 32'b00000000010000010000000100010011;
ROM[11852] <= 32'b00000000001100010010000000100011;
ROM[11853] <= 32'b00000000010000010000000100010011;
ROM[11854] <= 32'b00000000010000010010000000100011;
ROM[11855] <= 32'b00000000010000010000000100010011;
ROM[11856] <= 32'b00000000010100010010000000100011;
ROM[11857] <= 32'b00000000010000010000000100010011;
ROM[11858] <= 32'b00000000011000010010000000100011;
ROM[11859] <= 32'b00000000010000010000000100010011;
ROM[11860] <= 32'b00000001010000000000001110010011;
ROM[11861] <= 32'b00000000100000111000001110010011;
ROM[11862] <= 32'b01000000011100010000001110110011;
ROM[11863] <= 32'b00000000011100000000001000110011;
ROM[11864] <= 32'b00000000001000000000000110110011;
ROM[11865] <= 32'b00100100100000011110000011101111;
ROM[11866] <= 32'b00000010000000000000001110010011;
ROM[11867] <= 32'b00000000011100010010000000100011;
ROM[11868] <= 32'b00000000010000010000000100010011;
ROM[11869] <= 32'b00000000000000001100001110110111;
ROM[11870] <= 32'b10011100000000111000001110010011;
ROM[11871] <= 32'b00000000111000111000001110110011;
ROM[11872] <= 32'b00000000011100010010000000100011;
ROM[11873] <= 32'b00000000010000010000000100010011;
ROM[11874] <= 32'b00000000001100010010000000100011;
ROM[11875] <= 32'b00000000010000010000000100010011;
ROM[11876] <= 32'b00000000010000010010000000100011;
ROM[11877] <= 32'b00000000010000010000000100010011;
ROM[11878] <= 32'b00000000010100010010000000100011;
ROM[11879] <= 32'b00000000010000010000000100010011;
ROM[11880] <= 32'b00000000011000010010000000100011;
ROM[11881] <= 32'b00000000010000010000000100010011;
ROM[11882] <= 32'b00000001010000000000001110010011;
ROM[11883] <= 32'b00000000100000111000001110010011;
ROM[11884] <= 32'b01000000011100010000001110110011;
ROM[11885] <= 32'b00000000011100000000001000110011;
ROM[11886] <= 32'b00000000001000000000000110110011;
ROM[11887] <= 32'b00011111000000011110000011101111;
ROM[11888] <= 32'b00000110011100000000001110010011;
ROM[11889] <= 32'b00000000011100010010000000100011;
ROM[11890] <= 32'b00000000010000010000000100010011;
ROM[11891] <= 32'b00000000000000001100001110110111;
ROM[11892] <= 32'b10100001100000111000001110010011;
ROM[11893] <= 32'b00000000111000111000001110110011;
ROM[11894] <= 32'b00000000011100010010000000100011;
ROM[11895] <= 32'b00000000010000010000000100010011;
ROM[11896] <= 32'b00000000001100010010000000100011;
ROM[11897] <= 32'b00000000010000010000000100010011;
ROM[11898] <= 32'b00000000010000010010000000100011;
ROM[11899] <= 32'b00000000010000010000000100010011;
ROM[11900] <= 32'b00000000010100010010000000100011;
ROM[11901] <= 32'b00000000010000010000000100010011;
ROM[11902] <= 32'b00000000011000010010000000100011;
ROM[11903] <= 32'b00000000010000010000000100010011;
ROM[11904] <= 32'b00000001010000000000001110010011;
ROM[11905] <= 32'b00000000100000111000001110010011;
ROM[11906] <= 32'b01000000011100010000001110110011;
ROM[11907] <= 32'b00000000011100000000001000110011;
ROM[11908] <= 32'b00000000001000000000000110110011;
ROM[11909] <= 32'b00011001100000011110000011101111;
ROM[11910] <= 32'b00000111010100000000001110010011;
ROM[11911] <= 32'b00000000011100010010000000100011;
ROM[11912] <= 32'b00000000010000010000000100010011;
ROM[11913] <= 32'b00000000000000001100001110110111;
ROM[11914] <= 32'b10100111000000111000001110010011;
ROM[11915] <= 32'b00000000111000111000001110110011;
ROM[11916] <= 32'b00000000011100010010000000100011;
ROM[11917] <= 32'b00000000010000010000000100010011;
ROM[11918] <= 32'b00000000001100010010000000100011;
ROM[11919] <= 32'b00000000010000010000000100010011;
ROM[11920] <= 32'b00000000010000010010000000100011;
ROM[11921] <= 32'b00000000010000010000000100010011;
ROM[11922] <= 32'b00000000010100010010000000100011;
ROM[11923] <= 32'b00000000010000010000000100010011;
ROM[11924] <= 32'b00000000011000010010000000100011;
ROM[11925] <= 32'b00000000010000010000000100010011;
ROM[11926] <= 32'b00000001010000000000001110010011;
ROM[11927] <= 32'b00000000100000111000001110010011;
ROM[11928] <= 32'b01000000011100010000001110110011;
ROM[11929] <= 32'b00000000011100000000001000110011;
ROM[11930] <= 32'b00000000001000000000000110110011;
ROM[11931] <= 32'b00010100000000011110000011101111;
ROM[11932] <= 32'b00000110010100000000001110010011;
ROM[11933] <= 32'b00000000011100010010000000100011;
ROM[11934] <= 32'b00000000010000010000000100010011;
ROM[11935] <= 32'b00000000000000001100001110110111;
ROM[11936] <= 32'b10101100100000111000001110010011;
ROM[11937] <= 32'b00000000111000111000001110110011;
ROM[11938] <= 32'b00000000011100010010000000100011;
ROM[11939] <= 32'b00000000010000010000000100010011;
ROM[11940] <= 32'b00000000001100010010000000100011;
ROM[11941] <= 32'b00000000010000010000000100010011;
ROM[11942] <= 32'b00000000010000010010000000100011;
ROM[11943] <= 32'b00000000010000010000000100010011;
ROM[11944] <= 32'b00000000010100010010000000100011;
ROM[11945] <= 32'b00000000010000010000000100010011;
ROM[11946] <= 32'b00000000011000010010000000100011;
ROM[11947] <= 32'b00000000010000010000000100010011;
ROM[11948] <= 32'b00000001010000000000001110010011;
ROM[11949] <= 32'b00000000100000111000001110010011;
ROM[11950] <= 32'b01000000011100010000001110110011;
ROM[11951] <= 32'b00000000011100000000001000110011;
ROM[11952] <= 32'b00000000001000000000000110110011;
ROM[11953] <= 32'b00001110100000011110000011101111;
ROM[11954] <= 32'b00000111001100000000001110010011;
ROM[11955] <= 32'b00000000011100010010000000100011;
ROM[11956] <= 32'b00000000010000010000000100010011;
ROM[11957] <= 32'b00000000000000001100001110110111;
ROM[11958] <= 32'b10110010000000111000001110010011;
ROM[11959] <= 32'b00000000111000111000001110110011;
ROM[11960] <= 32'b00000000011100010010000000100011;
ROM[11961] <= 32'b00000000010000010000000100010011;
ROM[11962] <= 32'b00000000001100010010000000100011;
ROM[11963] <= 32'b00000000010000010000000100010011;
ROM[11964] <= 32'b00000000010000010010000000100011;
ROM[11965] <= 32'b00000000010000010000000100010011;
ROM[11966] <= 32'b00000000010100010010000000100011;
ROM[11967] <= 32'b00000000010000010000000100010011;
ROM[11968] <= 32'b00000000011000010010000000100011;
ROM[11969] <= 32'b00000000010000010000000100010011;
ROM[11970] <= 32'b00000001010000000000001110010011;
ROM[11971] <= 32'b00000000100000111000001110010011;
ROM[11972] <= 32'b01000000011100010000001110110011;
ROM[11973] <= 32'b00000000011100000000001000110011;
ROM[11974] <= 32'b00000000001000000000000110110011;
ROM[11975] <= 32'b00001001000000011110000011101111;
ROM[11976] <= 32'b00000111001100000000001110010011;
ROM[11977] <= 32'b00000000011100010010000000100011;
ROM[11978] <= 32'b00000000010000010000000100010011;
ROM[11979] <= 32'b00000000000000001100001110110111;
ROM[11980] <= 32'b10110111100000111000001110010011;
ROM[11981] <= 32'b00000000111000111000001110110011;
ROM[11982] <= 32'b00000000011100010010000000100011;
ROM[11983] <= 32'b00000000010000010000000100010011;
ROM[11984] <= 32'b00000000001100010010000000100011;
ROM[11985] <= 32'b00000000010000010000000100010011;
ROM[11986] <= 32'b00000000010000010010000000100011;
ROM[11987] <= 32'b00000000010000010000000100010011;
ROM[11988] <= 32'b00000000010100010010000000100011;
ROM[11989] <= 32'b00000000010000010000000100010011;
ROM[11990] <= 32'b00000000011000010010000000100011;
ROM[11991] <= 32'b00000000010000010000000100010011;
ROM[11992] <= 32'b00000001010000000000001110010011;
ROM[11993] <= 32'b00000000100000111000001110010011;
ROM[11994] <= 32'b01000000011100010000001110110011;
ROM[11995] <= 32'b00000000011100000000001000110011;
ROM[11996] <= 32'b00000000001000000000000110110011;
ROM[11997] <= 32'b00000011100000011110000011101111;
ROM[11998] <= 32'b00000010110000000000001110010011;
ROM[11999] <= 32'b00000000011100010010000000100011;
ROM[12000] <= 32'b00000000010000010000000100010011;
ROM[12001] <= 32'b00000000000000001100001110110111;
ROM[12002] <= 32'b10111101000000111000001110010011;
ROM[12003] <= 32'b00000000111000111000001110110011;
ROM[12004] <= 32'b00000000011100010010000000100011;
ROM[12005] <= 32'b00000000010000010000000100010011;
ROM[12006] <= 32'b00000000001100010010000000100011;
ROM[12007] <= 32'b00000000010000010000000100010011;
ROM[12008] <= 32'b00000000010000010010000000100011;
ROM[12009] <= 32'b00000000010000010000000100010011;
ROM[12010] <= 32'b00000000010100010010000000100011;
ROM[12011] <= 32'b00000000010000010000000100010011;
ROM[12012] <= 32'b00000000011000010010000000100011;
ROM[12013] <= 32'b00000000010000010000000100010011;
ROM[12014] <= 32'b00000001010000000000001110010011;
ROM[12015] <= 32'b00000000100000111000001110010011;
ROM[12016] <= 32'b01000000011100010000001110110011;
ROM[12017] <= 32'b00000000011100000000001000110011;
ROM[12018] <= 32'b00000000001000000000000110110011;
ROM[12019] <= 32'b01111110000100011101000011101111;
ROM[12020] <= 32'b00000010000000000000001110010011;
ROM[12021] <= 32'b00000000011100010010000000100011;
ROM[12022] <= 32'b00000000010000010000000100010011;
ROM[12023] <= 32'b00000000000000001100001110110111;
ROM[12024] <= 32'b11000010100000111000001110010011;
ROM[12025] <= 32'b00000000111000111000001110110011;
ROM[12026] <= 32'b00000000011100010010000000100011;
ROM[12027] <= 32'b00000000010000010000000100010011;
ROM[12028] <= 32'b00000000001100010010000000100011;
ROM[12029] <= 32'b00000000010000010000000100010011;
ROM[12030] <= 32'b00000000010000010010000000100011;
ROM[12031] <= 32'b00000000010000010000000100010011;
ROM[12032] <= 32'b00000000010100010010000000100011;
ROM[12033] <= 32'b00000000010000010000000100010011;
ROM[12034] <= 32'b00000000011000010010000000100011;
ROM[12035] <= 32'b00000000010000010000000100010011;
ROM[12036] <= 32'b00000001010000000000001110010011;
ROM[12037] <= 32'b00000000100000111000001110010011;
ROM[12038] <= 32'b01000000011100010000001110110011;
ROM[12039] <= 32'b00000000011100000000001000110011;
ROM[12040] <= 32'b00000000001000000000000110110011;
ROM[12041] <= 32'b01111000100100011101000011101111;
ROM[12042] <= 32'b00000110011100000000001110010011;
ROM[12043] <= 32'b00000000011100010010000000100011;
ROM[12044] <= 32'b00000000010000010000000100010011;
ROM[12045] <= 32'b00000000000000001100001110110111;
ROM[12046] <= 32'b11001000000000111000001110010011;
ROM[12047] <= 32'b00000000111000111000001110110011;
ROM[12048] <= 32'b00000000011100010010000000100011;
ROM[12049] <= 32'b00000000010000010000000100010011;
ROM[12050] <= 32'b00000000001100010010000000100011;
ROM[12051] <= 32'b00000000010000010000000100010011;
ROM[12052] <= 32'b00000000010000010010000000100011;
ROM[12053] <= 32'b00000000010000010000000100010011;
ROM[12054] <= 32'b00000000010100010010000000100011;
ROM[12055] <= 32'b00000000010000010000000100010011;
ROM[12056] <= 32'b00000000011000010010000000100011;
ROM[12057] <= 32'b00000000010000010000000100010011;
ROM[12058] <= 32'b00000001010000000000001110010011;
ROM[12059] <= 32'b00000000100000111000001110010011;
ROM[12060] <= 32'b01000000011100010000001110110011;
ROM[12061] <= 32'b00000000011100000000001000110011;
ROM[12062] <= 32'b00000000001000000000000110110011;
ROM[12063] <= 32'b01110011000100011101000011101111;
ROM[12064] <= 32'b00000110000100000000001110010011;
ROM[12065] <= 32'b00000000011100010010000000100011;
ROM[12066] <= 32'b00000000010000010000000100010011;
ROM[12067] <= 32'b00000000000000001100001110110111;
ROM[12068] <= 32'b11001101100000111000001110010011;
ROM[12069] <= 32'b00000000111000111000001110110011;
ROM[12070] <= 32'b00000000011100010010000000100011;
ROM[12071] <= 32'b00000000010000010000000100010011;
ROM[12072] <= 32'b00000000001100010010000000100011;
ROM[12073] <= 32'b00000000010000010000000100010011;
ROM[12074] <= 32'b00000000010000010010000000100011;
ROM[12075] <= 32'b00000000010000010000000100010011;
ROM[12076] <= 32'b00000000010100010010000000100011;
ROM[12077] <= 32'b00000000010000010000000100010011;
ROM[12078] <= 32'b00000000011000010010000000100011;
ROM[12079] <= 32'b00000000010000010000000100010011;
ROM[12080] <= 32'b00000001010000000000001110010011;
ROM[12081] <= 32'b00000000100000111000001110010011;
ROM[12082] <= 32'b01000000011100010000001110110011;
ROM[12083] <= 32'b00000000011100000000001000110011;
ROM[12084] <= 32'b00000000001000000000000110110011;
ROM[12085] <= 32'b01101101100100011101000011101111;
ROM[12086] <= 32'b00000110110100000000001110010011;
ROM[12087] <= 32'b00000000011100010010000000100011;
ROM[12088] <= 32'b00000000010000010000000100010011;
ROM[12089] <= 32'b00000000000000001100001110110111;
ROM[12090] <= 32'b11010011000000111000001110010011;
ROM[12091] <= 32'b00000000111000111000001110110011;
ROM[12092] <= 32'b00000000011100010010000000100011;
ROM[12093] <= 32'b00000000010000010000000100010011;
ROM[12094] <= 32'b00000000001100010010000000100011;
ROM[12095] <= 32'b00000000010000010000000100010011;
ROM[12096] <= 32'b00000000010000010010000000100011;
ROM[12097] <= 32'b00000000010000010000000100010011;
ROM[12098] <= 32'b00000000010100010010000000100011;
ROM[12099] <= 32'b00000000010000010000000100010011;
ROM[12100] <= 32'b00000000011000010010000000100011;
ROM[12101] <= 32'b00000000010000010000000100010011;
ROM[12102] <= 32'b00000001010000000000001110010011;
ROM[12103] <= 32'b00000000100000111000001110010011;
ROM[12104] <= 32'b01000000011100010000001110110011;
ROM[12105] <= 32'b00000000011100000000001000110011;
ROM[12106] <= 32'b00000000001000000000000110110011;
ROM[12107] <= 32'b01101000000100011101000011101111;
ROM[12108] <= 32'b00000110010100000000001110010011;
ROM[12109] <= 32'b00000000011100010010000000100011;
ROM[12110] <= 32'b00000000010000010000000100010011;
ROM[12111] <= 32'b00000000000000001100001110110111;
ROM[12112] <= 32'b11011000100000111000001110010011;
ROM[12113] <= 32'b00000000111000111000001110110011;
ROM[12114] <= 32'b00000000011100010010000000100011;
ROM[12115] <= 32'b00000000010000010000000100010011;
ROM[12116] <= 32'b00000000001100010010000000100011;
ROM[12117] <= 32'b00000000010000010000000100010011;
ROM[12118] <= 32'b00000000010000010010000000100011;
ROM[12119] <= 32'b00000000010000010000000100010011;
ROM[12120] <= 32'b00000000010100010010000000100011;
ROM[12121] <= 32'b00000000010000010000000100010011;
ROM[12122] <= 32'b00000000011000010010000000100011;
ROM[12123] <= 32'b00000000010000010000000100010011;
ROM[12124] <= 32'b00000001010000000000001110010011;
ROM[12125] <= 32'b00000000100000111000001110010011;
ROM[12126] <= 32'b01000000011100010000001110110011;
ROM[12127] <= 32'b00000000011100000000001000110011;
ROM[12128] <= 32'b00000000001000000000000110110011;
ROM[12129] <= 32'b01100010100100011101000011101111;
ROM[12130] <= 32'b00000010000000000000001110010011;
ROM[12131] <= 32'b00000000011100010010000000100011;
ROM[12132] <= 32'b00000000010000010000000100010011;
ROM[12133] <= 32'b00000000000000001100001110110111;
ROM[12134] <= 32'b11011110000000111000001110010011;
ROM[12135] <= 32'b00000000111000111000001110110011;
ROM[12136] <= 32'b00000000011100010010000000100011;
ROM[12137] <= 32'b00000000010000010000000100010011;
ROM[12138] <= 32'b00000000001100010010000000100011;
ROM[12139] <= 32'b00000000010000010000000100010011;
ROM[12140] <= 32'b00000000010000010010000000100011;
ROM[12141] <= 32'b00000000010000010000000100010011;
ROM[12142] <= 32'b00000000010100010010000000100011;
ROM[12143] <= 32'b00000000010000010000000100010011;
ROM[12144] <= 32'b00000000011000010010000000100011;
ROM[12145] <= 32'b00000000010000010000000100010011;
ROM[12146] <= 32'b00000001010000000000001110010011;
ROM[12147] <= 32'b00000000100000111000001110010011;
ROM[12148] <= 32'b01000000011100010000001110110011;
ROM[12149] <= 32'b00000000011100000000001000110011;
ROM[12150] <= 32'b00000000001000000000000110110011;
ROM[12151] <= 32'b01011101000100011101000011101111;
ROM[12152] <= 32'b00000110111100000000001110010011;
ROM[12153] <= 32'b00000000011100010010000000100011;
ROM[12154] <= 32'b00000000010000010000000100010011;
ROM[12155] <= 32'b00000000000000001100001110110111;
ROM[12156] <= 32'b11100011100000111000001110010011;
ROM[12157] <= 32'b00000000111000111000001110110011;
ROM[12158] <= 32'b00000000011100010010000000100011;
ROM[12159] <= 32'b00000000010000010000000100010011;
ROM[12160] <= 32'b00000000001100010010000000100011;
ROM[12161] <= 32'b00000000010000010000000100010011;
ROM[12162] <= 32'b00000000010000010010000000100011;
ROM[12163] <= 32'b00000000010000010000000100010011;
ROM[12164] <= 32'b00000000010100010010000000100011;
ROM[12165] <= 32'b00000000010000010000000100010011;
ROM[12166] <= 32'b00000000011000010010000000100011;
ROM[12167] <= 32'b00000000010000010000000100010011;
ROM[12168] <= 32'b00000001010000000000001110010011;
ROM[12169] <= 32'b00000000100000111000001110010011;
ROM[12170] <= 32'b01000000011100010000001110110011;
ROM[12171] <= 32'b00000000011100000000001000110011;
ROM[12172] <= 32'b00000000001000000000000110110011;
ROM[12173] <= 32'b01010111100100011101000011101111;
ROM[12174] <= 32'b00000111011000000000001110010011;
ROM[12175] <= 32'b00000000011100010010000000100011;
ROM[12176] <= 32'b00000000010000010000000100010011;
ROM[12177] <= 32'b00000000000000001100001110110111;
ROM[12178] <= 32'b11101001000000111000001110010011;
ROM[12179] <= 32'b00000000111000111000001110110011;
ROM[12180] <= 32'b00000000011100010010000000100011;
ROM[12181] <= 32'b00000000010000010000000100010011;
ROM[12182] <= 32'b00000000001100010010000000100011;
ROM[12183] <= 32'b00000000010000010000000100010011;
ROM[12184] <= 32'b00000000010000010010000000100011;
ROM[12185] <= 32'b00000000010000010000000100010011;
ROM[12186] <= 32'b00000000010100010010000000100011;
ROM[12187] <= 32'b00000000010000010000000100010011;
ROM[12188] <= 32'b00000000011000010010000000100011;
ROM[12189] <= 32'b00000000010000010000000100010011;
ROM[12190] <= 32'b00000001010000000000001110010011;
ROM[12191] <= 32'b00000000100000111000001110010011;
ROM[12192] <= 32'b01000000011100010000001110110011;
ROM[12193] <= 32'b00000000011100000000001000110011;
ROM[12194] <= 32'b00000000001000000000000110110011;
ROM[12195] <= 32'b01010010000100011101000011101111;
ROM[12196] <= 32'b00000110010100000000001110010011;
ROM[12197] <= 32'b00000000011100010010000000100011;
ROM[12198] <= 32'b00000000010000010000000100010011;
ROM[12199] <= 32'b00000000000000001100001110110111;
ROM[12200] <= 32'b11101110100000111000001110010011;
ROM[12201] <= 32'b00000000111000111000001110110011;
ROM[12202] <= 32'b00000000011100010010000000100011;
ROM[12203] <= 32'b00000000010000010000000100010011;
ROM[12204] <= 32'b00000000001100010010000000100011;
ROM[12205] <= 32'b00000000010000010000000100010011;
ROM[12206] <= 32'b00000000010000010010000000100011;
ROM[12207] <= 32'b00000000010000010000000100010011;
ROM[12208] <= 32'b00000000010100010010000000100011;
ROM[12209] <= 32'b00000000010000010000000100010011;
ROM[12210] <= 32'b00000000011000010010000000100011;
ROM[12211] <= 32'b00000000010000010000000100010011;
ROM[12212] <= 32'b00000001010000000000001110010011;
ROM[12213] <= 32'b00000000100000111000001110010011;
ROM[12214] <= 32'b01000000011100010000001110110011;
ROM[12215] <= 32'b00000000011100000000001000110011;
ROM[12216] <= 32'b00000000001000000000000110110011;
ROM[12217] <= 32'b01001100100100011101000011101111;
ROM[12218] <= 32'b00000111001000000000001110010011;
ROM[12219] <= 32'b00000000011100010010000000100011;
ROM[12220] <= 32'b00000000010000010000000100010011;
ROM[12221] <= 32'b00000000000000001100001110110111;
ROM[12222] <= 32'b11110100000000111000001110010011;
ROM[12223] <= 32'b00000000111000111000001110110011;
ROM[12224] <= 32'b00000000011100010010000000100011;
ROM[12225] <= 32'b00000000010000010000000100010011;
ROM[12226] <= 32'b00000000001100010010000000100011;
ROM[12227] <= 32'b00000000010000010000000100010011;
ROM[12228] <= 32'b00000000010000010010000000100011;
ROM[12229] <= 32'b00000000010000010000000100010011;
ROM[12230] <= 32'b00000000010100010010000000100011;
ROM[12231] <= 32'b00000000010000010000000100010011;
ROM[12232] <= 32'b00000000011000010010000000100011;
ROM[12233] <= 32'b00000000010000010000000100010011;
ROM[12234] <= 32'b00000001010000000000001110010011;
ROM[12235] <= 32'b00000000100000111000001110010011;
ROM[12236] <= 32'b01000000011100010000001110110011;
ROM[12237] <= 32'b00000000011100000000001000110011;
ROM[12238] <= 32'b00000000001000000000000110110011;
ROM[12239] <= 32'b01000111000100011101000011101111;
ROM[12240] <= 32'b00000010000100000000001110010011;
ROM[12241] <= 32'b00000000011100010010000000100011;
ROM[12242] <= 32'b00000000010000010000000100010011;
ROM[12243] <= 32'b00000000000000001100001110110111;
ROM[12244] <= 32'b11111001100000111000001110010011;
ROM[12245] <= 32'b00000000111000111000001110110011;
ROM[12246] <= 32'b00000000011100010010000000100011;
ROM[12247] <= 32'b00000000010000010000000100010011;
ROM[12248] <= 32'b00000000001100010010000000100011;
ROM[12249] <= 32'b00000000010000010000000100010011;
ROM[12250] <= 32'b00000000010000010010000000100011;
ROM[12251] <= 32'b00000000010000010000000100010011;
ROM[12252] <= 32'b00000000010100010010000000100011;
ROM[12253] <= 32'b00000000010000010000000100010011;
ROM[12254] <= 32'b00000000011000010010000000100011;
ROM[12255] <= 32'b00000000010000010000000100010011;
ROM[12256] <= 32'b00000001010000000000001110010011;
ROM[12257] <= 32'b00000000100000111000001110010011;
ROM[12258] <= 32'b01000000011100010000001110110011;
ROM[12259] <= 32'b00000000011100000000001000110011;
ROM[12260] <= 32'b00000000001000000000000110110011;
ROM[12261] <= 32'b01000001100100011101000011101111;
ROM[12262] <= 32'b00000000000000001100001110110111;
ROM[12263] <= 32'b11111110010000111000001110010011;
ROM[12264] <= 32'b00000000111000111000001110110011;
ROM[12265] <= 32'b00000000011100010010000000100011;
ROM[12266] <= 32'b00000000010000010000000100010011;
ROM[12267] <= 32'b00000000001100010010000000100011;
ROM[12268] <= 32'b00000000010000010000000100010011;
ROM[12269] <= 32'b00000000010000010010000000100011;
ROM[12270] <= 32'b00000000010000010000000100010011;
ROM[12271] <= 32'b00000000010100010010000000100011;
ROM[12272] <= 32'b00000000010000010000000100010011;
ROM[12273] <= 32'b00000000011000010010000000100011;
ROM[12274] <= 32'b00000000010000010000000100010011;
ROM[12275] <= 32'b00000001010000000000001110010011;
ROM[12276] <= 32'b00000000010000111000001110010011;
ROM[12277] <= 32'b01000000011100010000001110110011;
ROM[12278] <= 32'b00000000011100000000001000110011;
ROM[12279] <= 32'b00000000001000000000000110110011;
ROM[12280] <= 32'b01111000100100001010000011101111;
ROM[12281] <= 32'b11111111110000010000000100010011;
ROM[12282] <= 32'b00000000000000010010001110000011;
ROM[12283] <= 32'b00000000011101100010000000100011;
ROM[12284] <= 32'b00000000000000001100001110110111;
ROM[12285] <= 32'b00000011110000111000001110010011;
ROM[12286] <= 32'b00000000111000111000001110110011;
ROM[12287] <= 32'b00000000011100010010000000100011;
ROM[12288] <= 32'b00000000010000010000000100010011;
ROM[12289] <= 32'b00000000001100010010000000100011;
ROM[12290] <= 32'b00000000010000010000000100010011;
ROM[12291] <= 32'b00000000010000010010000000100011;
ROM[12292] <= 32'b00000000010000010000000100010011;
ROM[12293] <= 32'b00000000010100010010000000100011;
ROM[12294] <= 32'b00000000010000010000000100010011;
ROM[12295] <= 32'b00000000011000010010000000100011;
ROM[12296] <= 32'b00000000010000010000000100010011;
ROM[12297] <= 32'b00000001010000000000001110010011;
ROM[12298] <= 32'b00000000000000111000001110010011;
ROM[12299] <= 32'b01000000011100010000001110110011;
ROM[12300] <= 32'b00000000011100000000001000110011;
ROM[12301] <= 32'b00000000001000000000000110110011;
ROM[12302] <= 32'b00110011000000001011000011101111;
ROM[12303] <= 32'b11111111110000010000000100010011;
ROM[12304] <= 32'b00000000000000010010001110000011;
ROM[12305] <= 32'b00000000011101100010000000100011;
ROM[12306] <= 32'b00000000101100000000001110010011;
ROM[12307] <= 32'b00000000011100010010000000100011;
ROM[12308] <= 32'b00000000010000010000000100010011;
ROM[12309] <= 32'b00000000000000001100001110110111;
ROM[12310] <= 32'b00001010000000111000001110010011;
ROM[12311] <= 32'b00000000111000111000001110110011;
ROM[12312] <= 32'b00000000011100010010000000100011;
ROM[12313] <= 32'b00000000010000010000000100010011;
ROM[12314] <= 32'b00000000001100010010000000100011;
ROM[12315] <= 32'b00000000010000010000000100010011;
ROM[12316] <= 32'b00000000010000010010000000100011;
ROM[12317] <= 32'b00000000010000010000000100010011;
ROM[12318] <= 32'b00000000010100010010000000100011;
ROM[12319] <= 32'b00000000010000010000000100010011;
ROM[12320] <= 32'b00000000011000010010000000100011;
ROM[12321] <= 32'b00000000010000010000000100010011;
ROM[12322] <= 32'b00000001010000000000001110010011;
ROM[12323] <= 32'b00000000010000111000001110010011;
ROM[12324] <= 32'b01000000011100010000001110110011;
ROM[12325] <= 32'b00000000011100000000001000110011;
ROM[12326] <= 32'b00000000001000000000000110110011;
ROM[12327] <= 32'b01101010000000011101000011101111;
ROM[12328] <= 32'b00000101010000000000001110010011;
ROM[12329] <= 32'b00000000011100010010000000100011;
ROM[12330] <= 32'b00000000010000010000000100010011;
ROM[12331] <= 32'b00000000000000001100001110110111;
ROM[12332] <= 32'b00001111100000111000001110010011;
ROM[12333] <= 32'b00000000111000111000001110110011;
ROM[12334] <= 32'b00000000011100010010000000100011;
ROM[12335] <= 32'b00000000010000010000000100010011;
ROM[12336] <= 32'b00000000001100010010000000100011;
ROM[12337] <= 32'b00000000010000010000000100010011;
ROM[12338] <= 32'b00000000010000010010000000100011;
ROM[12339] <= 32'b00000000010000010000000100010011;
ROM[12340] <= 32'b00000000010100010010000000100011;
ROM[12341] <= 32'b00000000010000010000000100010011;
ROM[12342] <= 32'b00000000011000010010000000100011;
ROM[12343] <= 32'b00000000010000010000000100010011;
ROM[12344] <= 32'b00000001010000000000001110010011;
ROM[12345] <= 32'b00000000100000111000001110010011;
ROM[12346] <= 32'b01000000011100010000001110110011;
ROM[12347] <= 32'b00000000011100000000001000110011;
ROM[12348] <= 32'b00000000001000000000000110110011;
ROM[12349] <= 32'b00101011100100011101000011101111;
ROM[12350] <= 32'b00000110100000000000001110010011;
ROM[12351] <= 32'b00000000011100010010000000100011;
ROM[12352] <= 32'b00000000010000010000000100010011;
ROM[12353] <= 32'b00000000000000001100001110110111;
ROM[12354] <= 32'b00010101000000111000001110010011;
ROM[12355] <= 32'b00000000111000111000001110110011;
ROM[12356] <= 32'b00000000011100010010000000100011;
ROM[12357] <= 32'b00000000010000010000000100010011;
ROM[12358] <= 32'b00000000001100010010000000100011;
ROM[12359] <= 32'b00000000010000010000000100010011;
ROM[12360] <= 32'b00000000010000010010000000100011;
ROM[12361] <= 32'b00000000010000010000000100010011;
ROM[12362] <= 32'b00000000010100010010000000100011;
ROM[12363] <= 32'b00000000010000010000000100010011;
ROM[12364] <= 32'b00000000011000010010000000100011;
ROM[12365] <= 32'b00000000010000010000000100010011;
ROM[12366] <= 32'b00000001010000000000001110010011;
ROM[12367] <= 32'b00000000100000111000001110010011;
ROM[12368] <= 32'b01000000011100010000001110110011;
ROM[12369] <= 32'b00000000011100000000001000110011;
ROM[12370] <= 32'b00000000001000000000000110110011;
ROM[12371] <= 32'b00100110000100011101000011101111;
ROM[12372] <= 32'b00000110010100000000001110010011;
ROM[12373] <= 32'b00000000011100010010000000100011;
ROM[12374] <= 32'b00000000010000010000000100010011;
ROM[12375] <= 32'b00000000000000001100001110110111;
ROM[12376] <= 32'b00011010100000111000001110010011;
ROM[12377] <= 32'b00000000111000111000001110110011;
ROM[12378] <= 32'b00000000011100010010000000100011;
ROM[12379] <= 32'b00000000010000010000000100010011;
ROM[12380] <= 32'b00000000001100010010000000100011;
ROM[12381] <= 32'b00000000010000010000000100010011;
ROM[12382] <= 32'b00000000010000010010000000100011;
ROM[12383] <= 32'b00000000010000010000000100010011;
ROM[12384] <= 32'b00000000010100010010000000100011;
ROM[12385] <= 32'b00000000010000010000000100010011;
ROM[12386] <= 32'b00000000011000010010000000100011;
ROM[12387] <= 32'b00000000010000010000000100010011;
ROM[12388] <= 32'b00000001010000000000001110010011;
ROM[12389] <= 32'b00000000100000111000001110010011;
ROM[12390] <= 32'b01000000011100010000001110110011;
ROM[12391] <= 32'b00000000011100000000001000110011;
ROM[12392] <= 32'b00000000001000000000000110110011;
ROM[12393] <= 32'b00100000100100011101000011101111;
ROM[12394] <= 32'b00000010000000000000001110010011;
ROM[12395] <= 32'b00000000011100010010000000100011;
ROM[12396] <= 32'b00000000010000010000000100010011;
ROM[12397] <= 32'b00000000000000001100001110110111;
ROM[12398] <= 32'b00100000000000111000001110010011;
ROM[12399] <= 32'b00000000111000111000001110110011;
ROM[12400] <= 32'b00000000011100010010000000100011;
ROM[12401] <= 32'b00000000010000010000000100010011;
ROM[12402] <= 32'b00000000001100010010000000100011;
ROM[12403] <= 32'b00000000010000010000000100010011;
ROM[12404] <= 32'b00000000010000010010000000100011;
ROM[12405] <= 32'b00000000010000010000000100010011;
ROM[12406] <= 32'b00000000010100010010000000100011;
ROM[12407] <= 32'b00000000010000010000000100010011;
ROM[12408] <= 32'b00000000011000010010000000100011;
ROM[12409] <= 32'b00000000010000010000000100010011;
ROM[12410] <= 32'b00000001010000000000001110010011;
ROM[12411] <= 32'b00000000100000111000001110010011;
ROM[12412] <= 32'b01000000011100010000001110110011;
ROM[12413] <= 32'b00000000011100000000001000110011;
ROM[12414] <= 32'b00000000001000000000000110110011;
ROM[12415] <= 32'b00011011000100011101000011101111;
ROM[12416] <= 32'b00000111011100000000001110010011;
ROM[12417] <= 32'b00000000011100010010000000100011;
ROM[12418] <= 32'b00000000010000010000000100010011;
ROM[12419] <= 32'b00000000000000001100001110110111;
ROM[12420] <= 32'b00100101100000111000001110010011;
ROM[12421] <= 32'b00000000111000111000001110110011;
ROM[12422] <= 32'b00000000011100010010000000100011;
ROM[12423] <= 32'b00000000010000010000000100010011;
ROM[12424] <= 32'b00000000001100010010000000100011;
ROM[12425] <= 32'b00000000010000010000000100010011;
ROM[12426] <= 32'b00000000010000010010000000100011;
ROM[12427] <= 32'b00000000010000010000000100010011;
ROM[12428] <= 32'b00000000010100010010000000100011;
ROM[12429] <= 32'b00000000010000010000000100010011;
ROM[12430] <= 32'b00000000011000010010000000100011;
ROM[12431] <= 32'b00000000010000010000000100010011;
ROM[12432] <= 32'b00000001010000000000001110010011;
ROM[12433] <= 32'b00000000100000111000001110010011;
ROM[12434] <= 32'b01000000011100010000001110110011;
ROM[12435] <= 32'b00000000011100000000001000110011;
ROM[12436] <= 32'b00000000001000000000000110110011;
ROM[12437] <= 32'b00010101100100011101000011101111;
ROM[12438] <= 32'b00000110111100000000001110010011;
ROM[12439] <= 32'b00000000011100010010000000100011;
ROM[12440] <= 32'b00000000010000010000000100010011;
ROM[12441] <= 32'b00000000000000001100001110110111;
ROM[12442] <= 32'b00101011000000111000001110010011;
ROM[12443] <= 32'b00000000111000111000001110110011;
ROM[12444] <= 32'b00000000011100010010000000100011;
ROM[12445] <= 32'b00000000010000010000000100010011;
ROM[12446] <= 32'b00000000001100010010000000100011;
ROM[12447] <= 32'b00000000010000010000000100010011;
ROM[12448] <= 32'b00000000010000010010000000100011;
ROM[12449] <= 32'b00000000010000010000000100010011;
ROM[12450] <= 32'b00000000010100010010000000100011;
ROM[12451] <= 32'b00000000010000010000000100010011;
ROM[12452] <= 32'b00000000011000010010000000100011;
ROM[12453] <= 32'b00000000010000010000000100010011;
ROM[12454] <= 32'b00000001010000000000001110010011;
ROM[12455] <= 32'b00000000100000111000001110010011;
ROM[12456] <= 32'b01000000011100010000001110110011;
ROM[12457] <= 32'b00000000011100000000001000110011;
ROM[12458] <= 32'b00000000001000000000000110110011;
ROM[12459] <= 32'b00010000000100011101000011101111;
ROM[12460] <= 32'b00000111001000000000001110010011;
ROM[12461] <= 32'b00000000011100010010000000100011;
ROM[12462] <= 32'b00000000010000010000000100010011;
ROM[12463] <= 32'b00000000000000001100001110110111;
ROM[12464] <= 32'b00110000100000111000001110010011;
ROM[12465] <= 32'b00000000111000111000001110110011;
ROM[12466] <= 32'b00000000011100010010000000100011;
ROM[12467] <= 32'b00000000010000010000000100010011;
ROM[12468] <= 32'b00000000001100010010000000100011;
ROM[12469] <= 32'b00000000010000010000000100010011;
ROM[12470] <= 32'b00000000010000010010000000100011;
ROM[12471] <= 32'b00000000010000010000000100010011;
ROM[12472] <= 32'b00000000010100010010000000100011;
ROM[12473] <= 32'b00000000010000010000000100010011;
ROM[12474] <= 32'b00000000011000010010000000100011;
ROM[12475] <= 32'b00000000010000010000000100010011;
ROM[12476] <= 32'b00000001010000000000001110010011;
ROM[12477] <= 32'b00000000100000111000001110010011;
ROM[12478] <= 32'b01000000011100010000001110110011;
ROM[12479] <= 32'b00000000011100000000001000110011;
ROM[12480] <= 32'b00000000001000000000000110110011;
ROM[12481] <= 32'b00001010100100011101000011101111;
ROM[12482] <= 32'b00000110010000000000001110010011;
ROM[12483] <= 32'b00000000011100010010000000100011;
ROM[12484] <= 32'b00000000010000010000000100010011;
ROM[12485] <= 32'b00000000000000001100001110110111;
ROM[12486] <= 32'b00110110000000111000001110010011;
ROM[12487] <= 32'b00000000111000111000001110110011;
ROM[12488] <= 32'b00000000011100010010000000100011;
ROM[12489] <= 32'b00000000010000010000000100010011;
ROM[12490] <= 32'b00000000001100010010000000100011;
ROM[12491] <= 32'b00000000010000010000000100010011;
ROM[12492] <= 32'b00000000010000010010000000100011;
ROM[12493] <= 32'b00000000010000010000000100010011;
ROM[12494] <= 32'b00000000010100010010000000100011;
ROM[12495] <= 32'b00000000010000010000000100010011;
ROM[12496] <= 32'b00000000011000010010000000100011;
ROM[12497] <= 32'b00000000010000010000000100010011;
ROM[12498] <= 32'b00000001010000000000001110010011;
ROM[12499] <= 32'b00000000100000111000001110010011;
ROM[12500] <= 32'b01000000011100010000001110110011;
ROM[12501] <= 32'b00000000011100000000001000110011;
ROM[12502] <= 32'b00000000001000000000000110110011;
ROM[12503] <= 32'b00000101000100011101000011101111;
ROM[12504] <= 32'b00000010000000000000001110010011;
ROM[12505] <= 32'b00000000011100010010000000100011;
ROM[12506] <= 32'b00000000010000010000000100010011;
ROM[12507] <= 32'b00000000000000001100001110110111;
ROM[12508] <= 32'b00111011100000111000001110010011;
ROM[12509] <= 32'b00000000111000111000001110110011;
ROM[12510] <= 32'b00000000011100010010000000100011;
ROM[12511] <= 32'b00000000010000010000000100010011;
ROM[12512] <= 32'b00000000001100010010000000100011;
ROM[12513] <= 32'b00000000010000010000000100010011;
ROM[12514] <= 32'b00000000010000010010000000100011;
ROM[12515] <= 32'b00000000010000010000000100010011;
ROM[12516] <= 32'b00000000010100010010000000100011;
ROM[12517] <= 32'b00000000010000010000000100010011;
ROM[12518] <= 32'b00000000011000010010000000100011;
ROM[12519] <= 32'b00000000010000010000000100010011;
ROM[12520] <= 32'b00000001010000000000001110010011;
ROM[12521] <= 32'b00000000100000111000001110010011;
ROM[12522] <= 32'b01000000011100010000001110110011;
ROM[12523] <= 32'b00000000011100000000001000110011;
ROM[12524] <= 32'b00000000001000000000000110110011;
ROM[12525] <= 32'b01111111100000011101000011101111;
ROM[12526] <= 32'b00000110100100000000001110010011;
ROM[12527] <= 32'b00000000011100010010000000100011;
ROM[12528] <= 32'b00000000010000010000000100010011;
ROM[12529] <= 32'b00000000000000001100001110110111;
ROM[12530] <= 32'b01000001000000111000001110010011;
ROM[12531] <= 32'b00000000111000111000001110110011;
ROM[12532] <= 32'b00000000011100010010000000100011;
ROM[12533] <= 32'b00000000010000010000000100010011;
ROM[12534] <= 32'b00000000001100010010000000100011;
ROM[12535] <= 32'b00000000010000010000000100010011;
ROM[12536] <= 32'b00000000010000010010000000100011;
ROM[12537] <= 32'b00000000010000010000000100010011;
ROM[12538] <= 32'b00000000010100010010000000100011;
ROM[12539] <= 32'b00000000010000010000000100010011;
ROM[12540] <= 32'b00000000011000010010000000100011;
ROM[12541] <= 32'b00000000010000010000000100010011;
ROM[12542] <= 32'b00000001010000000000001110010011;
ROM[12543] <= 32'b00000000100000111000001110010011;
ROM[12544] <= 32'b01000000011100010000001110110011;
ROM[12545] <= 32'b00000000011100000000001000110011;
ROM[12546] <= 32'b00000000001000000000000110110011;
ROM[12547] <= 32'b01111010000000011101000011101111;
ROM[12548] <= 32'b00000111001100000000001110010011;
ROM[12549] <= 32'b00000000011100010010000000100011;
ROM[12550] <= 32'b00000000010000010000000100010011;
ROM[12551] <= 32'b00000000000000001100001110110111;
ROM[12552] <= 32'b01000110100000111000001110010011;
ROM[12553] <= 32'b00000000111000111000001110110011;
ROM[12554] <= 32'b00000000011100010010000000100011;
ROM[12555] <= 32'b00000000010000010000000100010011;
ROM[12556] <= 32'b00000000001100010010000000100011;
ROM[12557] <= 32'b00000000010000010000000100010011;
ROM[12558] <= 32'b00000000010000010010000000100011;
ROM[12559] <= 32'b00000000010000010000000100010011;
ROM[12560] <= 32'b00000000010100010010000000100011;
ROM[12561] <= 32'b00000000010000010000000100010011;
ROM[12562] <= 32'b00000000011000010010000000100011;
ROM[12563] <= 32'b00000000010000010000000100010011;
ROM[12564] <= 32'b00000001010000000000001110010011;
ROM[12565] <= 32'b00000000100000111000001110010011;
ROM[12566] <= 32'b01000000011100010000001110110011;
ROM[12567] <= 32'b00000000011100000000001000110011;
ROM[12568] <= 32'b00000000001000000000000110110011;
ROM[12569] <= 32'b01110100100000011101000011101111;
ROM[12570] <= 32'b00000000000000001100001110110111;
ROM[12571] <= 32'b01001011010000111000001110010011;
ROM[12572] <= 32'b00000000111000111000001110110011;
ROM[12573] <= 32'b00000000011100010010000000100011;
ROM[12574] <= 32'b00000000010000010000000100010011;
ROM[12575] <= 32'b00000000001100010010000000100011;
ROM[12576] <= 32'b00000000010000010000000100010011;
ROM[12577] <= 32'b00000000010000010010000000100011;
ROM[12578] <= 32'b00000000010000010000000100010011;
ROM[12579] <= 32'b00000000010100010010000000100011;
ROM[12580] <= 32'b00000000010000010000000100010011;
ROM[12581] <= 32'b00000000011000010010000000100011;
ROM[12582] <= 32'b00000000010000010000000100010011;
ROM[12583] <= 32'b00000001010000000000001110010011;
ROM[12584] <= 32'b00000000010000111000001110010011;
ROM[12585] <= 32'b01000000011100010000001110110011;
ROM[12586] <= 32'b00000000011100000000001000110011;
ROM[12587] <= 32'b00000000001000000000000110110011;
ROM[12588] <= 32'b00101011100100001010000011101111;
ROM[12589] <= 32'b11111111110000010000000100010011;
ROM[12590] <= 32'b00000000000000010010001110000011;
ROM[12591] <= 32'b00000000011101100010000000100011;
ROM[12592] <= 32'b00000000000000011010001110000011;
ROM[12593] <= 32'b00000000011100010010000000100011;
ROM[12594] <= 32'b00000000010000010000000100010011;
ROM[12595] <= 32'b00000000100000011010001110000011;
ROM[12596] <= 32'b00000000011100010010000000100011;
ROM[12597] <= 32'b00000000010000010000000100010011;
ROM[12598] <= 32'b00000000010000000000001110010011;
ROM[12599] <= 32'b00000000011100010010000000100011;
ROM[12600] <= 32'b00000000010000010000000100010011;
ROM[12601] <= 32'b00000000000000001100001110110111;
ROM[12602] <= 32'b01010011000000111000001110010011;
ROM[12603] <= 32'b00000000111000111000001110110011;
ROM[12604] <= 32'b00000000011100010010000000100011;
ROM[12605] <= 32'b00000000010000010000000100010011;
ROM[12606] <= 32'b00000000001100010010000000100011;
ROM[12607] <= 32'b00000000010000010000000100010011;
ROM[12608] <= 32'b00000000010000010010000000100011;
ROM[12609] <= 32'b00000000010000010000000100010011;
ROM[12610] <= 32'b00000000010100010010000000100011;
ROM[12611] <= 32'b00000000010000010000000100010011;
ROM[12612] <= 32'b00000000011000010010000000100011;
ROM[12613] <= 32'b00000000010000010000000100010011;
ROM[12614] <= 32'b00000001010000000000001110010011;
ROM[12615] <= 32'b00000000100000111000001110010011;
ROM[12616] <= 32'b01000000011100010000001110110011;
ROM[12617] <= 32'b00000000011100000000001000110011;
ROM[12618] <= 32'b00000000001000000000000110110011;
ROM[12619] <= 32'b00110000000000000101000011101111;
ROM[12620] <= 32'b11111111110000010000000100010011;
ROM[12621] <= 32'b00000000000000010010001110000011;
ROM[12622] <= 32'b11111111110000010000000100010011;
ROM[12623] <= 32'b00000000000000010010010000000011;
ROM[12624] <= 32'b00000000011101000000001110110011;
ROM[12625] <= 32'b00000000011100010010000000100011;
ROM[12626] <= 32'b00000000010000010000000100010011;
ROM[12627] <= 32'b11111111110000010000000100010011;
ROM[12628] <= 32'b00000000000000010010001110000011;
ROM[12629] <= 32'b00000000000000111000001100010011;
ROM[12630] <= 32'b00000000110100110000010000110011;
ROM[12631] <= 32'b00000000000001000010001110000011;
ROM[12632] <= 32'b00000000011100010010000000100011;
ROM[12633] <= 32'b00000000010000010000000100010011;
ROM[12634] <= 32'b00000000000000001100001110110111;
ROM[12635] <= 32'b01011011010000111000001110010011;
ROM[12636] <= 32'b00000000111000111000001110110011;
ROM[12637] <= 32'b00000000011100010010000000100011;
ROM[12638] <= 32'b00000000010000010000000100010011;
ROM[12639] <= 32'b00000000001100010010000000100011;
ROM[12640] <= 32'b00000000010000010000000100010011;
ROM[12641] <= 32'b00000000010000010010000000100011;
ROM[12642] <= 32'b00000000010000010000000100010011;
ROM[12643] <= 32'b00000000010100010010000000100011;
ROM[12644] <= 32'b00000000010000010000000100010011;
ROM[12645] <= 32'b00000000011000010010000000100011;
ROM[12646] <= 32'b00000000010000010000000100010011;
ROM[12647] <= 32'b00000001010000000000001110010011;
ROM[12648] <= 32'b00000000010000111000001110010011;
ROM[12649] <= 32'b01000000011100010000001110110011;
ROM[12650] <= 32'b00000000011100000000001000110011;
ROM[12651] <= 32'b00000000001000000000000110110011;
ROM[12652] <= 32'b00011011100100001010000011101111;
ROM[12653] <= 32'b11111111110000010000000100010011;
ROM[12654] <= 32'b00000000000000010010001110000011;
ROM[12655] <= 32'b00000000011101100010000000100011;
ROM[12656] <= 32'b00000000000000001100001110110111;
ROM[12657] <= 32'b01100000110000111000001110010011;
ROM[12658] <= 32'b00000000111000111000001110110011;
ROM[12659] <= 32'b00000000011100010010000000100011;
ROM[12660] <= 32'b00000000010000010000000100010011;
ROM[12661] <= 32'b00000000001100010010000000100011;
ROM[12662] <= 32'b00000000010000010000000100010011;
ROM[12663] <= 32'b00000000010000010010000000100011;
ROM[12664] <= 32'b00000000010000010000000100010011;
ROM[12665] <= 32'b00000000010100010010000000100011;
ROM[12666] <= 32'b00000000010000010000000100010011;
ROM[12667] <= 32'b00000000011000010010000000100011;
ROM[12668] <= 32'b00000000010000010000000100010011;
ROM[12669] <= 32'b00000001010000000000001110010011;
ROM[12670] <= 32'b00000000000000111000001110010011;
ROM[12671] <= 32'b01000000011100010000001110110011;
ROM[12672] <= 32'b00000000011100000000001000110011;
ROM[12673] <= 32'b00000000001000000000000110110011;
ROM[12674] <= 32'b01010110000100001010000011101111;
ROM[12675] <= 32'b11111111110000010000000100010011;
ROM[12676] <= 32'b00000000000000010010001110000011;
ROM[12677] <= 32'b00000000011101100010000000100011;
ROM[12678] <= 32'b00000001010000011010001110000011;
ROM[12679] <= 32'b00000000011100010010000000100011;
ROM[12680] <= 32'b00000000010000010000000100010011;
ROM[12681] <= 32'b00000000000100000000001110010011;
ROM[12682] <= 32'b00000000011100010010000000100011;
ROM[12683] <= 32'b00000000010000010000000100010011;
ROM[12684] <= 32'b11111111110000010000000100010011;
ROM[12685] <= 32'b00000000000000010010001110000011;
ROM[12686] <= 32'b11111111110000010000000100010011;
ROM[12687] <= 32'b00000000000000010010010000000011;
ROM[12688] <= 32'b01000000011101000000001110110011;
ROM[12689] <= 32'b00000000011100010010000000100011;
ROM[12690] <= 32'b00000000010000010000000100010011;
ROM[12691] <= 32'b11111111110000010000000100010011;
ROM[12692] <= 32'b00000000000000010010001110000011;
ROM[12693] <= 32'b00000000011100011010101000100011;
ROM[12694] <= 32'b00000010110000000001000011101111;
ROM[12695] <= 32'b00000010110000000000001110010011;
ROM[12696] <= 32'b00000000011100010010000000100011;
ROM[12697] <= 32'b00000000010000010000000100010011;
ROM[12698] <= 32'b00000000000000001100001110110111;
ROM[12699] <= 32'b01101011010000111000001110010011;
ROM[12700] <= 32'b00000000111000111000001110110011;
ROM[12701] <= 32'b00000000011100010010000000100011;
ROM[12702] <= 32'b00000000010000010000000100010011;
ROM[12703] <= 32'b00000000001100010010000000100011;
ROM[12704] <= 32'b00000000010000010000000100010011;
ROM[12705] <= 32'b00000000010000010010000000100011;
ROM[12706] <= 32'b00000000010000010000000100010011;
ROM[12707] <= 32'b00000000010100010010000000100011;
ROM[12708] <= 32'b00000000010000010000000100010011;
ROM[12709] <= 32'b00000000011000010010000000100011;
ROM[12710] <= 32'b00000000010000010000000100010011;
ROM[12711] <= 32'b00000001010000000000001110010011;
ROM[12712] <= 32'b00000000010000111000001110010011;
ROM[12713] <= 32'b01000000011100010000001110110011;
ROM[12714] <= 32'b00000000011100000000001000110011;
ROM[12715] <= 32'b00000000001000000000000110110011;
ROM[12716] <= 32'b00001000110000011101000011101111;
ROM[12717] <= 32'b00000110110000000000001110010011;
ROM[12718] <= 32'b00000000011100010010000000100011;
ROM[12719] <= 32'b00000000010000010000000100010011;
ROM[12720] <= 32'b00000000000000001100001110110111;
ROM[12721] <= 32'b01110000110000111000001110010011;
ROM[12722] <= 32'b00000000111000111000001110110011;
ROM[12723] <= 32'b00000000011100010010000000100011;
ROM[12724] <= 32'b00000000010000010000000100010011;
ROM[12725] <= 32'b00000000001100010010000000100011;
ROM[12726] <= 32'b00000000010000010000000100010011;
ROM[12727] <= 32'b00000000010000010010000000100011;
ROM[12728] <= 32'b00000000010000010000000100010011;
ROM[12729] <= 32'b00000000010100010010000000100011;
ROM[12730] <= 32'b00000000010000010000000100010011;
ROM[12731] <= 32'b00000000011000010010000000100011;
ROM[12732] <= 32'b00000000010000010000000100010011;
ROM[12733] <= 32'b00000001010000000000001110010011;
ROM[12734] <= 32'b00000000100000111000001110010011;
ROM[12735] <= 32'b01000000011100010000001110110011;
ROM[12736] <= 32'b00000000011100000000001000110011;
ROM[12737] <= 32'b00000000001000000000000110110011;
ROM[12738] <= 32'b01001010010000011101000011101111;
ROM[12739] <= 32'b00000110010100000000001110010011;
ROM[12740] <= 32'b00000000011100010010000000100011;
ROM[12741] <= 32'b00000000010000010000000100010011;
ROM[12742] <= 32'b00000000000000001100001110110111;
ROM[12743] <= 32'b01110110010000111000001110010011;
ROM[12744] <= 32'b00000000111000111000001110110011;
ROM[12745] <= 32'b00000000011100010010000000100011;
ROM[12746] <= 32'b00000000010000010000000100010011;
ROM[12747] <= 32'b00000000001100010010000000100011;
ROM[12748] <= 32'b00000000010000010000000100010011;
ROM[12749] <= 32'b00000000010000010010000000100011;
ROM[12750] <= 32'b00000000010000010000000100010011;
ROM[12751] <= 32'b00000000010100010010000000100011;
ROM[12752] <= 32'b00000000010000010000000100010011;
ROM[12753] <= 32'b00000000011000010010000000100011;
ROM[12754] <= 32'b00000000010000010000000100010011;
ROM[12755] <= 32'b00000001010000000000001110010011;
ROM[12756] <= 32'b00000000100000111000001110010011;
ROM[12757] <= 32'b01000000011100010000001110110011;
ROM[12758] <= 32'b00000000011100000000001000110011;
ROM[12759] <= 32'b00000000001000000000000110110011;
ROM[12760] <= 32'b01000100110000011101000011101111;
ROM[12761] <= 32'b00000111010000000000001110010011;
ROM[12762] <= 32'b00000000011100010010000000100011;
ROM[12763] <= 32'b00000000010000010000000100010011;
ROM[12764] <= 32'b00000000000000001100001110110111;
ROM[12765] <= 32'b01111011110000111000001110010011;
ROM[12766] <= 32'b00000000111000111000001110110011;
ROM[12767] <= 32'b00000000011100010010000000100011;
ROM[12768] <= 32'b00000000010000010000000100010011;
ROM[12769] <= 32'b00000000001100010010000000100011;
ROM[12770] <= 32'b00000000010000010000000100010011;
ROM[12771] <= 32'b00000000010000010010000000100011;
ROM[12772] <= 32'b00000000010000010000000100010011;
ROM[12773] <= 32'b00000000010100010010000000100011;
ROM[12774] <= 32'b00000000010000010000000100010011;
ROM[12775] <= 32'b00000000011000010010000000100011;
ROM[12776] <= 32'b00000000010000010000000100010011;
ROM[12777] <= 32'b00000001010000000000001110010011;
ROM[12778] <= 32'b00000000100000111000001110010011;
ROM[12779] <= 32'b01000000011100010000001110110011;
ROM[12780] <= 32'b00000000011100000000001000110011;
ROM[12781] <= 32'b00000000001000000000000110110011;
ROM[12782] <= 32'b00111111010000011101000011101111;
ROM[12783] <= 32'b00000111010000000000001110010011;
ROM[12784] <= 32'b00000000011100010010000000100011;
ROM[12785] <= 32'b00000000010000010000000100010011;
ROM[12786] <= 32'b00000000000000001101001110110111;
ROM[12787] <= 32'b10000001010000111000001110010011;
ROM[12788] <= 32'b00000000111000111000001110110011;
ROM[12789] <= 32'b00000000011100010010000000100011;
ROM[12790] <= 32'b00000000010000010000000100010011;
ROM[12791] <= 32'b00000000001100010010000000100011;
ROM[12792] <= 32'b00000000010000010000000100010011;
ROM[12793] <= 32'b00000000010000010010000000100011;
ROM[12794] <= 32'b00000000010000010000000100010011;
ROM[12795] <= 32'b00000000010100010010000000100011;
ROM[12796] <= 32'b00000000010000010000000100010011;
ROM[12797] <= 32'b00000000011000010010000000100011;
ROM[12798] <= 32'b00000000010000010000000100010011;
ROM[12799] <= 32'b00000001010000000000001110010011;
ROM[12800] <= 32'b00000000100000111000001110010011;
ROM[12801] <= 32'b01000000011100010000001110110011;
ROM[12802] <= 32'b00000000011100000000001000110011;
ROM[12803] <= 32'b00000000001000000000000110110011;
ROM[12804] <= 32'b00111001110000011101000011101111;
ROM[12805] <= 32'b00000110010100000000001110010011;
ROM[12806] <= 32'b00000000011100010010000000100011;
ROM[12807] <= 32'b00000000010000010000000100010011;
ROM[12808] <= 32'b00000000000000001101001110110111;
ROM[12809] <= 32'b10000110110000111000001110010011;
ROM[12810] <= 32'b00000000111000111000001110110011;
ROM[12811] <= 32'b00000000011100010010000000100011;
ROM[12812] <= 32'b00000000010000010000000100010011;
ROM[12813] <= 32'b00000000001100010010000000100011;
ROM[12814] <= 32'b00000000010000010000000100010011;
ROM[12815] <= 32'b00000000010000010010000000100011;
ROM[12816] <= 32'b00000000010000010000000100010011;
ROM[12817] <= 32'b00000000010100010010000000100011;
ROM[12818] <= 32'b00000000010000010000000100010011;
ROM[12819] <= 32'b00000000011000010010000000100011;
ROM[12820] <= 32'b00000000010000010000000100010011;
ROM[12821] <= 32'b00000001010000000000001110010011;
ROM[12822] <= 32'b00000000100000111000001110010011;
ROM[12823] <= 32'b01000000011100010000001110110011;
ROM[12824] <= 32'b00000000011100000000001000110011;
ROM[12825] <= 32'b00000000001000000000000110110011;
ROM[12826] <= 32'b00110100010000011101000011101111;
ROM[12827] <= 32'b00000111001000000000001110010011;
ROM[12828] <= 32'b00000000011100010010000000100011;
ROM[12829] <= 32'b00000000010000010000000100010011;
ROM[12830] <= 32'b00000000000000001101001110110111;
ROM[12831] <= 32'b10001100010000111000001110010011;
ROM[12832] <= 32'b00000000111000111000001110110011;
ROM[12833] <= 32'b00000000011100010010000000100011;
ROM[12834] <= 32'b00000000010000010000000100010011;
ROM[12835] <= 32'b00000000001100010010000000100011;
ROM[12836] <= 32'b00000000010000010000000100010011;
ROM[12837] <= 32'b00000000010000010010000000100011;
ROM[12838] <= 32'b00000000010000010000000100010011;
ROM[12839] <= 32'b00000000010100010010000000100011;
ROM[12840] <= 32'b00000000010000010000000100010011;
ROM[12841] <= 32'b00000000011000010010000000100011;
ROM[12842] <= 32'b00000000010000010000000100010011;
ROM[12843] <= 32'b00000001010000000000001110010011;
ROM[12844] <= 32'b00000000100000111000001110010011;
ROM[12845] <= 32'b01000000011100010000001110110011;
ROM[12846] <= 32'b00000000011100000000001000110011;
ROM[12847] <= 32'b00000000001000000000000110110011;
ROM[12848] <= 32'b00101110110000011101000011101111;
ROM[12849] <= 32'b00000010000000000000001110010011;
ROM[12850] <= 32'b00000000011100010010000000100011;
ROM[12851] <= 32'b00000000010000010000000100010011;
ROM[12852] <= 32'b00000000000000001101001110110111;
ROM[12853] <= 32'b10010001110000111000001110010011;
ROM[12854] <= 32'b00000000111000111000001110110011;
ROM[12855] <= 32'b00000000011100010010000000100011;
ROM[12856] <= 32'b00000000010000010000000100010011;
ROM[12857] <= 32'b00000000001100010010000000100011;
ROM[12858] <= 32'b00000000010000010000000100010011;
ROM[12859] <= 32'b00000000010000010010000000100011;
ROM[12860] <= 32'b00000000010000010000000100010011;
ROM[12861] <= 32'b00000000010100010010000000100011;
ROM[12862] <= 32'b00000000010000010000000100010011;
ROM[12863] <= 32'b00000000011000010010000000100011;
ROM[12864] <= 32'b00000000010000010000000100010011;
ROM[12865] <= 32'b00000001010000000000001110010011;
ROM[12866] <= 32'b00000000100000111000001110010011;
ROM[12867] <= 32'b01000000011100010000001110110011;
ROM[12868] <= 32'b00000000011100000000001000110011;
ROM[12869] <= 32'b00000000001000000000000110110011;
ROM[12870] <= 32'b00101001010000011101000011101111;
ROM[12871] <= 32'b00000110000100000000001110010011;
ROM[12872] <= 32'b00000000011100010010000000100011;
ROM[12873] <= 32'b00000000010000010000000100010011;
ROM[12874] <= 32'b00000000000000001101001110110111;
ROM[12875] <= 32'b10010111010000111000001110010011;
ROM[12876] <= 32'b00000000111000111000001110110011;
ROM[12877] <= 32'b00000000011100010010000000100011;
ROM[12878] <= 32'b00000000010000010000000100010011;
ROM[12879] <= 32'b00000000001100010010000000100011;
ROM[12880] <= 32'b00000000010000010000000100010011;
ROM[12881] <= 32'b00000000010000010010000000100011;
ROM[12882] <= 32'b00000000010000010000000100010011;
ROM[12883] <= 32'b00000000010100010010000000100011;
ROM[12884] <= 32'b00000000010000010000000100010011;
ROM[12885] <= 32'b00000000011000010010000000100011;
ROM[12886] <= 32'b00000000010000010000000100010011;
ROM[12887] <= 32'b00000001010000000000001110010011;
ROM[12888] <= 32'b00000000100000111000001110010011;
ROM[12889] <= 32'b01000000011100010000001110110011;
ROM[12890] <= 32'b00000000011100000000001000110011;
ROM[12891] <= 32'b00000000001000000000000110110011;
ROM[12892] <= 32'b00100011110000011101000011101111;
ROM[12893] <= 32'b00000110110000000000001110010011;
ROM[12894] <= 32'b00000000011100010010000000100011;
ROM[12895] <= 32'b00000000010000010000000100010011;
ROM[12896] <= 32'b00000000000000001101001110110111;
ROM[12897] <= 32'b10011100110000111000001110010011;
ROM[12898] <= 32'b00000000111000111000001110110011;
ROM[12899] <= 32'b00000000011100010010000000100011;
ROM[12900] <= 32'b00000000010000010000000100010011;
ROM[12901] <= 32'b00000000001100010010000000100011;
ROM[12902] <= 32'b00000000010000010000000100010011;
ROM[12903] <= 32'b00000000010000010010000000100011;
ROM[12904] <= 32'b00000000010000010000000100010011;
ROM[12905] <= 32'b00000000010100010010000000100011;
ROM[12906] <= 32'b00000000010000010000000100010011;
ROM[12907] <= 32'b00000000011000010010000000100011;
ROM[12908] <= 32'b00000000010000010000000100010011;
ROM[12909] <= 32'b00000001010000000000001110010011;
ROM[12910] <= 32'b00000000100000111000001110010011;
ROM[12911] <= 32'b01000000011100010000001110110011;
ROM[12912] <= 32'b00000000011100000000001000110011;
ROM[12913] <= 32'b00000000001000000000000110110011;
ROM[12914] <= 32'b00011110010000011101000011101111;
ROM[12915] <= 32'b00000111001000000000001110010011;
ROM[12916] <= 32'b00000000011100010010000000100011;
ROM[12917] <= 32'b00000000010000010000000100010011;
ROM[12918] <= 32'b00000000000000001101001110110111;
ROM[12919] <= 32'b10100010010000111000001110010011;
ROM[12920] <= 32'b00000000111000111000001110110011;
ROM[12921] <= 32'b00000000011100010010000000100011;
ROM[12922] <= 32'b00000000010000010000000100010011;
ROM[12923] <= 32'b00000000001100010010000000100011;
ROM[12924] <= 32'b00000000010000010000000100010011;
ROM[12925] <= 32'b00000000010000010010000000100011;
ROM[12926] <= 32'b00000000010000010000000100010011;
ROM[12927] <= 32'b00000000010100010010000000100011;
ROM[12928] <= 32'b00000000010000010000000100010011;
ROM[12929] <= 32'b00000000011000010010000000100011;
ROM[12930] <= 32'b00000000010000010000000100010011;
ROM[12931] <= 32'b00000001010000000000001110010011;
ROM[12932] <= 32'b00000000100000111000001110010011;
ROM[12933] <= 32'b01000000011100010000001110110011;
ROM[12934] <= 32'b00000000011100000000001000110011;
ROM[12935] <= 32'b00000000001000000000000110110011;
ROM[12936] <= 32'b00011000110000011101000011101111;
ROM[12937] <= 32'b00000110010100000000001110010011;
ROM[12938] <= 32'b00000000011100010010000000100011;
ROM[12939] <= 32'b00000000010000010000000100010011;
ROM[12940] <= 32'b00000000000000001101001110110111;
ROM[12941] <= 32'b10100111110000111000001110010011;
ROM[12942] <= 32'b00000000111000111000001110110011;
ROM[12943] <= 32'b00000000011100010010000000100011;
ROM[12944] <= 32'b00000000010000010000000100010011;
ROM[12945] <= 32'b00000000001100010010000000100011;
ROM[12946] <= 32'b00000000010000010000000100010011;
ROM[12947] <= 32'b00000000010000010010000000100011;
ROM[12948] <= 32'b00000000010000010000000100010011;
ROM[12949] <= 32'b00000000010100010010000000100011;
ROM[12950] <= 32'b00000000010000010000000100010011;
ROM[12951] <= 32'b00000000011000010010000000100011;
ROM[12952] <= 32'b00000000010000010000000100010011;
ROM[12953] <= 32'b00000001010000000000001110010011;
ROM[12954] <= 32'b00000000100000111000001110010011;
ROM[12955] <= 32'b01000000011100010000001110110011;
ROM[12956] <= 32'b00000000011100000000001000110011;
ROM[12957] <= 32'b00000000001000000000000110110011;
ROM[12958] <= 32'b00010011010000011101000011101111;
ROM[12959] <= 32'b00000110000100000000001110010011;
ROM[12960] <= 32'b00000000011100010010000000100011;
ROM[12961] <= 32'b00000000010000010000000100010011;
ROM[12962] <= 32'b00000000000000001101001110110111;
ROM[12963] <= 32'b10101101010000111000001110010011;
ROM[12964] <= 32'b00000000111000111000001110110011;
ROM[12965] <= 32'b00000000011100010010000000100011;
ROM[12966] <= 32'b00000000010000010000000100010011;
ROM[12967] <= 32'b00000000001100010010000000100011;
ROM[12968] <= 32'b00000000010000010000000100010011;
ROM[12969] <= 32'b00000000010000010010000000100011;
ROM[12970] <= 32'b00000000010000010000000100010011;
ROM[12971] <= 32'b00000000010100010010000000100011;
ROM[12972] <= 32'b00000000010000010000000100010011;
ROM[12973] <= 32'b00000000011000010010000000100011;
ROM[12974] <= 32'b00000000010000010000000100010011;
ROM[12975] <= 32'b00000001010000000000001110010011;
ROM[12976] <= 32'b00000000100000111000001110010011;
ROM[12977] <= 32'b01000000011100010000001110110011;
ROM[12978] <= 32'b00000000011100000000001000110011;
ROM[12979] <= 32'b00000000001000000000000110110011;
ROM[12980] <= 32'b00001101110000011101000011101111;
ROM[12981] <= 32'b00000110010000000000001110010011;
ROM[12982] <= 32'b00000000011100010010000000100011;
ROM[12983] <= 32'b00000000010000010000000100010011;
ROM[12984] <= 32'b00000000000000001101001110110111;
ROM[12985] <= 32'b10110010110000111000001110010011;
ROM[12986] <= 32'b00000000111000111000001110110011;
ROM[12987] <= 32'b00000000011100010010000000100011;
ROM[12988] <= 32'b00000000010000010000000100010011;
ROM[12989] <= 32'b00000000001100010010000000100011;
ROM[12990] <= 32'b00000000010000010000000100010011;
ROM[12991] <= 32'b00000000010000010010000000100011;
ROM[12992] <= 32'b00000000010000010000000100010011;
ROM[12993] <= 32'b00000000010100010010000000100011;
ROM[12994] <= 32'b00000000010000010000000100010011;
ROM[12995] <= 32'b00000000011000010010000000100011;
ROM[12996] <= 32'b00000000010000010000000100010011;
ROM[12997] <= 32'b00000001010000000000001110010011;
ROM[12998] <= 32'b00000000100000111000001110010011;
ROM[12999] <= 32'b01000000011100010000001110110011;
ROM[13000] <= 32'b00000000011100000000001000110011;
ROM[13001] <= 32'b00000000001000000000000110110011;
ROM[13002] <= 32'b00001000010000011101000011101111;
ROM[13003] <= 32'b00000111100100000000001110010011;
ROM[13004] <= 32'b00000000011100010010000000100011;
ROM[13005] <= 32'b00000000010000010000000100010011;
ROM[13006] <= 32'b00000000000000001101001110110111;
ROM[13007] <= 32'b10111000010000111000001110010011;
ROM[13008] <= 32'b00000000111000111000001110110011;
ROM[13009] <= 32'b00000000011100010010000000100011;
ROM[13010] <= 32'b00000000010000010000000100010011;
ROM[13011] <= 32'b00000000001100010010000000100011;
ROM[13012] <= 32'b00000000010000010000000100010011;
ROM[13013] <= 32'b00000000010000010010000000100011;
ROM[13014] <= 32'b00000000010000010000000100010011;
ROM[13015] <= 32'b00000000010100010010000000100011;
ROM[13016] <= 32'b00000000010000010000000100010011;
ROM[13017] <= 32'b00000000011000010010000000100011;
ROM[13018] <= 32'b00000000010000010000000100010011;
ROM[13019] <= 32'b00000001010000000000001110010011;
ROM[13020] <= 32'b00000000100000111000001110010011;
ROM[13021] <= 32'b01000000011100010000001110110011;
ROM[13022] <= 32'b00000000011100000000001000110011;
ROM[13023] <= 32'b00000000001000000000000110110011;
ROM[13024] <= 32'b00000010110000011101000011101111;
ROM[13025] <= 32'b00000010000000000000001110010011;
ROM[13026] <= 32'b00000000011100010010000000100011;
ROM[13027] <= 32'b00000000010000010000000100010011;
ROM[13028] <= 32'b00000000000000001101001110110111;
ROM[13029] <= 32'b10111101110000111000001110010011;
ROM[13030] <= 32'b00000000111000111000001110110011;
ROM[13031] <= 32'b00000000011100010010000000100011;
ROM[13032] <= 32'b00000000010000010000000100010011;
ROM[13033] <= 32'b00000000001100010010000000100011;
ROM[13034] <= 32'b00000000010000010000000100010011;
ROM[13035] <= 32'b00000000010000010010000000100011;
ROM[13036] <= 32'b00000000010000010000000100010011;
ROM[13037] <= 32'b00000000010100010010000000100011;
ROM[13038] <= 32'b00000000010000010000000100010011;
ROM[13039] <= 32'b00000000011000010010000000100011;
ROM[13040] <= 32'b00000000010000010000000100010011;
ROM[13041] <= 32'b00000001010000000000001110010011;
ROM[13042] <= 32'b00000000100000111000001110010011;
ROM[13043] <= 32'b01000000011100010000001110110011;
ROM[13044] <= 32'b00000000011100000000001000110011;
ROM[13045] <= 32'b00000000001000000000000110110011;
ROM[13046] <= 32'b01111101010100011100000011101111;
ROM[13047] <= 32'b00000110011100000000001110010011;
ROM[13048] <= 32'b00000000011100010010000000100011;
ROM[13049] <= 32'b00000000010000010000000100010011;
ROM[13050] <= 32'b00000000000000001101001110110111;
ROM[13051] <= 32'b11000011010000111000001110010011;
ROM[13052] <= 32'b00000000111000111000001110110011;
ROM[13053] <= 32'b00000000011100010010000000100011;
ROM[13054] <= 32'b00000000010000010000000100010011;
ROM[13055] <= 32'b00000000001100010010000000100011;
ROM[13056] <= 32'b00000000010000010000000100010011;
ROM[13057] <= 32'b00000000010000010010000000100011;
ROM[13058] <= 32'b00000000010000010000000100010011;
ROM[13059] <= 32'b00000000010100010010000000100011;
ROM[13060] <= 32'b00000000010000010000000100010011;
ROM[13061] <= 32'b00000000011000010010000000100011;
ROM[13062] <= 32'b00000000010000010000000100010011;
ROM[13063] <= 32'b00000001010000000000001110010011;
ROM[13064] <= 32'b00000000100000111000001110010011;
ROM[13065] <= 32'b01000000011100010000001110110011;
ROM[13066] <= 32'b00000000011100000000001000110011;
ROM[13067] <= 32'b00000000001000000000000110110011;
ROM[13068] <= 32'b01110111110100011100000011101111;
ROM[13069] <= 32'b00000111010100000000001110010011;
ROM[13070] <= 32'b00000000011100010010000000100011;
ROM[13071] <= 32'b00000000010000010000000100010011;
ROM[13072] <= 32'b00000000000000001101001110110111;
ROM[13073] <= 32'b11001000110000111000001110010011;
ROM[13074] <= 32'b00000000111000111000001110110011;
ROM[13075] <= 32'b00000000011100010010000000100011;
ROM[13076] <= 32'b00000000010000010000000100010011;
ROM[13077] <= 32'b00000000001100010010000000100011;
ROM[13078] <= 32'b00000000010000010000000100010011;
ROM[13079] <= 32'b00000000010000010010000000100011;
ROM[13080] <= 32'b00000000010000010000000100010011;
ROM[13081] <= 32'b00000000010100010010000000100011;
ROM[13082] <= 32'b00000000010000010000000100010011;
ROM[13083] <= 32'b00000000011000010010000000100011;
ROM[13084] <= 32'b00000000010000010000000100010011;
ROM[13085] <= 32'b00000001010000000000001110010011;
ROM[13086] <= 32'b00000000100000111000001110010011;
ROM[13087] <= 32'b01000000011100010000001110110011;
ROM[13088] <= 32'b00000000011100000000001000110011;
ROM[13089] <= 32'b00000000001000000000000110110011;
ROM[13090] <= 32'b01110010010100011100000011101111;
ROM[13091] <= 32'b00000110010100000000001110010011;
ROM[13092] <= 32'b00000000011100010010000000100011;
ROM[13093] <= 32'b00000000010000010000000100010011;
ROM[13094] <= 32'b00000000000000001101001110110111;
ROM[13095] <= 32'b11001110010000111000001110010011;
ROM[13096] <= 32'b00000000111000111000001110110011;
ROM[13097] <= 32'b00000000011100010010000000100011;
ROM[13098] <= 32'b00000000010000010000000100010011;
ROM[13099] <= 32'b00000000001100010010000000100011;
ROM[13100] <= 32'b00000000010000010000000100010011;
ROM[13101] <= 32'b00000000010000010010000000100011;
ROM[13102] <= 32'b00000000010000010000000100010011;
ROM[13103] <= 32'b00000000010100010010000000100011;
ROM[13104] <= 32'b00000000010000010000000100010011;
ROM[13105] <= 32'b00000000011000010010000000100011;
ROM[13106] <= 32'b00000000010000010000000100010011;
ROM[13107] <= 32'b00000001010000000000001110010011;
ROM[13108] <= 32'b00000000100000111000001110010011;
ROM[13109] <= 32'b01000000011100010000001110110011;
ROM[13110] <= 32'b00000000011100000000001000110011;
ROM[13111] <= 32'b00000000001000000000000110110011;
ROM[13112] <= 32'b01101100110100011100000011101111;
ROM[13113] <= 32'b00000111001100000000001110010011;
ROM[13114] <= 32'b00000000011100010010000000100011;
ROM[13115] <= 32'b00000000010000010000000100010011;
ROM[13116] <= 32'b00000000000000001101001110110111;
ROM[13117] <= 32'b11010011110000111000001110010011;
ROM[13118] <= 32'b00000000111000111000001110110011;
ROM[13119] <= 32'b00000000011100010010000000100011;
ROM[13120] <= 32'b00000000010000010000000100010011;
ROM[13121] <= 32'b00000000001100010010000000100011;
ROM[13122] <= 32'b00000000010000010000000100010011;
ROM[13123] <= 32'b00000000010000010010000000100011;
ROM[13124] <= 32'b00000000010000010000000100010011;
ROM[13125] <= 32'b00000000010100010010000000100011;
ROM[13126] <= 32'b00000000010000010000000100010011;
ROM[13127] <= 32'b00000000011000010010000000100011;
ROM[13128] <= 32'b00000000010000010000000100010011;
ROM[13129] <= 32'b00000001010000000000001110010011;
ROM[13130] <= 32'b00000000100000111000001110010011;
ROM[13131] <= 32'b01000000011100010000001110110011;
ROM[13132] <= 32'b00000000011100000000001000110011;
ROM[13133] <= 32'b00000000001000000000000110110011;
ROM[13134] <= 32'b01100111010100011100000011101111;
ROM[13135] <= 32'b00000111001100000000001110010011;
ROM[13136] <= 32'b00000000011100010010000000100011;
ROM[13137] <= 32'b00000000010000010000000100010011;
ROM[13138] <= 32'b00000000000000001101001110110111;
ROM[13139] <= 32'b11011001010000111000001110010011;
ROM[13140] <= 32'b00000000111000111000001110110011;
ROM[13141] <= 32'b00000000011100010010000000100011;
ROM[13142] <= 32'b00000000010000010000000100010011;
ROM[13143] <= 32'b00000000001100010010000000100011;
ROM[13144] <= 32'b00000000010000010000000100010011;
ROM[13145] <= 32'b00000000010000010010000000100011;
ROM[13146] <= 32'b00000000010000010000000100010011;
ROM[13147] <= 32'b00000000010100010010000000100011;
ROM[13148] <= 32'b00000000010000010000000100010011;
ROM[13149] <= 32'b00000000011000010010000000100011;
ROM[13150] <= 32'b00000000010000010000000100010011;
ROM[13151] <= 32'b00000001010000000000001110010011;
ROM[13152] <= 32'b00000000100000111000001110010011;
ROM[13153] <= 32'b01000000011100010000001110110011;
ROM[13154] <= 32'b00000000011100000000001000110011;
ROM[13155] <= 32'b00000000001000000000000110110011;
ROM[13156] <= 32'b01100001110100011100000011101111;
ROM[13157] <= 32'b00000110010100000000001110010011;
ROM[13158] <= 32'b00000000011100010010000000100011;
ROM[13159] <= 32'b00000000010000010000000100010011;
ROM[13160] <= 32'b00000000000000001101001110110111;
ROM[13161] <= 32'b11011110110000111000001110010011;
ROM[13162] <= 32'b00000000111000111000001110110011;
ROM[13163] <= 32'b00000000011100010010000000100011;
ROM[13164] <= 32'b00000000010000010000000100010011;
ROM[13165] <= 32'b00000000001100010010000000100011;
ROM[13166] <= 32'b00000000010000010000000100010011;
ROM[13167] <= 32'b00000000010000010010000000100011;
ROM[13168] <= 32'b00000000010000010000000100010011;
ROM[13169] <= 32'b00000000010100010010000000100011;
ROM[13170] <= 32'b00000000010000010000000100010011;
ROM[13171] <= 32'b00000000011000010010000000100011;
ROM[13172] <= 32'b00000000010000010000000100010011;
ROM[13173] <= 32'b00000001010000000000001110010011;
ROM[13174] <= 32'b00000000100000111000001110010011;
ROM[13175] <= 32'b01000000011100010000001110110011;
ROM[13176] <= 32'b00000000011100000000001000110011;
ROM[13177] <= 32'b00000000001000000000000110110011;
ROM[13178] <= 32'b01011100010100011100000011101111;
ROM[13179] <= 32'b00000110010000000000001110010011;
ROM[13180] <= 32'b00000000011100010010000000100011;
ROM[13181] <= 32'b00000000010000010000000100010011;
ROM[13182] <= 32'b00000000000000001101001110110111;
ROM[13183] <= 32'b11100100010000111000001110010011;
ROM[13184] <= 32'b00000000111000111000001110110011;
ROM[13185] <= 32'b00000000011100010010000000100011;
ROM[13186] <= 32'b00000000010000010000000100010011;
ROM[13187] <= 32'b00000000001100010010000000100011;
ROM[13188] <= 32'b00000000010000010000000100010011;
ROM[13189] <= 32'b00000000010000010010000000100011;
ROM[13190] <= 32'b00000000010000010000000100010011;
ROM[13191] <= 32'b00000000010100010010000000100011;
ROM[13192] <= 32'b00000000010000010000000100010011;
ROM[13193] <= 32'b00000000011000010010000000100011;
ROM[13194] <= 32'b00000000010000010000000100010011;
ROM[13195] <= 32'b00000001010000000000001110010011;
ROM[13196] <= 32'b00000000100000111000001110010011;
ROM[13197] <= 32'b01000000011100010000001110110011;
ROM[13198] <= 32'b00000000011100000000001000110011;
ROM[13199] <= 32'b00000000001000000000000110110011;
ROM[13200] <= 32'b01010110110100011100000011101111;
ROM[13201] <= 32'b00000010110000000000001110010011;
ROM[13202] <= 32'b00000000011100010010000000100011;
ROM[13203] <= 32'b00000000010000010000000100010011;
ROM[13204] <= 32'b00000000000000001101001110110111;
ROM[13205] <= 32'b11101001110000111000001110010011;
ROM[13206] <= 32'b00000000111000111000001110110011;
ROM[13207] <= 32'b00000000011100010010000000100011;
ROM[13208] <= 32'b00000000010000010000000100010011;
ROM[13209] <= 32'b00000000001100010010000000100011;
ROM[13210] <= 32'b00000000010000010000000100010011;
ROM[13211] <= 32'b00000000010000010010000000100011;
ROM[13212] <= 32'b00000000010000010000000100010011;
ROM[13213] <= 32'b00000000010100010010000000100011;
ROM[13214] <= 32'b00000000010000010000000100010011;
ROM[13215] <= 32'b00000000011000010010000000100011;
ROM[13216] <= 32'b00000000010000010000000100010011;
ROM[13217] <= 32'b00000001010000000000001110010011;
ROM[13218] <= 32'b00000000100000111000001110010011;
ROM[13219] <= 32'b01000000011100010000001110110011;
ROM[13220] <= 32'b00000000011100000000001000110011;
ROM[13221] <= 32'b00000000001000000000000110110011;
ROM[13222] <= 32'b01010001010100011100000011101111;
ROM[13223] <= 32'b00000010000000000000001110010011;
ROM[13224] <= 32'b00000000011100010010000000100011;
ROM[13225] <= 32'b00000000010000010000000100010011;
ROM[13226] <= 32'b00000000000000001101001110110111;
ROM[13227] <= 32'b11101111010000111000001110010011;
ROM[13228] <= 32'b00000000111000111000001110110011;
ROM[13229] <= 32'b00000000011100010010000000100011;
ROM[13230] <= 32'b00000000010000010000000100010011;
ROM[13231] <= 32'b00000000001100010010000000100011;
ROM[13232] <= 32'b00000000010000010000000100010011;
ROM[13233] <= 32'b00000000010000010010000000100011;
ROM[13234] <= 32'b00000000010000010000000100010011;
ROM[13235] <= 32'b00000000010100010010000000100011;
ROM[13236] <= 32'b00000000010000010000000100010011;
ROM[13237] <= 32'b00000000011000010010000000100011;
ROM[13238] <= 32'b00000000010000010000000100010011;
ROM[13239] <= 32'b00000001010000000000001110010011;
ROM[13240] <= 32'b00000000100000111000001110010011;
ROM[13241] <= 32'b01000000011100010000001110110011;
ROM[13242] <= 32'b00000000011100000000001000110011;
ROM[13243] <= 32'b00000000001000000000000110110011;
ROM[13244] <= 32'b01001011110100011100000011101111;
ROM[13245] <= 32'b00000110011100000000001110010011;
ROM[13246] <= 32'b00000000011100010010000000100011;
ROM[13247] <= 32'b00000000010000010000000100010011;
ROM[13248] <= 32'b00000000000000001101001110110111;
ROM[13249] <= 32'b11110100110000111000001110010011;
ROM[13250] <= 32'b00000000111000111000001110110011;
ROM[13251] <= 32'b00000000011100010010000000100011;
ROM[13252] <= 32'b00000000010000010000000100010011;
ROM[13253] <= 32'b00000000001100010010000000100011;
ROM[13254] <= 32'b00000000010000010000000100010011;
ROM[13255] <= 32'b00000000010000010010000000100011;
ROM[13256] <= 32'b00000000010000010000000100010011;
ROM[13257] <= 32'b00000000010100010010000000100011;
ROM[13258] <= 32'b00000000010000010000000100010011;
ROM[13259] <= 32'b00000000011000010010000000100011;
ROM[13260] <= 32'b00000000010000010000000100010011;
ROM[13261] <= 32'b00000001010000000000001110010011;
ROM[13262] <= 32'b00000000100000111000001110010011;
ROM[13263] <= 32'b01000000011100010000001110110011;
ROM[13264] <= 32'b00000000011100000000001000110011;
ROM[13265] <= 32'b00000000001000000000000110110011;
ROM[13266] <= 32'b01000110010100011100000011101111;
ROM[13267] <= 32'b00000111010100000000001110010011;
ROM[13268] <= 32'b00000000011100010010000000100011;
ROM[13269] <= 32'b00000000010000010000000100010011;
ROM[13270] <= 32'b00000000000000001101001110110111;
ROM[13271] <= 32'b11111010010000111000001110010011;
ROM[13272] <= 32'b00000000111000111000001110110011;
ROM[13273] <= 32'b00000000011100010010000000100011;
ROM[13274] <= 32'b00000000010000010000000100010011;
ROM[13275] <= 32'b00000000001100010010000000100011;
ROM[13276] <= 32'b00000000010000010000000100010011;
ROM[13277] <= 32'b00000000010000010010000000100011;
ROM[13278] <= 32'b00000000010000010000000100010011;
ROM[13279] <= 32'b00000000010100010010000000100011;
ROM[13280] <= 32'b00000000010000010000000100010011;
ROM[13281] <= 32'b00000000011000010010000000100011;
ROM[13282] <= 32'b00000000010000010000000100010011;
ROM[13283] <= 32'b00000001010000000000001110010011;
ROM[13284] <= 32'b00000000100000111000001110010011;
ROM[13285] <= 32'b01000000011100010000001110110011;
ROM[13286] <= 32'b00000000011100000000001000110011;
ROM[13287] <= 32'b00000000001000000000000110110011;
ROM[13288] <= 32'b01000000110100011100000011101111;
ROM[13289] <= 32'b00000110010100000000001110010011;
ROM[13290] <= 32'b00000000011100010010000000100011;
ROM[13291] <= 32'b00000000010000010000000100010011;
ROM[13292] <= 32'b00000000000000001101001110110111;
ROM[13293] <= 32'b11111111110000111000001110010011;
ROM[13294] <= 32'b00000000111000111000001110110011;
ROM[13295] <= 32'b00000000011100010010000000100011;
ROM[13296] <= 32'b00000000010000010000000100010011;
ROM[13297] <= 32'b00000000001100010010000000100011;
ROM[13298] <= 32'b00000000010000010000000100010011;
ROM[13299] <= 32'b00000000010000010010000000100011;
ROM[13300] <= 32'b00000000010000010000000100010011;
ROM[13301] <= 32'b00000000010100010010000000100011;
ROM[13302] <= 32'b00000000010000010000000100010011;
ROM[13303] <= 32'b00000000011000010010000000100011;
ROM[13304] <= 32'b00000000010000010000000100010011;
ROM[13305] <= 32'b00000001010000000000001110010011;
ROM[13306] <= 32'b00000000100000111000001110010011;
ROM[13307] <= 32'b01000000011100010000001110110011;
ROM[13308] <= 32'b00000000011100000000001000110011;
ROM[13309] <= 32'b00000000001000000000000110110011;
ROM[13310] <= 32'b00111011010100011100000011101111;
ROM[13311] <= 32'b00000111001100000000001110010011;
ROM[13312] <= 32'b00000000011100010010000000100011;
ROM[13313] <= 32'b00000000010000010000000100010011;
ROM[13314] <= 32'b00000000000000001101001110110111;
ROM[13315] <= 32'b00000101010000111000001110010011;
ROM[13316] <= 32'b00000000111000111000001110110011;
ROM[13317] <= 32'b00000000011100010010000000100011;
ROM[13318] <= 32'b00000000010000010000000100010011;
ROM[13319] <= 32'b00000000001100010010000000100011;
ROM[13320] <= 32'b00000000010000010000000100010011;
ROM[13321] <= 32'b00000000010000010010000000100011;
ROM[13322] <= 32'b00000000010000010000000100010011;
ROM[13323] <= 32'b00000000010100010010000000100011;
ROM[13324] <= 32'b00000000010000010000000100010011;
ROM[13325] <= 32'b00000000011000010010000000100011;
ROM[13326] <= 32'b00000000010000010000000100010011;
ROM[13327] <= 32'b00000001010000000000001110010011;
ROM[13328] <= 32'b00000000100000111000001110010011;
ROM[13329] <= 32'b01000000011100010000001110110011;
ROM[13330] <= 32'b00000000011100000000001000110011;
ROM[13331] <= 32'b00000000001000000000000110110011;
ROM[13332] <= 32'b00110101110100011100000011101111;
ROM[13333] <= 32'b00000111001100000000001110010011;
ROM[13334] <= 32'b00000000011100010010000000100011;
ROM[13335] <= 32'b00000000010000010000000100010011;
ROM[13336] <= 32'b00000000000000001101001110110111;
ROM[13337] <= 32'b00001010110000111000001110010011;
ROM[13338] <= 32'b00000000111000111000001110110011;
ROM[13339] <= 32'b00000000011100010010000000100011;
ROM[13340] <= 32'b00000000010000010000000100010011;
ROM[13341] <= 32'b00000000001100010010000000100011;
ROM[13342] <= 32'b00000000010000010000000100010011;
ROM[13343] <= 32'b00000000010000010010000000100011;
ROM[13344] <= 32'b00000000010000010000000100010011;
ROM[13345] <= 32'b00000000010100010010000000100011;
ROM[13346] <= 32'b00000000010000010000000100010011;
ROM[13347] <= 32'b00000000011000010010000000100011;
ROM[13348] <= 32'b00000000010000010000000100010011;
ROM[13349] <= 32'b00000001010000000000001110010011;
ROM[13350] <= 32'b00000000100000111000001110010011;
ROM[13351] <= 32'b01000000011100010000001110110011;
ROM[13352] <= 32'b00000000011100000000001000110011;
ROM[13353] <= 32'b00000000001000000000000110110011;
ROM[13354] <= 32'b00110000010100011100000011101111;
ROM[13355] <= 32'b00000010000000000000001110010011;
ROM[13356] <= 32'b00000000011100010010000000100011;
ROM[13357] <= 32'b00000000010000010000000100010011;
ROM[13358] <= 32'b00000000000000001101001110110111;
ROM[13359] <= 32'b00010000010000111000001110010011;
ROM[13360] <= 32'b00000000111000111000001110110011;
ROM[13361] <= 32'b00000000011100010010000000100011;
ROM[13362] <= 32'b00000000010000010000000100010011;
ROM[13363] <= 32'b00000000001100010010000000100011;
ROM[13364] <= 32'b00000000010000010000000100010011;
ROM[13365] <= 32'b00000000010000010010000000100011;
ROM[13366] <= 32'b00000000010000010000000100010011;
ROM[13367] <= 32'b00000000010100010010000000100011;
ROM[13368] <= 32'b00000000010000010000000100010011;
ROM[13369] <= 32'b00000000011000010010000000100011;
ROM[13370] <= 32'b00000000010000010000000100010011;
ROM[13371] <= 32'b00000001010000000000001110010011;
ROM[13372] <= 32'b00000000100000111000001110010011;
ROM[13373] <= 32'b01000000011100010000001110110011;
ROM[13374] <= 32'b00000000011100000000001000110011;
ROM[13375] <= 32'b00000000001000000000000110110011;
ROM[13376] <= 32'b00101010110100011100000011101111;
ROM[13377] <= 32'b00000110000100000000001110010011;
ROM[13378] <= 32'b00000000011100010010000000100011;
ROM[13379] <= 32'b00000000010000010000000100010011;
ROM[13380] <= 32'b00000000000000001101001110110111;
ROM[13381] <= 32'b00010101110000111000001110010011;
ROM[13382] <= 32'b00000000111000111000001110110011;
ROM[13383] <= 32'b00000000011100010010000000100011;
ROM[13384] <= 32'b00000000010000010000000100010011;
ROM[13385] <= 32'b00000000001100010010000000100011;
ROM[13386] <= 32'b00000000010000010000000100010011;
ROM[13387] <= 32'b00000000010000010010000000100011;
ROM[13388] <= 32'b00000000010000010000000100010011;
ROM[13389] <= 32'b00000000010100010010000000100011;
ROM[13390] <= 32'b00000000010000010000000100010011;
ROM[13391] <= 32'b00000000011000010010000000100011;
ROM[13392] <= 32'b00000000010000010000000100010011;
ROM[13393] <= 32'b00000001010000000000001110010011;
ROM[13394] <= 32'b00000000100000111000001110010011;
ROM[13395] <= 32'b01000000011100010000001110110011;
ROM[13396] <= 32'b00000000011100000000001000110011;
ROM[13397] <= 32'b00000000001000000000000110110011;
ROM[13398] <= 32'b00100101010100011100000011101111;
ROM[13399] <= 32'b00000110111000000000001110010011;
ROM[13400] <= 32'b00000000011100010010000000100011;
ROM[13401] <= 32'b00000000010000010000000100010011;
ROM[13402] <= 32'b00000000000000001101001110110111;
ROM[13403] <= 32'b00011011010000111000001110010011;
ROM[13404] <= 32'b00000000111000111000001110110011;
ROM[13405] <= 32'b00000000011100010010000000100011;
ROM[13406] <= 32'b00000000010000010000000100010011;
ROM[13407] <= 32'b00000000001100010010000000100011;
ROM[13408] <= 32'b00000000010000010000000100010011;
ROM[13409] <= 32'b00000000010000010010000000100011;
ROM[13410] <= 32'b00000000010000010000000100010011;
ROM[13411] <= 32'b00000000010100010010000000100011;
ROM[13412] <= 32'b00000000010000010000000100010011;
ROM[13413] <= 32'b00000000011000010010000000100011;
ROM[13414] <= 32'b00000000010000010000000100010011;
ROM[13415] <= 32'b00000001010000000000001110010011;
ROM[13416] <= 32'b00000000100000111000001110010011;
ROM[13417] <= 32'b01000000011100010000001110110011;
ROM[13418] <= 32'b00000000011100000000001000110011;
ROM[13419] <= 32'b00000000001000000000000110110011;
ROM[13420] <= 32'b00011111110100011100000011101111;
ROM[13421] <= 32'b00000110111100000000001110010011;
ROM[13422] <= 32'b00000000011100010010000000100011;
ROM[13423] <= 32'b00000000010000010000000100010011;
ROM[13424] <= 32'b00000000000000001101001110110111;
ROM[13425] <= 32'b00100000110000111000001110010011;
ROM[13426] <= 32'b00000000111000111000001110110011;
ROM[13427] <= 32'b00000000011100010010000000100011;
ROM[13428] <= 32'b00000000010000010000000100010011;
ROM[13429] <= 32'b00000000001100010010000000100011;
ROM[13430] <= 32'b00000000010000010000000100010011;
ROM[13431] <= 32'b00000000010000010010000000100011;
ROM[13432] <= 32'b00000000010000010000000100010011;
ROM[13433] <= 32'b00000000010100010010000000100011;
ROM[13434] <= 32'b00000000010000010000000100010011;
ROM[13435] <= 32'b00000000011000010010000000100011;
ROM[13436] <= 32'b00000000010000010000000100010011;
ROM[13437] <= 32'b00000001010000000000001110010011;
ROM[13438] <= 32'b00000000100000111000001110010011;
ROM[13439] <= 32'b01000000011100010000001110110011;
ROM[13440] <= 32'b00000000011100000000001000110011;
ROM[13441] <= 32'b00000000001000000000000110110011;
ROM[13442] <= 32'b00011010010100011100000011101111;
ROM[13443] <= 32'b00000111010000000000001110010011;
ROM[13444] <= 32'b00000000011100010010000000100011;
ROM[13445] <= 32'b00000000010000010000000100010011;
ROM[13446] <= 32'b00000000000000001101001110110111;
ROM[13447] <= 32'b00100110010000111000001110010011;
ROM[13448] <= 32'b00000000111000111000001110110011;
ROM[13449] <= 32'b00000000011100010010000000100011;
ROM[13450] <= 32'b00000000010000010000000100010011;
ROM[13451] <= 32'b00000000001100010010000000100011;
ROM[13452] <= 32'b00000000010000010000000100010011;
ROM[13453] <= 32'b00000000010000010010000000100011;
ROM[13454] <= 32'b00000000010000010000000100010011;
ROM[13455] <= 32'b00000000010100010010000000100011;
ROM[13456] <= 32'b00000000010000010000000100010011;
ROM[13457] <= 32'b00000000011000010010000000100011;
ROM[13458] <= 32'b00000000010000010000000100010011;
ROM[13459] <= 32'b00000001010000000000001110010011;
ROM[13460] <= 32'b00000000100000111000001110010011;
ROM[13461] <= 32'b01000000011100010000001110110011;
ROM[13462] <= 32'b00000000011100000000001000110011;
ROM[13463] <= 32'b00000000001000000000000110110011;
ROM[13464] <= 32'b00010100110100011100000011101111;
ROM[13465] <= 32'b00000110100000000000001110010011;
ROM[13466] <= 32'b00000000011100010010000000100011;
ROM[13467] <= 32'b00000000010000010000000100010011;
ROM[13468] <= 32'b00000000000000001101001110110111;
ROM[13469] <= 32'b00101011110000111000001110010011;
ROM[13470] <= 32'b00000000111000111000001110110011;
ROM[13471] <= 32'b00000000011100010010000000100011;
ROM[13472] <= 32'b00000000010000010000000100010011;
ROM[13473] <= 32'b00000000001100010010000000100011;
ROM[13474] <= 32'b00000000010000010000000100010011;
ROM[13475] <= 32'b00000000010000010010000000100011;
ROM[13476] <= 32'b00000000010000010000000100010011;
ROM[13477] <= 32'b00000000010100010010000000100011;
ROM[13478] <= 32'b00000000010000010000000100010011;
ROM[13479] <= 32'b00000000011000010010000000100011;
ROM[13480] <= 32'b00000000010000010000000100010011;
ROM[13481] <= 32'b00000001010000000000001110010011;
ROM[13482] <= 32'b00000000100000111000001110010011;
ROM[13483] <= 32'b01000000011100010000001110110011;
ROM[13484] <= 32'b00000000011100000000001000110011;
ROM[13485] <= 32'b00000000001000000000000110110011;
ROM[13486] <= 32'b00001111010100011100000011101111;
ROM[13487] <= 32'b00000110010100000000001110010011;
ROM[13488] <= 32'b00000000011100010010000000100011;
ROM[13489] <= 32'b00000000010000010000000100010011;
ROM[13490] <= 32'b00000000000000001101001110110111;
ROM[13491] <= 32'b00110001010000111000001110010011;
ROM[13492] <= 32'b00000000111000111000001110110011;
ROM[13493] <= 32'b00000000011100010010000000100011;
ROM[13494] <= 32'b00000000010000010000000100010011;
ROM[13495] <= 32'b00000000001100010010000000100011;
ROM[13496] <= 32'b00000000010000010000000100010011;
ROM[13497] <= 32'b00000000010000010010000000100011;
ROM[13498] <= 32'b00000000010000010000000100010011;
ROM[13499] <= 32'b00000000010100010010000000100011;
ROM[13500] <= 32'b00000000010000010000000100010011;
ROM[13501] <= 32'b00000000011000010010000000100011;
ROM[13502] <= 32'b00000000010000010000000100010011;
ROM[13503] <= 32'b00000001010000000000001110010011;
ROM[13504] <= 32'b00000000100000111000001110010011;
ROM[13505] <= 32'b01000000011100010000001110110011;
ROM[13506] <= 32'b00000000011100000000001000110011;
ROM[13507] <= 32'b00000000001000000000000110110011;
ROM[13508] <= 32'b00001001110100011100000011101111;
ROM[13509] <= 32'b00000111001000000000001110010011;
ROM[13510] <= 32'b00000000011100010010000000100011;
ROM[13511] <= 32'b00000000010000010000000100010011;
ROM[13512] <= 32'b00000000000000001101001110110111;
ROM[13513] <= 32'b00110110110000111000001110010011;
ROM[13514] <= 32'b00000000111000111000001110110011;
ROM[13515] <= 32'b00000000011100010010000000100011;
ROM[13516] <= 32'b00000000010000010000000100010011;
ROM[13517] <= 32'b00000000001100010010000000100011;
ROM[13518] <= 32'b00000000010000010000000100010011;
ROM[13519] <= 32'b00000000010000010010000000100011;
ROM[13520] <= 32'b00000000010000010000000100010011;
ROM[13521] <= 32'b00000000010100010010000000100011;
ROM[13522] <= 32'b00000000010000010000000100010011;
ROM[13523] <= 32'b00000000011000010010000000100011;
ROM[13524] <= 32'b00000000010000010000000100010011;
ROM[13525] <= 32'b00000001010000000000001110010011;
ROM[13526] <= 32'b00000000100000111000001110010011;
ROM[13527] <= 32'b01000000011100010000001110110011;
ROM[13528] <= 32'b00000000011100000000001000110011;
ROM[13529] <= 32'b00000000001000000000000110110011;
ROM[13530] <= 32'b00000100010100011100000011101111;
ROM[13531] <= 32'b00000010000000000000001110010011;
ROM[13532] <= 32'b00000000011100010010000000100011;
ROM[13533] <= 32'b00000000010000010000000100010011;
ROM[13534] <= 32'b00000000000000001101001110110111;
ROM[13535] <= 32'b00111100010000111000001110010011;
ROM[13536] <= 32'b00000000111000111000001110110011;
ROM[13537] <= 32'b00000000011100010010000000100011;
ROM[13538] <= 32'b00000000010000010000000100010011;
ROM[13539] <= 32'b00000000001100010010000000100011;
ROM[13540] <= 32'b00000000010000010000000100010011;
ROM[13541] <= 32'b00000000010000010010000000100011;
ROM[13542] <= 32'b00000000010000010000000100010011;
ROM[13543] <= 32'b00000000010100010010000000100011;
ROM[13544] <= 32'b00000000010000010000000100010011;
ROM[13545] <= 32'b00000000011000010010000000100011;
ROM[13546] <= 32'b00000000010000010000000100010011;
ROM[13547] <= 32'b00000001010000000000001110010011;
ROM[13548] <= 32'b00000000100000111000001110010011;
ROM[13549] <= 32'b01000000011100010000001110110011;
ROM[13550] <= 32'b00000000011100000000001000110011;
ROM[13551] <= 32'b00000000001000000000000110110011;
ROM[13552] <= 32'b01111110110000011100000011101111;
ROM[13553] <= 32'b00000110110000000000001110010011;
ROM[13554] <= 32'b00000000011100010010000000100011;
ROM[13555] <= 32'b00000000010000010000000100010011;
ROM[13556] <= 32'b00000000000000001101001110110111;
ROM[13557] <= 32'b01000001110000111000001110010011;
ROM[13558] <= 32'b00000000111000111000001110110011;
ROM[13559] <= 32'b00000000011100010010000000100011;
ROM[13560] <= 32'b00000000010000010000000100010011;
ROM[13561] <= 32'b00000000001100010010000000100011;
ROM[13562] <= 32'b00000000010000010000000100010011;
ROM[13563] <= 32'b00000000010000010010000000100011;
ROM[13564] <= 32'b00000000010000010000000100010011;
ROM[13565] <= 32'b00000000010100010010000000100011;
ROM[13566] <= 32'b00000000010000010000000100010011;
ROM[13567] <= 32'b00000000011000010010000000100011;
ROM[13568] <= 32'b00000000010000010000000100010011;
ROM[13569] <= 32'b00000001010000000000001110010011;
ROM[13570] <= 32'b00000000100000111000001110010011;
ROM[13571] <= 32'b01000000011100010000001110110011;
ROM[13572] <= 32'b00000000011100000000001000110011;
ROM[13573] <= 32'b00000000001000000000000110110011;
ROM[13574] <= 32'b01111001010000011100000011101111;
ROM[13575] <= 32'b00000110010100000000001110010011;
ROM[13576] <= 32'b00000000011100010010000000100011;
ROM[13577] <= 32'b00000000010000010000000100010011;
ROM[13578] <= 32'b00000000000000001101001110110111;
ROM[13579] <= 32'b01000111010000111000001110010011;
ROM[13580] <= 32'b00000000111000111000001110110011;
ROM[13581] <= 32'b00000000011100010010000000100011;
ROM[13582] <= 32'b00000000010000010000000100010011;
ROM[13583] <= 32'b00000000001100010010000000100011;
ROM[13584] <= 32'b00000000010000010000000100010011;
ROM[13585] <= 32'b00000000010000010010000000100011;
ROM[13586] <= 32'b00000000010000010000000100010011;
ROM[13587] <= 32'b00000000010100010010000000100011;
ROM[13588] <= 32'b00000000010000010000000100010011;
ROM[13589] <= 32'b00000000011000010010000000100011;
ROM[13590] <= 32'b00000000010000010000000100010011;
ROM[13591] <= 32'b00000001010000000000001110010011;
ROM[13592] <= 32'b00000000100000111000001110010011;
ROM[13593] <= 32'b01000000011100010000001110110011;
ROM[13594] <= 32'b00000000011100000000001000110011;
ROM[13595] <= 32'b00000000001000000000000110110011;
ROM[13596] <= 32'b01110011110000011100000011101111;
ROM[13597] <= 32'b00000111010000000000001110010011;
ROM[13598] <= 32'b00000000011100010010000000100011;
ROM[13599] <= 32'b00000000010000010000000100010011;
ROM[13600] <= 32'b00000000000000001101001110110111;
ROM[13601] <= 32'b01001100110000111000001110010011;
ROM[13602] <= 32'b00000000111000111000001110110011;
ROM[13603] <= 32'b00000000011100010010000000100011;
ROM[13604] <= 32'b00000000010000010000000100010011;
ROM[13605] <= 32'b00000000001100010010000000100011;
ROM[13606] <= 32'b00000000010000010000000100010011;
ROM[13607] <= 32'b00000000010000010010000000100011;
ROM[13608] <= 32'b00000000010000010000000100010011;
ROM[13609] <= 32'b00000000010100010010000000100011;
ROM[13610] <= 32'b00000000010000010000000100010011;
ROM[13611] <= 32'b00000000011000010010000000100011;
ROM[13612] <= 32'b00000000010000010000000100010011;
ROM[13613] <= 32'b00000001010000000000001110010011;
ROM[13614] <= 32'b00000000100000111000001110010011;
ROM[13615] <= 32'b01000000011100010000001110110011;
ROM[13616] <= 32'b00000000011100000000001000110011;
ROM[13617] <= 32'b00000000001000000000000110110011;
ROM[13618] <= 32'b01101110010000011100000011101111;
ROM[13619] <= 32'b00000111010000000000001110010011;
ROM[13620] <= 32'b00000000011100010010000000100011;
ROM[13621] <= 32'b00000000010000010000000100010011;
ROM[13622] <= 32'b00000000000000001101001110110111;
ROM[13623] <= 32'b01010010010000111000001110010011;
ROM[13624] <= 32'b00000000111000111000001110110011;
ROM[13625] <= 32'b00000000011100010010000000100011;
ROM[13626] <= 32'b00000000010000010000000100010011;
ROM[13627] <= 32'b00000000001100010010000000100011;
ROM[13628] <= 32'b00000000010000010000000100010011;
ROM[13629] <= 32'b00000000010000010010000000100011;
ROM[13630] <= 32'b00000000010000010000000100010011;
ROM[13631] <= 32'b00000000010100010010000000100011;
ROM[13632] <= 32'b00000000010000010000000100010011;
ROM[13633] <= 32'b00000000011000010010000000100011;
ROM[13634] <= 32'b00000000010000010000000100010011;
ROM[13635] <= 32'b00000001010000000000001110010011;
ROM[13636] <= 32'b00000000100000111000001110010011;
ROM[13637] <= 32'b01000000011100010000001110110011;
ROM[13638] <= 32'b00000000011100000000001000110011;
ROM[13639] <= 32'b00000000001000000000000110110011;
ROM[13640] <= 32'b01101000110000011100000011101111;
ROM[13641] <= 32'b00000110010100000000001110010011;
ROM[13642] <= 32'b00000000011100010010000000100011;
ROM[13643] <= 32'b00000000010000010000000100010011;
ROM[13644] <= 32'b00000000000000001101001110110111;
ROM[13645] <= 32'b01010111110000111000001110010011;
ROM[13646] <= 32'b00000000111000111000001110110011;
ROM[13647] <= 32'b00000000011100010010000000100011;
ROM[13648] <= 32'b00000000010000010000000100010011;
ROM[13649] <= 32'b00000000001100010010000000100011;
ROM[13650] <= 32'b00000000010000010000000100010011;
ROM[13651] <= 32'b00000000010000010010000000100011;
ROM[13652] <= 32'b00000000010000010000000100010011;
ROM[13653] <= 32'b00000000010100010010000000100011;
ROM[13654] <= 32'b00000000010000010000000100010011;
ROM[13655] <= 32'b00000000011000010010000000100011;
ROM[13656] <= 32'b00000000010000010000000100010011;
ROM[13657] <= 32'b00000001010000000000001110010011;
ROM[13658] <= 32'b00000000100000111000001110010011;
ROM[13659] <= 32'b01000000011100010000001110110011;
ROM[13660] <= 32'b00000000011100000000001000110011;
ROM[13661] <= 32'b00000000001000000000000110110011;
ROM[13662] <= 32'b01100011010000011100000011101111;
ROM[13663] <= 32'b00000111001000000000001110010011;
ROM[13664] <= 32'b00000000011100010010000000100011;
ROM[13665] <= 32'b00000000010000010000000100010011;
ROM[13666] <= 32'b00000000000000001101001110110111;
ROM[13667] <= 32'b01011101010000111000001110010011;
ROM[13668] <= 32'b00000000111000111000001110110011;
ROM[13669] <= 32'b00000000011100010010000000100011;
ROM[13670] <= 32'b00000000010000010000000100010011;
ROM[13671] <= 32'b00000000001100010010000000100011;
ROM[13672] <= 32'b00000000010000010000000100010011;
ROM[13673] <= 32'b00000000010000010010000000100011;
ROM[13674] <= 32'b00000000010000010000000100010011;
ROM[13675] <= 32'b00000000010100010010000000100011;
ROM[13676] <= 32'b00000000010000010000000100010011;
ROM[13677] <= 32'b00000000011000010010000000100011;
ROM[13678] <= 32'b00000000010000010000000100010011;
ROM[13679] <= 32'b00000001010000000000001110010011;
ROM[13680] <= 32'b00000000100000111000001110010011;
ROM[13681] <= 32'b01000000011100010000001110110011;
ROM[13682] <= 32'b00000000011100000000001000110011;
ROM[13683] <= 32'b00000000001000000000000110110011;
ROM[13684] <= 32'b01011101110000011100000011101111;
ROM[13685] <= 32'b00000000000000001101001110110111;
ROM[13686] <= 32'b01100010000000111000001110010011;
ROM[13687] <= 32'b00000000111000111000001110110011;
ROM[13688] <= 32'b00000000011100010010000000100011;
ROM[13689] <= 32'b00000000010000010000000100010011;
ROM[13690] <= 32'b00000000001100010010000000100011;
ROM[13691] <= 32'b00000000010000010000000100010011;
ROM[13692] <= 32'b00000000010000010010000000100011;
ROM[13693] <= 32'b00000000010000010000000100010011;
ROM[13694] <= 32'b00000000010100010010000000100011;
ROM[13695] <= 32'b00000000010000010000000100010011;
ROM[13696] <= 32'b00000000011000010010000000100011;
ROM[13697] <= 32'b00000000010000010000000100010011;
ROM[13698] <= 32'b00000001010000000000001110010011;
ROM[13699] <= 32'b00000000010000111000001110010011;
ROM[13700] <= 32'b01000000011100010000001110110011;
ROM[13701] <= 32'b00000000011100000000001000110011;
ROM[13702] <= 32'b00000000001000000000000110110011;
ROM[13703] <= 32'b00010100110100001001000011101111;
ROM[13704] <= 32'b11111111110000010000000100010011;
ROM[13705] <= 32'b00000000000000010010001110000011;
ROM[13706] <= 32'b00000000011101100010000000100011;
ROM[13707] <= 32'b00000000000000001101001110110111;
ROM[13708] <= 32'b01100111100000111000001110010011;
ROM[13709] <= 32'b00000000111000111000001110110011;
ROM[13710] <= 32'b00000000011100010010000000100011;
ROM[13711] <= 32'b00000000010000010000000100010011;
ROM[13712] <= 32'b00000000001100010010000000100011;
ROM[13713] <= 32'b00000000010000010000000100010011;
ROM[13714] <= 32'b00000000010000010010000000100011;
ROM[13715] <= 32'b00000000010000010000000100010011;
ROM[13716] <= 32'b00000000010100010010000000100011;
ROM[13717] <= 32'b00000000010000010000000100010011;
ROM[13718] <= 32'b00000000011000010010000000100011;
ROM[13719] <= 32'b00000000010000010000000100010011;
ROM[13720] <= 32'b00000001010000000000001110010011;
ROM[13721] <= 32'b00000000000000111000001110010011;
ROM[13722] <= 32'b01000000011100010000001110110011;
ROM[13723] <= 32'b00000000011100000000001000110011;
ROM[13724] <= 32'b00000000001000000000000110110011;
ROM[13725] <= 32'b01001111010100001001000011101111;
ROM[13726] <= 32'b11111111110000010000000100010011;
ROM[13727] <= 32'b00000000000000010010001110000011;
ROM[13728] <= 32'b00000000011101100010000000100011;
ROM[13729] <= 32'b00000000000000001101001110110111;
ROM[13730] <= 32'b01101101000000111000001110010011;
ROM[13731] <= 32'b00000000111000111000001110110011;
ROM[13732] <= 32'b00000000011100010010000000100011;
ROM[13733] <= 32'b00000000010000010000000100010011;
ROM[13734] <= 32'b00000000001100010010000000100011;
ROM[13735] <= 32'b00000000010000010000000100010011;
ROM[13736] <= 32'b00000000010000010010000000100011;
ROM[13737] <= 32'b00000000010000010000000100010011;
ROM[13738] <= 32'b00000000010100010010000000100011;
ROM[13739] <= 32'b00000000010000010000000100010011;
ROM[13740] <= 32'b00000000011000010010000000100011;
ROM[13741] <= 32'b00000000010000010000000100010011;
ROM[13742] <= 32'b00000001010000000000001110010011;
ROM[13743] <= 32'b00000000000000111000001110010011;
ROM[13744] <= 32'b01000000011100010000001110110011;
ROM[13745] <= 32'b00000000011100000000001000110011;
ROM[13746] <= 32'b00000000001000000000000110110011;
ROM[13747] <= 32'b01001001110100001001000011101111;
ROM[13748] <= 32'b11111111110000010000000100010011;
ROM[13749] <= 32'b00000000000000010010001110000011;
ROM[13750] <= 32'b00000000011101100010000000100011;
ROM[13751] <= 32'b10101000100011111010000011101111;
ROM[13752] <= 32'b00000000100000011010001110000011;
ROM[13753] <= 32'b00000000011100010010000000100011;
ROM[13754] <= 32'b00000000010000010000000100010011;
ROM[13755] <= 32'b00000000000100000000001110010011;
ROM[13756] <= 32'b00000000011100010010000000100011;
ROM[13757] <= 32'b00000000010000010000000100010011;
ROM[13758] <= 32'b11111111110000010000000100010011;
ROM[13759] <= 32'b00000000000000010010001110000011;
ROM[13760] <= 32'b11111111110000010000000100010011;
ROM[13761] <= 32'b00000000000000010010010000000011;
ROM[13762] <= 32'b00000000011101000000001110110011;
ROM[13763] <= 32'b00000000011100010010000000100011;
ROM[13764] <= 32'b00000000010000010000000100010011;
ROM[13765] <= 32'b11111111110000010000000100010011;
ROM[13766] <= 32'b00000000000000010010001110000011;
ROM[13767] <= 32'b00000000011100011010010000100011;
ROM[13768] <= 32'b11101000100111111000000011101111;
ROM[13769] <= 32'b00000000000000000000001110010011;
ROM[13770] <= 32'b00000000011100010010000000100011;
ROM[13771] <= 32'b00000000010000010000000100010011;
ROM[13772] <= 32'b00000001010000000000001110010011;
ROM[13773] <= 32'b01000000011100011000001110110011;
ROM[13774] <= 32'b00000000000000111010000010000011;
ROM[13775] <= 32'b11111111110000010000000100010011;
ROM[13776] <= 32'b00000000000000010010001110000011;
ROM[13777] <= 32'b00000000011100100010000000100011;
ROM[13778] <= 32'b00000000010000100000000100010011;
ROM[13779] <= 32'b00000001010000000000001110010011;
ROM[13780] <= 32'b01000000011100011000001110110011;
ROM[13781] <= 32'b00000000010000111010000110000011;
ROM[13782] <= 32'b00000000100000111010001000000011;
ROM[13783] <= 32'b00000000110000111010001010000011;
ROM[13784] <= 32'b00000001000000111010001100000011;
ROM[13785] <= 32'b00000000000000001000000011100111;
ROM[13786] <= 32'b00000000000000000100001110110111;
ROM[13787] <= 32'b11111111111100111000001110010011;
ROM[13788] <= 32'b00000000011100010010000000100011;
ROM[13789] <= 32'b00000000010000010000000100010011;
ROM[13790] <= 32'b11111111110000010000000100010011;
ROM[13791] <= 32'b00000000000000010010001110000011;
ROM[13792] <= 32'b00000100011101101010000000100011;
ROM[13793] <= 32'b00000100000001101010001110000011;
ROM[13794] <= 32'b00000000011100010010000000100011;
ROM[13795] <= 32'b00000000010000010000000100010011;
ROM[13796] <= 32'b00000100000001101010001110000011;
ROM[13797] <= 32'b00000000011100010010000000100011;
ROM[13798] <= 32'b00000000010000010000000100010011;
ROM[13799] <= 32'b11111111110000010000000100010011;
ROM[13800] <= 32'b00000000000000010010001110000011;
ROM[13801] <= 32'b11111111110000010000000100010011;
ROM[13802] <= 32'b00000000000000010010010000000011;
ROM[13803] <= 32'b00000000011101000000001110110011;
ROM[13804] <= 32'b00000000011100010010000000100011;
ROM[13805] <= 32'b00000000010000010000000100010011;
ROM[13806] <= 32'b00000100000001101010001110000011;
ROM[13807] <= 32'b00000000011100010010000000100011;
ROM[13808] <= 32'b00000000010000010000000100010011;
ROM[13809] <= 32'b11111111110000010000000100010011;
ROM[13810] <= 32'b00000000000000010010001110000011;
ROM[13811] <= 32'b11111111110000010000000100010011;
ROM[13812] <= 32'b00000000000000010010010000000011;
ROM[13813] <= 32'b00000000011101000000001110110011;
ROM[13814] <= 32'b00000000011100010010000000100011;
ROM[13815] <= 32'b00000000010000010000000100010011;
ROM[13816] <= 32'b00000100000001101010001110000011;
ROM[13817] <= 32'b00000000011100010010000000100011;
ROM[13818] <= 32'b00000000010000010000000100010011;
ROM[13819] <= 32'b11111111110000010000000100010011;
ROM[13820] <= 32'b00000000000000010010001110000011;
ROM[13821] <= 32'b11111111110000010000000100010011;
ROM[13822] <= 32'b00000000000000010010010000000011;
ROM[13823] <= 32'b00000000011101000000001110110011;
ROM[13824] <= 32'b00000000011100010010000000100011;
ROM[13825] <= 32'b00000000010000010000000100010011;
ROM[13826] <= 32'b11111111110000010000000100010011;
ROM[13827] <= 32'b00000000000000010010001110000011;
ROM[13828] <= 32'b00000100011101101010000000100011;
ROM[13829] <= 32'b00000000000000000000001110010011;
ROM[13830] <= 32'b00000000011100010010000000100011;
ROM[13831] <= 32'b00000000010000010000000100010011;
ROM[13832] <= 32'b00000001010000000000001110010011;
ROM[13833] <= 32'b01000000011100011000001110110011;
ROM[13834] <= 32'b00000000000000111010000010000011;
ROM[13835] <= 32'b11111111110000010000000100010011;
ROM[13836] <= 32'b00000000000000010010001110000011;
ROM[13837] <= 32'b00000000011100100010000000100011;
ROM[13838] <= 32'b00000000010000100000000100010011;
ROM[13839] <= 32'b00000001010000000000001110010011;
ROM[13840] <= 32'b01000000011100011000001110110011;
ROM[13841] <= 32'b00000000010000111010000110000011;
ROM[13842] <= 32'b00000000100000111010001000000011;
ROM[13843] <= 32'b00000000110000111010001010000011;
ROM[13844] <= 32'b00000001000000111010001100000011;
ROM[13845] <= 32'b00000000000000001000000011100111;
ROM[13846] <= 32'b00000100000001101010001110000011;
ROM[13847] <= 32'b00000000011100010010000000100011;
ROM[13848] <= 32'b00000000010000010000000100010011;
ROM[13849] <= 32'b00000000000000000000001110010011;
ROM[13850] <= 32'b00000000011100010010000000100011;
ROM[13851] <= 32'b00000000010000010000000100010011;
ROM[13852] <= 32'b11111111110000010000000100010011;
ROM[13853] <= 32'b00000000000000010010001110000011;
ROM[13854] <= 32'b11111111110000010000000100010011;
ROM[13855] <= 32'b00000000000000010010010000000011;
ROM[13856] <= 32'b00000000011101000000001110110011;
ROM[13857] <= 32'b00000000011100010010000000100011;
ROM[13858] <= 32'b00000000010000010000000100010011;
ROM[13859] <= 32'b11111111110000010000000100010011;
ROM[13860] <= 32'b00000000000000010010001110000011;
ROM[13861] <= 32'b00000000000000111000001100010011;
ROM[13862] <= 32'b00000000110100110000010000110011;
ROM[13863] <= 32'b00000000000001000010001110000011;
ROM[13864] <= 32'b00000000011100010010000000100011;
ROM[13865] <= 32'b00000000010000010000000100010011;
ROM[13866] <= 32'b00000001010000000000001110010011;
ROM[13867] <= 32'b01000000011100011000001110110011;
ROM[13868] <= 32'b00000000000000111010000010000011;
ROM[13869] <= 32'b11111111110000010000000100010011;
ROM[13870] <= 32'b00000000000000010010001110000011;
ROM[13871] <= 32'b00000000011100100010000000100011;
ROM[13872] <= 32'b00000000010000100000000100010011;
ROM[13873] <= 32'b00000001010000000000001110010011;
ROM[13874] <= 32'b01000000011100011000001110110011;
ROM[13875] <= 32'b00000000010000111010000110000011;
ROM[13876] <= 32'b00000000100000111010001000000011;
ROM[13877] <= 32'b00000000110000111010001010000011;
ROM[13878] <= 32'b00000001000000111010001100000011;
ROM[13879] <= 32'b00000000000000001000000011100111;
ROM[13880] <= 32'b00000000000000010010000000100011;
ROM[13881] <= 32'b00000000010000010000000100010011;
ROM[13882] <= 32'b00000000000000010010000000100011;
ROM[13883] <= 32'b00000000010000010000000100010011;
ROM[13884] <= 32'b00000000000000000000001110010011;
ROM[13885] <= 32'b00000000011100010010000000100011;
ROM[13886] <= 32'b00000000010000010000000100010011;
ROM[13887] <= 32'b11111111110000010000000100010011;
ROM[13888] <= 32'b00000000000000010010001110000011;
ROM[13889] <= 32'b00000000011100011010001000100011;
ROM[13890] <= 32'b00000000010000011010001110000011;
ROM[13891] <= 32'b00000000011100010010000000100011;
ROM[13892] <= 32'b00000000010000010000000100010011;
ROM[13893] <= 32'b00000000000000000000001110010011;
ROM[13894] <= 32'b00000000011100010010000000100011;
ROM[13895] <= 32'b00000000010000010000000100010011;
ROM[13896] <= 32'b11111111110000010000000100010011;
ROM[13897] <= 32'b00000000000000010010001110000011;
ROM[13898] <= 32'b11111111110000010000000100010011;
ROM[13899] <= 32'b00000000000000010010010000000011;
ROM[13900] <= 32'b00000000011101000010010010110011;
ROM[13901] <= 32'b00000000100000111010010100110011;
ROM[13902] <= 32'b00000000101001001000001110110011;
ROM[13903] <= 32'b00000000000100111000001110010011;
ROM[13904] <= 32'b00000000000100111111001110010011;
ROM[13905] <= 32'b00000000011100010010000000100011;
ROM[13906] <= 32'b00000000010000010000000100010011;
ROM[13907] <= 32'b11111111110000010000000100010011;
ROM[13908] <= 32'b00000000000000010010001110000011;
ROM[13909] <= 32'b01000000011100000000001110110011;
ROM[13910] <= 32'b00000000000100111000001110010011;
ROM[13911] <= 32'b00000000011100010010000000100011;
ROM[13912] <= 32'b00000000010000010000000100010011;
ROM[13913] <= 32'b11111111110000010000000100010011;
ROM[13914] <= 32'b00000000000000010010001110000011;
ROM[13915] <= 32'b00000000000000111000101001100011;
ROM[13916] <= 32'b00000000000000001110001110110111;
ROM[13917] <= 32'b10100101100000111000001110010011;
ROM[13918] <= 32'b00000000111000111000001110110011;
ROM[13919] <= 32'b00000000000000111000000011100111;
ROM[13920] <= 32'b00000000000000001110001110110111;
ROM[13921] <= 32'b10011100110000111000001110010011;
ROM[13922] <= 32'b00000000111000111000001110110011;
ROM[13923] <= 32'b00000000011100010010000000100011;
ROM[13924] <= 32'b00000000010000010000000100010011;
ROM[13925] <= 32'b00000000001100010010000000100011;
ROM[13926] <= 32'b00000000010000010000000100010011;
ROM[13927] <= 32'b00000000010000010010000000100011;
ROM[13928] <= 32'b00000000010000010000000100010011;
ROM[13929] <= 32'b00000000010100010010000000100011;
ROM[13930] <= 32'b00000000010000010000000100010011;
ROM[13931] <= 32'b00000000011000010010000000100011;
ROM[13932] <= 32'b00000000010000010000000100010011;
ROM[13933] <= 32'b00000001010000000000001110010011;
ROM[13934] <= 32'b00000000000000111000001110010011;
ROM[13935] <= 32'b01000000011100010000001110110011;
ROM[13936] <= 32'b00000000011100000000001000110011;
ROM[13937] <= 32'b00000000001000000000000110110011;
ROM[13938] <= 32'b11101001000111111111000011101111;
ROM[13939] <= 32'b11111111110000010000000100010011;
ROM[13940] <= 32'b00000000000000010010001110000011;
ROM[13941] <= 32'b00000000011100011010000000100011;
ROM[13942] <= 32'b00000000000000011010001110000011;
ROM[13943] <= 32'b00000000011100010010000000100011;
ROM[13944] <= 32'b00000000010000010000000100010011;
ROM[13945] <= 32'b00000000000000000000001110010011;
ROM[13946] <= 32'b00000000011100010010000000100011;
ROM[13947] <= 32'b00000000010000010000000100010011;
ROM[13948] <= 32'b11111111110000010000000100010011;
ROM[13949] <= 32'b00000000000000010010001110000011;
ROM[13950] <= 32'b11111111110000010000000100010011;
ROM[13951] <= 32'b00000000000000010010010000000011;
ROM[13952] <= 32'b00000000011101000010010010110011;
ROM[13953] <= 32'b00000000100000111010010100110011;
ROM[13954] <= 32'b00000000101001001000001110110011;
ROM[13955] <= 32'b00000000000100111000001110010011;
ROM[13956] <= 32'b00000000000100111111001110010011;
ROM[13957] <= 32'b00000000011100010010000000100011;
ROM[13958] <= 32'b00000000010000010000000100010011;
ROM[13959] <= 32'b11111111110000010000000100010011;
ROM[13960] <= 32'b00000000000000010010001110000011;
ROM[13961] <= 32'b00000000000000111000101001100011;
ROM[13962] <= 32'b00000000000000001110001110110111;
ROM[13963] <= 32'b10100101010000111000001110010011;
ROM[13964] <= 32'b00000000111000111000001110110011;
ROM[13965] <= 32'b00000000000000111000000011100111;
ROM[13966] <= 32'b00000000000100000000001110010011;
ROM[13967] <= 32'b00000000011100010010000000100011;
ROM[13968] <= 32'b00000000010000010000000100010011;
ROM[13969] <= 32'b11111111110000010000000100010011;
ROM[13970] <= 32'b00000000000000010010001110000011;
ROM[13971] <= 32'b00000000011100011010001000100011;
ROM[13972] <= 32'b00000000010000000000000011101111;
ROM[13973] <= 32'b11101011010111111111000011101111;
ROM[13974] <= 32'b00000000000000011010001110000011;
ROM[13975] <= 32'b00000000011100010010000000100011;
ROM[13976] <= 32'b00000000010000010000000100010011;
ROM[13977] <= 32'b00000110000000000000001110010011;
ROM[13978] <= 32'b00000000011100010010000000100011;
ROM[13979] <= 32'b00000000010000010000000100010011;
ROM[13980] <= 32'b11111111110000010000000100010011;
ROM[13981] <= 32'b00000000000000010010001110000011;
ROM[13982] <= 32'b11111111110000010000000100010011;
ROM[13983] <= 32'b00000000000000010010010000000011;
ROM[13984] <= 32'b00000000100000111010001110110011;
ROM[13985] <= 32'b00000000011100010010000000100011;
ROM[13986] <= 32'b00000000010000010000000100010011;
ROM[13987] <= 32'b11111111110000010000000100010011;
ROM[13988] <= 32'b00000000000000010010001110000011;
ROM[13989] <= 32'b00000000000000111000101001100011;
ROM[13990] <= 32'b00000000000000001110001110110111;
ROM[13991] <= 32'b10101010110000111000001110010011;
ROM[13992] <= 32'b00000000111000111000001110110011;
ROM[13993] <= 32'b00000000000000111000000011100111;
ROM[13994] <= 32'b00001001100000000000000011101111;
ROM[13995] <= 32'b00000000000000011010001110000011;
ROM[13996] <= 32'b00000000011100010010000000100011;
ROM[13997] <= 32'b00000000010000010000000100010011;
ROM[13998] <= 32'b00000111101100000000001110010011;
ROM[13999] <= 32'b00000000011100010010000000100011;
ROM[14000] <= 32'b00000000010000010000000100010011;
ROM[14001] <= 32'b11111111110000010000000100010011;
ROM[14002] <= 32'b00000000000000010010001110000011;
ROM[14003] <= 32'b11111111110000010000000100010011;
ROM[14004] <= 32'b00000000000000010010010000000011;
ROM[14005] <= 32'b00000000011101000010001110110011;
ROM[14006] <= 32'b00000000011100010010000000100011;
ROM[14007] <= 32'b00000000010000010000000100010011;
ROM[14008] <= 32'b11111111110000010000000100010011;
ROM[14009] <= 32'b00000000000000010010001110000011;
ROM[14010] <= 32'b00000000000000111000101001100011;
ROM[14011] <= 32'b00000000000000001110001110110111;
ROM[14012] <= 32'b10110000000000111000001110010011;
ROM[14013] <= 32'b00000000111000111000001110110011;
ROM[14014] <= 32'b00000000000000111000000011100111;
ROM[14015] <= 32'b00000100010000000000000011101111;
ROM[14016] <= 32'b00000000000000011010001110000011;
ROM[14017] <= 32'b00000000011100010010000000100011;
ROM[14018] <= 32'b00000000010000010000000100010011;
ROM[14019] <= 32'b00000010000000000000001110010011;
ROM[14020] <= 32'b00000000011100010010000000100011;
ROM[14021] <= 32'b00000000010000010000000100010011;
ROM[14022] <= 32'b11111111110000010000000100010011;
ROM[14023] <= 32'b00000000000000010010001110000011;
ROM[14024] <= 32'b11111111110000010000000100010011;
ROM[14025] <= 32'b00000000000000010010010000000011;
ROM[14026] <= 32'b01000000011101000000001110110011;
ROM[14027] <= 32'b00000000011100010010000000100011;
ROM[14028] <= 32'b00000000010000010000000100010011;
ROM[14029] <= 32'b11111111110000010000000100010011;
ROM[14030] <= 32'b00000000000000010010001110000011;
ROM[14031] <= 32'b00000000011100011010000000100011;
ROM[14032] <= 32'b00000000000000011010001110000011;
ROM[14033] <= 32'b00000000011100010010000000100011;
ROM[14034] <= 32'b00000000010000010000000100010011;
ROM[14035] <= 32'b00000000000000001110001110110111;
ROM[14036] <= 32'b10111001100000111000001110010011;
ROM[14037] <= 32'b00000000111000111000001110110011;
ROM[14038] <= 32'b00000000011100010010000000100011;
ROM[14039] <= 32'b00000000010000010000000100010011;
ROM[14040] <= 32'b00000000001100010010000000100011;
ROM[14041] <= 32'b00000000010000010000000100010011;
ROM[14042] <= 32'b00000000010000010010000000100011;
ROM[14043] <= 32'b00000000010000010000000100010011;
ROM[14044] <= 32'b00000000010100010010000000100011;
ROM[14045] <= 32'b00000000010000010000000100010011;
ROM[14046] <= 32'b00000000011000010010000000100011;
ROM[14047] <= 32'b00000000010000010000000100010011;
ROM[14048] <= 32'b00000001010000000000001110010011;
ROM[14049] <= 32'b00000000010000111000001110010011;
ROM[14050] <= 32'b01000000011100010000001110110011;
ROM[14051] <= 32'b00000000011100000000001000110011;
ROM[14052] <= 32'b00000000001000000000000110110011;
ROM[14053] <= 32'b00001110000000001000000011101111;
ROM[14054] <= 32'b11111111110000010000000100010011;
ROM[14055] <= 32'b00000000000000010010001110000011;
ROM[14056] <= 32'b00000000011101100010000000100011;
ROM[14057] <= 32'b00000000000000011010001110000011;
ROM[14058] <= 32'b00000000011100010010000000100011;
ROM[14059] <= 32'b00000000010000010000000100010011;
ROM[14060] <= 32'b00000001010000000000001110010011;
ROM[14061] <= 32'b01000000011100011000001110110011;
ROM[14062] <= 32'b00000000000000111010000010000011;
ROM[14063] <= 32'b11111111110000010000000100010011;
ROM[14064] <= 32'b00000000000000010010001110000011;
ROM[14065] <= 32'b00000000011100100010000000100011;
ROM[14066] <= 32'b00000000010000100000000100010011;
ROM[14067] <= 32'b00000001010000000000001110010011;
ROM[14068] <= 32'b01000000011100011000001110110011;
ROM[14069] <= 32'b00000000010000111010000110000011;
ROM[14070] <= 32'b00000000100000111010001000000011;
ROM[14071] <= 32'b00000000110000111010001010000011;
ROM[14072] <= 32'b00000001000000111010001100000011;
ROM[14073] <= 32'b00000000000000001000000011100111;
ROM[14074] <= 32'b00000000000000010010000000100011;
ROM[14075] <= 32'b00000000010000010000000100010011;
ROM[14076] <= 32'b00000000000000010010000000100011;
ROM[14077] <= 32'b00000000010000010000000100010011;
ROM[14078] <= 32'b00000100001000000000001110010011;
ROM[14079] <= 32'b00000000011100010010000000100011;
ROM[14080] <= 32'b00000000010000010000000100010011;
ROM[14081] <= 32'b00000000000000001110001110110111;
ROM[14082] <= 32'b11000101000000111000001110010011;
ROM[14083] <= 32'b00000000111000111000001110110011;
ROM[14084] <= 32'b00000000011100010010000000100011;
ROM[14085] <= 32'b00000000010000010000000100010011;
ROM[14086] <= 32'b00000000001100010010000000100011;
ROM[14087] <= 32'b00000000010000010000000100010011;
ROM[14088] <= 32'b00000000010000010010000000100011;
ROM[14089] <= 32'b00000000010000010000000100010011;
ROM[14090] <= 32'b00000000010100010010000000100011;
ROM[14091] <= 32'b00000000010000010000000100010011;
ROM[14092] <= 32'b00000000011000010010000000100011;
ROM[14093] <= 32'b00000000010000010000000100010011;
ROM[14094] <= 32'b00000001010000000000001110010011;
ROM[14095] <= 32'b00000000010000111000001110010011;
ROM[14096] <= 32'b01000000011100010000001110110011;
ROM[14097] <= 32'b00000000011100000000001000110011;
ROM[14098] <= 32'b00000000001000000000000110110011;
ROM[14099] <= 32'b00000010100000001000000011101111;
ROM[14100] <= 32'b11111111110000010000000100010011;
ROM[14101] <= 32'b00000000000000010010001110000011;
ROM[14102] <= 32'b00000000011101100010000000100011;
ROM[14103] <= 32'b00000000000000100010001110000011;
ROM[14104] <= 32'b00000000011100010010000000100011;
ROM[14105] <= 32'b00000000010000010000000100010011;
ROM[14106] <= 32'b00000000000000001110001110110111;
ROM[14107] <= 32'b11001011010000111000001110010011;
ROM[14108] <= 32'b00000000111000111000001110110011;
ROM[14109] <= 32'b00000000011100010010000000100011;
ROM[14110] <= 32'b00000000010000010000000100010011;
ROM[14111] <= 32'b00000000001100010010000000100011;
ROM[14112] <= 32'b00000000010000010000000100010011;
ROM[14113] <= 32'b00000000010000010010000000100011;
ROM[14114] <= 32'b00000000010000010000000100010011;
ROM[14115] <= 32'b00000000010100010010000000100011;
ROM[14116] <= 32'b00000000010000010000000100010011;
ROM[14117] <= 32'b00000000011000010010000000100011;
ROM[14118] <= 32'b00000000010000010000000100010011;
ROM[14119] <= 32'b00000001010000000000001110010011;
ROM[14120] <= 32'b00000000010000111000001110010011;
ROM[14121] <= 32'b01000000011100010000001110110011;
ROM[14122] <= 32'b00000000011100000000001000110011;
ROM[14123] <= 32'b00000000001000000000000110110011;
ROM[14124] <= 32'b00101011100000001001000011101111;
ROM[14125] <= 32'b11111111110000010000000100010011;
ROM[14126] <= 32'b00000000000000010010001110000011;
ROM[14127] <= 32'b00000000011101100010000000100011;
ROM[14128] <= 32'b00000011001000000000001110010011;
ROM[14129] <= 32'b00000000011100010010000000100011;
ROM[14130] <= 32'b00000000010000010000000100010011;
ROM[14131] <= 32'b00000000000000001110001110110111;
ROM[14132] <= 32'b11010001100000111000001110010011;
ROM[14133] <= 32'b00000000111000111000001110110011;
ROM[14134] <= 32'b00000000011100010010000000100011;
ROM[14135] <= 32'b00000000010000010000000100010011;
ROM[14136] <= 32'b00000000001100010010000000100011;
ROM[14137] <= 32'b00000000010000010000000100010011;
ROM[14138] <= 32'b00000000010000010010000000100011;
ROM[14139] <= 32'b00000000010000010000000100010011;
ROM[14140] <= 32'b00000000010100010010000000100011;
ROM[14141] <= 32'b00000000010000010000000100010011;
ROM[14142] <= 32'b00000000011000010010000000100011;
ROM[14143] <= 32'b00000000010000010000000100010011;
ROM[14144] <= 32'b00000001010000000000001110010011;
ROM[14145] <= 32'b00000000010000111000001110010011;
ROM[14146] <= 32'b01000000011100010000001110110011;
ROM[14147] <= 32'b00000000011100000000001000110011;
ROM[14148] <= 32'b00000000001000000000000110110011;
ROM[14149] <= 32'b00100010100100011011000011101111;
ROM[14150] <= 32'b11111111110000010000000100010011;
ROM[14151] <= 32'b00000000000000010010001110000011;
ROM[14152] <= 32'b00000000011100011010000000100011;
ROM[14153] <= 32'b00000000000000001110001110110111;
ROM[14154] <= 32'b11010111000000111000001110010011;
ROM[14155] <= 32'b00000000111000111000001110110011;
ROM[14156] <= 32'b00000000011100010010000000100011;
ROM[14157] <= 32'b00000000010000010000000100010011;
ROM[14158] <= 32'b00000000001100010010000000100011;
ROM[14159] <= 32'b00000000010000010000000100010011;
ROM[14160] <= 32'b00000000010000010010000000100011;
ROM[14161] <= 32'b00000000010000010000000100010011;
ROM[14162] <= 32'b00000000010100010010000000100011;
ROM[14163] <= 32'b00000000010000010000000100010011;
ROM[14164] <= 32'b00000000011000010010000000100011;
ROM[14165] <= 32'b00000000010000010000000100010011;
ROM[14166] <= 32'b00000001010000000000001110010011;
ROM[14167] <= 32'b00000000000000111000001110010011;
ROM[14168] <= 32'b01000000011100010000001110110011;
ROM[14169] <= 32'b00000000011100000000001000110011;
ROM[14170] <= 32'b00000000001000000000000110110011;
ROM[14171] <= 32'b10110111010111111111000011101111;
ROM[14172] <= 32'b11111111110000010000000100010011;
ROM[14173] <= 32'b00000000000000010010001110000011;
ROM[14174] <= 32'b00000000011100011010001000100011;
ROM[14175] <= 32'b00000000010000011010001110000011;
ROM[14176] <= 32'b00000000011100010010000000100011;
ROM[14177] <= 32'b00000000010000010000000100010011;
ROM[14178] <= 32'b00000000000000001110001110110111;
ROM[14179] <= 32'b11011101010000111000001110010011;
ROM[14180] <= 32'b00000000111000111000001110110011;
ROM[14181] <= 32'b00000000011100010010000000100011;
ROM[14182] <= 32'b00000000010000010000000100010011;
ROM[14183] <= 32'b00000000001100010010000000100011;
ROM[14184] <= 32'b00000000010000010000000100010011;
ROM[14185] <= 32'b00000000010000010010000000100011;
ROM[14186] <= 32'b00000000010000010000000100010011;
ROM[14187] <= 32'b00000000010100010010000000100011;
ROM[14188] <= 32'b00000000010000010000000100010011;
ROM[14189] <= 32'b00000000011000010010000000100011;
ROM[14190] <= 32'b00000000010000010000000100010011;
ROM[14191] <= 32'b00000001010000000000001110010011;
ROM[14192] <= 32'b00000000000000111000001110010011;
ROM[14193] <= 32'b01000000011100010000001110110011;
ROM[14194] <= 32'b00000000011100000000001000110011;
ROM[14195] <= 32'b00000000001000000000000110110011;
ROM[14196] <= 32'b01100111010100011100000011101111;
ROM[14197] <= 32'b11111111110000010000000100010011;
ROM[14198] <= 32'b00000000000000010010001110000011;
ROM[14199] <= 32'b11111111110000010000000100010011;
ROM[14200] <= 32'b00000000000000010010010000000011;
ROM[14201] <= 32'b00000000011101000010010010110011;
ROM[14202] <= 32'b00000000100000111010010100110011;
ROM[14203] <= 32'b00000000101001001000001110110011;
ROM[14204] <= 32'b00000000000100111000001110010011;
ROM[14205] <= 32'b00000000000100111111001110010011;
ROM[14206] <= 32'b00000000011100010010000000100011;
ROM[14207] <= 32'b00000000010000010000000100010011;
ROM[14208] <= 32'b11111111110000010000000100010011;
ROM[14209] <= 32'b00000000000000010010001110000011;
ROM[14210] <= 32'b01000000011100000000001110110011;
ROM[14211] <= 32'b00000000000100111000001110010011;
ROM[14212] <= 32'b00000000011100010010000000100011;
ROM[14213] <= 32'b00000000010000010000000100010011;
ROM[14214] <= 32'b11111111110000010000000100010011;
ROM[14215] <= 32'b00000000000000010010001110000011;
ROM[14216] <= 32'b01000000011100000000001110110011;
ROM[14217] <= 32'b00000000000100111000001110010011;
ROM[14218] <= 32'b00000000011100010010000000100011;
ROM[14219] <= 32'b00000000010000010000000100010011;
ROM[14220] <= 32'b11111111110000010000000100010011;
ROM[14221] <= 32'b00000000000000010010001110000011;
ROM[14222] <= 32'b00000000000000111000101001100011;
ROM[14223] <= 32'b00000000000000001110001110110111;
ROM[14224] <= 32'b00000010000000111000001110010011;
ROM[14225] <= 32'b00000000111000111000001110110011;
ROM[14226] <= 32'b00000000000000111000000011100111;
ROM[14227] <= 32'b00000000010000011010001110000011;
ROM[14228] <= 32'b00000000011100010010000000100011;
ROM[14229] <= 32'b00000000010000010000000100010011;
ROM[14230] <= 32'b00000000000000001110001110110111;
ROM[14231] <= 32'b11101010010000111000001110010011;
ROM[14232] <= 32'b00000000111000111000001110110011;
ROM[14233] <= 32'b00000000011100010010000000100011;
ROM[14234] <= 32'b00000000010000010000000100010011;
ROM[14235] <= 32'b00000000001100010010000000100011;
ROM[14236] <= 32'b00000000010000010000000100010011;
ROM[14237] <= 32'b00000000010000010010000000100011;
ROM[14238] <= 32'b00000000010000010000000100010011;
ROM[14239] <= 32'b00000000010100010010000000100011;
ROM[14240] <= 32'b00000000010000010000000100010011;
ROM[14241] <= 32'b00000000011000010010000000100011;
ROM[14242] <= 32'b00000000010000010000000100010011;
ROM[14243] <= 32'b00000001010000000000001110010011;
ROM[14244] <= 32'b00000000000000111000001110010011;
ROM[14245] <= 32'b01000000011100010000001110110011;
ROM[14246] <= 32'b00000000011100000000001000110011;
ROM[14247] <= 32'b00000000001000000000000110110011;
ROM[14248] <= 32'b01011110100100011100000011101111;
ROM[14249] <= 32'b11111111110000010000000100010011;
ROM[14250] <= 32'b00000000000000010010001110000011;
ROM[14251] <= 32'b11111111110000010000000100010011;
ROM[14252] <= 32'b00000000000000010010010000000011;
ROM[14253] <= 32'b00000000011101000010010010110011;
ROM[14254] <= 32'b00000000100000111010010100110011;
ROM[14255] <= 32'b00000000101001001000001110110011;
ROM[14256] <= 32'b00000000000100111000001110010011;
ROM[14257] <= 32'b00000000000100111111001110010011;
ROM[14258] <= 32'b00000000011100010010000000100011;
ROM[14259] <= 32'b00000000010000010000000100010011;
ROM[14260] <= 32'b11111111110000010000000100010011;
ROM[14261] <= 32'b00000000000000010010001110000011;
ROM[14262] <= 32'b00000000000000111000101001100011;
ROM[14263] <= 32'b00000000000000001110001110110111;
ROM[14264] <= 32'b11110110000000111000001110010011;
ROM[14265] <= 32'b00000000111000111000001110110011;
ROM[14266] <= 32'b00000000000000111000000011100111;
ROM[14267] <= 32'b00000000000000011010001110000011;
ROM[14268] <= 32'b00000000011100010010000000100011;
ROM[14269] <= 32'b00000000010000010000000100010011;
ROM[14270] <= 32'b00000000010000011010001110000011;
ROM[14271] <= 32'b00000000011100010010000000100011;
ROM[14272] <= 32'b00000000010000010000000100010011;
ROM[14273] <= 32'b00000000000000001110001110110111;
ROM[14274] <= 32'b11110101000000111000001110010011;
ROM[14275] <= 32'b00000000111000111000001110110011;
ROM[14276] <= 32'b00000000011100010010000000100011;
ROM[14277] <= 32'b00000000010000010000000100010011;
ROM[14278] <= 32'b00000000001100010010000000100011;
ROM[14279] <= 32'b00000000010000010000000100010011;
ROM[14280] <= 32'b00000000010000010010000000100011;
ROM[14281] <= 32'b00000000010000010000000100010011;
ROM[14282] <= 32'b00000000010100010010000000100011;
ROM[14283] <= 32'b00000000010000010000000100010011;
ROM[14284] <= 32'b00000000011000010010000000100011;
ROM[14285] <= 32'b00000000010000010000000100010011;
ROM[14286] <= 32'b00000001010000000000001110010011;
ROM[14287] <= 32'b00000000100000111000001110010011;
ROM[14288] <= 32'b01000000011100010000001110110011;
ROM[14289] <= 32'b00000000011100000000001000110011;
ROM[14290] <= 32'b00000000001000000000000110110011;
ROM[14291] <= 32'b01000110000100011011000011101111;
ROM[14292] <= 32'b11111111110000010000000100010011;
ROM[14293] <= 32'b00000000000000010010001110000011;
ROM[14294] <= 32'b00000000011101100010000000100011;
ROM[14295] <= 32'b00000110100000000000000011101111;
ROM[14296] <= 32'b00000000000000011010001110000011;
ROM[14297] <= 32'b00000000011100010010000000100011;
ROM[14298] <= 32'b00000000010000010000000100010011;
ROM[14299] <= 32'b00000000000000001110001110110111;
ROM[14300] <= 32'b11111011100000111000001110010011;
ROM[14301] <= 32'b00000000111000111000001110110011;
ROM[14302] <= 32'b00000000011100010010000000100011;
ROM[14303] <= 32'b00000000010000010000000100010011;
ROM[14304] <= 32'b00000000001100010010000000100011;
ROM[14305] <= 32'b00000000010000010000000100010011;
ROM[14306] <= 32'b00000000010000010010000000100011;
ROM[14307] <= 32'b00000000010000010000000100010011;
ROM[14308] <= 32'b00000000010100010010000000100011;
ROM[14309] <= 32'b00000000010000010000000100010011;
ROM[14310] <= 32'b00000000011000010010000000100011;
ROM[14311] <= 32'b00000000010000010000000100010011;
ROM[14312] <= 32'b00000001010000000000001110010011;
ROM[14313] <= 32'b00000000010000111000001110010011;
ROM[14314] <= 32'b01000000011100010000001110110011;
ROM[14315] <= 32'b00000000011100000000001000110011;
ROM[14316] <= 32'b00000000001000000000000110110011;
ROM[14317] <= 32'b01011101100100011011000011101111;
ROM[14318] <= 32'b11111111110000010000000100010011;
ROM[14319] <= 32'b00000000000000010010001110000011;
ROM[14320] <= 32'b00000000011101100010000000100011;
ROM[14321] <= 32'b00000000000000001110001110110111;
ROM[14322] <= 32'b00000001000000111000001110010011;
ROM[14323] <= 32'b00000000111000111000001110110011;
ROM[14324] <= 32'b00000000011100010010000000100011;
ROM[14325] <= 32'b00000000010000010000000100010011;
ROM[14326] <= 32'b00000000001100010010000000100011;
ROM[14327] <= 32'b00000000010000010000000100010011;
ROM[14328] <= 32'b00000000010000010010000000100011;
ROM[14329] <= 32'b00000000010000010000000100010011;
ROM[14330] <= 32'b00000000010100010010000000100011;
ROM[14331] <= 32'b00000000010000010000000100010011;
ROM[14332] <= 32'b00000000011000010010000000100011;
ROM[14333] <= 32'b00000000010000010000000100010011;
ROM[14334] <= 32'b00000001010000000000001110010011;
ROM[14335] <= 32'b00000000000000111000001110010011;
ROM[14336] <= 32'b01000000011100010000001110110011;
ROM[14337] <= 32'b00000000011100000000001000110011;
ROM[14338] <= 32'b00000000001000000000000110110011;
ROM[14339] <= 32'b10001101010111111111000011101111;
ROM[14340] <= 32'b11111111110000010000000100010011;
ROM[14341] <= 32'b00000000000000010010001110000011;
ROM[14342] <= 32'b00000000011100011010001000100011;
ROM[14343] <= 32'b11010110000111111111000011101111;
ROM[14344] <= 32'b00000100001100000000001110010011;
ROM[14345] <= 32'b00000000011100010010000000100011;
ROM[14346] <= 32'b00000000010000010000000100010011;
ROM[14347] <= 32'b00000000000000001110001110110111;
ROM[14348] <= 32'b00000111100000111000001110010011;
ROM[14349] <= 32'b00000000111000111000001110110011;
ROM[14350] <= 32'b00000000011100010010000000100011;
ROM[14351] <= 32'b00000000010000010000000100010011;
ROM[14352] <= 32'b00000000001100010010000000100011;
ROM[14353] <= 32'b00000000010000010000000100010011;
ROM[14354] <= 32'b00000000010000010010000000100011;
ROM[14355] <= 32'b00000000010000010000000100010011;
ROM[14356] <= 32'b00000000010100010010000000100011;
ROM[14357] <= 32'b00000000010000010000000100010011;
ROM[14358] <= 32'b00000000011000010010000000100011;
ROM[14359] <= 32'b00000000010000010000000100010011;
ROM[14360] <= 32'b00000001010000000000001110010011;
ROM[14361] <= 32'b00000000010000111000001110010011;
ROM[14362] <= 32'b01000000011100010000001110110011;
ROM[14363] <= 32'b00000000011100000000001000110011;
ROM[14364] <= 32'b00000000001000000000000110110011;
ROM[14365] <= 32'b01000000000100000111000011101111;
ROM[14366] <= 32'b11111111110000010000000100010011;
ROM[14367] <= 32'b00000000000000010010001110000011;
ROM[14368] <= 32'b00000000011101100010000000100011;
ROM[14369] <= 32'b00000000000000011010001110000011;
ROM[14370] <= 32'b00000000011100010010000000100011;
ROM[14371] <= 32'b00000000010000010000000100010011;
ROM[14372] <= 32'b00000001010000000000001110010011;
ROM[14373] <= 32'b01000000011100011000001110110011;
ROM[14374] <= 32'b00000000000000111010000010000011;
ROM[14375] <= 32'b11111111110000010000000100010011;
ROM[14376] <= 32'b00000000000000010010001110000011;
ROM[14377] <= 32'b00000000011100100010000000100011;
ROM[14378] <= 32'b00000000010000100000000100010011;
ROM[14379] <= 32'b00000001010000000000001110010011;
ROM[14380] <= 32'b01000000011100011000001110110011;
ROM[14381] <= 32'b00000000010000111010000110000011;
ROM[14382] <= 32'b00000000100000111010001000000011;
ROM[14383] <= 32'b00000000110000111010001010000011;
ROM[14384] <= 32'b00000001000000111010001100000011;
ROM[14385] <= 32'b00000000000000001000000011100111;
ROM[14386] <= 32'b00000000000000010010000000100011;
ROM[14387] <= 32'b00000000010000010000000100010011;
ROM[14388] <= 32'b00000000000000100010001110000011;
ROM[14389] <= 32'b00000000011100010010000000100011;
ROM[14390] <= 32'b00000000010000010000000100010011;
ROM[14391] <= 32'b00000000000000001110001110110111;
ROM[14392] <= 32'b00010010100000111000001110010011;
ROM[14393] <= 32'b00000000111000111000001110110011;
ROM[14394] <= 32'b00000000011100010010000000100011;
ROM[14395] <= 32'b00000000010000010000000100010011;
ROM[14396] <= 32'b00000000001100010010000000100011;
ROM[14397] <= 32'b00000000010000010000000100010011;
ROM[14398] <= 32'b00000000010000010010000000100011;
ROM[14399] <= 32'b00000000010000010000000100010011;
ROM[14400] <= 32'b00000000010100010010000000100011;
ROM[14401] <= 32'b00000000010000010000000100010011;
ROM[14402] <= 32'b00000000011000010010000000100011;
ROM[14403] <= 32'b00000000010000010000000100010011;
ROM[14404] <= 32'b00000001010000000000001110010011;
ROM[14405] <= 32'b00000000010000111000001110010011;
ROM[14406] <= 32'b01000000011100010000001110110011;
ROM[14407] <= 32'b00000000011100000000001000110011;
ROM[14408] <= 32'b00000000001000000000000110110011;
ROM[14409] <= 32'b10101100010111111111000011101111;
ROM[14410] <= 32'b11111111110000010000000100010011;
ROM[14411] <= 32'b00000000000000010010001110000011;
ROM[14412] <= 32'b00000000011100011010000000100011;
ROM[14413] <= 32'b00000000000000011010001110000011;
ROM[14414] <= 32'b00000000011100010010000000100011;
ROM[14415] <= 32'b00000000010000010000000100010011;
ROM[14416] <= 32'b00000000000000001110001110110111;
ROM[14417] <= 32'b00011000110000111000001110010011;
ROM[14418] <= 32'b00000000111000111000001110110011;
ROM[14419] <= 32'b00000000011100010010000000100011;
ROM[14420] <= 32'b00000000010000010000000100010011;
ROM[14421] <= 32'b00000000001100010010000000100011;
ROM[14422] <= 32'b00000000010000010000000100010011;
ROM[14423] <= 32'b00000000010000010010000000100011;
ROM[14424] <= 32'b00000000010000010000000100010011;
ROM[14425] <= 32'b00000000010100010010000000100011;
ROM[14426] <= 32'b00000000010000010000000100010011;
ROM[14427] <= 32'b00000000011000010010000000100011;
ROM[14428] <= 32'b00000000010000010000000100010011;
ROM[14429] <= 32'b00000001010000000000001110010011;
ROM[14430] <= 32'b00000000010000111000001110010011;
ROM[14431] <= 32'b01000000011100010000001110110011;
ROM[14432] <= 32'b00000000011100000000001000110011;
ROM[14433] <= 32'b00000000001000000000000110110011;
ROM[14434] <= 32'b01010000000100011011000011101111;
ROM[14435] <= 32'b00000001010000000000001110010011;
ROM[14436] <= 32'b01000000011100011000001110110011;
ROM[14437] <= 32'b00000000000000111010000010000011;
ROM[14438] <= 32'b11111111110000010000000100010011;
ROM[14439] <= 32'b00000000000000010010001110000011;
ROM[14440] <= 32'b00000000011100100010000000100011;
ROM[14441] <= 32'b00000000010000100000000100010011;
ROM[14442] <= 32'b00000001010000000000001110010011;
ROM[14443] <= 32'b01000000011100011000001110110011;
ROM[14444] <= 32'b00000000010000111010000110000011;
ROM[14445] <= 32'b00000000100000111010001000000011;
ROM[14446] <= 32'b00000000110000111010001010000011;
ROM[14447] <= 32'b00000001000000111010001100000011;
ROM[14448] <= 32'b00000000000000001000000011100111;
ROM[14449] <= 32'b00000000000000010010000000100011;
ROM[14450] <= 32'b00000000010000010000000100010011;
ROM[14451] <= 32'b00000000000000010010000000100011;
ROM[14452] <= 32'b00000000010000010000000100010011;
ROM[14453] <= 32'b00000000000000010010000000100011;
ROM[14454] <= 32'b00000000010000010000000100010011;
ROM[14455] <= 32'b00000000000000010010000000100011;
ROM[14456] <= 32'b00000000010000010000000100010011;
ROM[14457] <= 32'b00000000000000010010000000100011;
ROM[14458] <= 32'b00000000010000010000000100010011;
ROM[14459] <= 32'b00000000000000010010000000100011;
ROM[14460] <= 32'b00000000010000010000000100010011;
ROM[14461] <= 32'b00000000000000010010000000100011;
ROM[14462] <= 32'b00000000010000010000000100010011;
ROM[14463] <= 32'b00000000000000010010000000100011;
ROM[14464] <= 32'b00000000010000010000000100010011;
ROM[14465] <= 32'b00000000000000010010000000100011;
ROM[14466] <= 32'b00000000010000010000000100010011;
ROM[14467] <= 32'b00000000000000010010000000100011;
ROM[14468] <= 32'b00000000010000010000000100010011;
ROM[14469] <= 32'b00000000000000010010000000100011;
ROM[14470] <= 32'b00000000010000010000000100010011;
ROM[14471] <= 32'b00000000000000010010000000100011;
ROM[14472] <= 32'b00000000010000010000000100010011;
ROM[14473] <= 32'b00000000000000010010000000100011;
ROM[14474] <= 32'b00000000010000010000000100010011;
ROM[14475] <= 32'b00000000000000010010000000100011;
ROM[14476] <= 32'b00000000010000010000000100010011;
ROM[14477] <= 32'b00000100001100000000001110010011;
ROM[14478] <= 32'b00000000011100010010000000100011;
ROM[14479] <= 32'b00000000010000010000000100010011;
ROM[14480] <= 32'b11111111110000010000000100010011;
ROM[14481] <= 32'b00000000000000010010001110000011;
ROM[14482] <= 32'b00000010011100011010000000100011;
ROM[14483] <= 32'b00000100110000000000001110010011;
ROM[14484] <= 32'b00000000011100010010000000100011;
ROM[14485] <= 32'b00000000010000010000000100010011;
ROM[14486] <= 32'b11111111110000010000000100010011;
ROM[14487] <= 32'b00000000000000010010001110000011;
ROM[14488] <= 32'b00000000011100011010111000100011;
ROM[14489] <= 32'b00000100011000000000001110010011;
ROM[14490] <= 32'b00000000011100010010000000100011;
ROM[14491] <= 32'b00000000010000010000000100010011;
ROM[14492] <= 32'b11111111110000010000000100010011;
ROM[14493] <= 32'b00000000000000010010001110000011;
ROM[14494] <= 32'b00000010011100011010010000100011;
ROM[14495] <= 32'b00000101000100000000001110010011;
ROM[14496] <= 32'b00000000011100010010000000100011;
ROM[14497] <= 32'b00000000010000010000000100010011;
ROM[14498] <= 32'b11111111110000010000000100010011;
ROM[14499] <= 32'b00000000000000010010001110000011;
ROM[14500] <= 32'b00000010011100011010011000100011;
ROM[14501] <= 32'b00000100010100000000001110010011;
ROM[14502] <= 32'b00000000011100010010000000100011;
ROM[14503] <= 32'b00000000010000010000000100010011;
ROM[14504] <= 32'b11111111110000010000000100010011;
ROM[14505] <= 32'b00000000000000010010001110000011;
ROM[14506] <= 32'b00000010011100011010001000100011;
ROM[14507] <= 32'b00000101001100000000001110010011;
ROM[14508] <= 32'b00000000011100010010000000100011;
ROM[14509] <= 32'b00000000010000010000000100010011;
ROM[14510] <= 32'b11111111110000010000000100010011;
ROM[14511] <= 32'b00000000000000010010001110000011;
ROM[14512] <= 32'b00000010011100011010100000100011;
ROM[14513] <= 32'b00000100100000000000001110010011;
ROM[14514] <= 32'b00000000011100010010000000100011;
ROM[14515] <= 32'b00000000010000010000000100010011;
ROM[14516] <= 32'b11111111110000010000000100010011;
ROM[14517] <= 32'b00000000000000010010001110000011;
ROM[14518] <= 32'b00000010011100011010101000100011;
ROM[14519] <= 32'b00000000000100000000001110010011;
ROM[14520] <= 32'b00000000011100010010000000100011;
ROM[14521] <= 32'b00000000010000010000000100010011;
ROM[14522] <= 32'b00000000000000001110001110110111;
ROM[14523] <= 32'b00110011010000111000001110010011;
ROM[14524] <= 32'b00000000111000111000001110110011;
ROM[14525] <= 32'b00000000011100010010000000100011;
ROM[14526] <= 32'b00000000010000010000000100010011;
ROM[14527] <= 32'b00000000001100010010000000100011;
ROM[14528] <= 32'b00000000010000010000000100010011;
ROM[14529] <= 32'b00000000010000010010000000100011;
ROM[14530] <= 32'b00000000010000010000000100010011;
ROM[14531] <= 32'b00000000010100010010000000100011;
ROM[14532] <= 32'b00000000010000010000000100010011;
ROM[14533] <= 32'b00000000011000010010000000100011;
ROM[14534] <= 32'b00000000010000010000000100010011;
ROM[14535] <= 32'b00000001010000000000001110010011;
ROM[14536] <= 32'b00000000010000111000001110010011;
ROM[14537] <= 32'b01000000011100010000001110110011;
ROM[14538] <= 32'b00000000011100000000001000110011;
ROM[14539] <= 32'b00000000001000000000000110110011;
ROM[14540] <= 32'b01000000110000011011000011101111;
ROM[14541] <= 32'b00000010000000000000001110010011;
ROM[14542] <= 32'b00000000011100010010000000100011;
ROM[14543] <= 32'b00000000010000010000000100010011;
ROM[14544] <= 32'b00000000000000001110001110110111;
ROM[14545] <= 32'b00111000110000111000001110010011;
ROM[14546] <= 32'b00000000111000111000001110110011;
ROM[14547] <= 32'b00000000011100010010000000100011;
ROM[14548] <= 32'b00000000010000010000000100010011;
ROM[14549] <= 32'b00000000001100010010000000100011;
ROM[14550] <= 32'b00000000010000010000000100010011;
ROM[14551] <= 32'b00000000010000010010000000100011;
ROM[14552] <= 32'b00000000010000010000000100010011;
ROM[14553] <= 32'b00000000010100010010000000100011;
ROM[14554] <= 32'b00000000010000010000000100010011;
ROM[14555] <= 32'b00000000011000010010000000100011;
ROM[14556] <= 32'b00000000010000010000000100010011;
ROM[14557] <= 32'b00000001010000000000001110010011;
ROM[14558] <= 32'b00000000100000111000001110010011;
ROM[14559] <= 32'b01000000011100010000001110110011;
ROM[14560] <= 32'b00000000011100000000001000110011;
ROM[14561] <= 32'b00000000001000000000000110110011;
ROM[14562] <= 32'b00000010010100011011000011101111;
ROM[14563] <= 32'b11111111110000010000000100010011;
ROM[14564] <= 32'b00000000000000010010001110000011;
ROM[14565] <= 32'b00000000011100011010011000100011;
ROM[14566] <= 32'b00000000010100000000001110010011;
ROM[14567] <= 32'b00000000011100010010000000100011;
ROM[14568] <= 32'b00000000010000010000000100010011;
ROM[14569] <= 32'b00000000000000001110001110110111;
ROM[14570] <= 32'b00111111000000111000001110010011;
ROM[14571] <= 32'b00000000111000111000001110110011;
ROM[14572] <= 32'b00000000011100010010000000100011;
ROM[14573] <= 32'b00000000010000010000000100010011;
ROM[14574] <= 32'b00000000001100010010000000100011;
ROM[14575] <= 32'b00000000010000010000000100010011;
ROM[14576] <= 32'b00000000010000010010000000100011;
ROM[14577] <= 32'b00000000010000010000000100010011;
ROM[14578] <= 32'b00000000010100010010000000100011;
ROM[14579] <= 32'b00000000010000010000000100010011;
ROM[14580] <= 32'b00000000011000010010000000100011;
ROM[14581] <= 32'b00000000010000010000000100010011;
ROM[14582] <= 32'b00000001010000000000001110010011;
ROM[14583] <= 32'b00000000010000111000001110010011;
ROM[14584] <= 32'b01000000011100010000001110110011;
ROM[14585] <= 32'b00000000011100000000001000110011;
ROM[14586] <= 32'b00000000001000000000000110110011;
ROM[14587] <= 32'b00110101000000011011000011101111;
ROM[14588] <= 32'b00000010110100000000001110010011;
ROM[14589] <= 32'b00000000011100010010000000100011;
ROM[14590] <= 32'b00000000010000010000000100010011;
ROM[14591] <= 32'b00000000000000001110001110110111;
ROM[14592] <= 32'b01000100100000111000001110010011;
ROM[14593] <= 32'b00000000111000111000001110110011;
ROM[14594] <= 32'b00000000011100010010000000100011;
ROM[14595] <= 32'b00000000010000010000000100010011;
ROM[14596] <= 32'b00000000001100010010000000100011;
ROM[14597] <= 32'b00000000010000010000000100010011;
ROM[14598] <= 32'b00000000010000010010000000100011;
ROM[14599] <= 32'b00000000010000010000000100010011;
ROM[14600] <= 32'b00000000010100010010000000100011;
ROM[14601] <= 32'b00000000010000010000000100010011;
ROM[14602] <= 32'b00000000011000010010000000100011;
ROM[14603] <= 32'b00000000010000010000000100010011;
ROM[14604] <= 32'b00000001010000000000001110010011;
ROM[14605] <= 32'b00000000100000111000001110010011;
ROM[14606] <= 32'b01000000011100010000001110110011;
ROM[14607] <= 32'b00000000011100000000001000110011;
ROM[14608] <= 32'b00000000001000000000000110110011;
ROM[14609] <= 32'b01110110100000011011000011101111;
ROM[14610] <= 32'b00000010110100000000001110010011;
ROM[14611] <= 32'b00000000011100010010000000100011;
ROM[14612] <= 32'b00000000010000010000000100010011;
ROM[14613] <= 32'b00000000000000001110001110110111;
ROM[14614] <= 32'b01001010000000111000001110010011;
ROM[14615] <= 32'b00000000111000111000001110110011;
ROM[14616] <= 32'b00000000011100010010000000100011;
ROM[14617] <= 32'b00000000010000010000000100010011;
ROM[14618] <= 32'b00000000001100010010000000100011;
ROM[14619] <= 32'b00000000010000010000000100010011;
ROM[14620] <= 32'b00000000010000010010000000100011;
ROM[14621] <= 32'b00000000010000010000000100010011;
ROM[14622] <= 32'b00000000010100010010000000100011;
ROM[14623] <= 32'b00000000010000010000000100010011;
ROM[14624] <= 32'b00000000011000010010000000100011;
ROM[14625] <= 32'b00000000010000010000000100010011;
ROM[14626] <= 32'b00000001010000000000001110010011;
ROM[14627] <= 32'b00000000100000111000001110010011;
ROM[14628] <= 32'b01000000011100010000001110110011;
ROM[14629] <= 32'b00000000011100000000001000110011;
ROM[14630] <= 32'b00000000001000000000000110110011;
ROM[14631] <= 32'b01110001000000011011000011101111;
ROM[14632] <= 32'b00000010110100000000001110010011;
ROM[14633] <= 32'b00000000011100010010000000100011;
ROM[14634] <= 32'b00000000010000010000000100010011;
ROM[14635] <= 32'b00000000000000001110001110110111;
ROM[14636] <= 32'b01001111100000111000001110010011;
ROM[14637] <= 32'b00000000111000111000001110110011;
ROM[14638] <= 32'b00000000011100010010000000100011;
ROM[14639] <= 32'b00000000010000010000000100010011;
ROM[14640] <= 32'b00000000001100010010000000100011;
ROM[14641] <= 32'b00000000010000010000000100010011;
ROM[14642] <= 32'b00000000010000010010000000100011;
ROM[14643] <= 32'b00000000010000010000000100010011;
ROM[14644] <= 32'b00000000010100010010000000100011;
ROM[14645] <= 32'b00000000010000010000000100010011;
ROM[14646] <= 32'b00000000011000010010000000100011;
ROM[14647] <= 32'b00000000010000010000000100010011;
ROM[14648] <= 32'b00000001010000000000001110010011;
ROM[14649] <= 32'b00000000100000111000001110010011;
ROM[14650] <= 32'b01000000011100010000001110110011;
ROM[14651] <= 32'b00000000011100000000001000110011;
ROM[14652] <= 32'b00000000001000000000000110110011;
ROM[14653] <= 32'b01101011100000011011000011101111;
ROM[14654] <= 32'b00000011111000000000001110010011;
ROM[14655] <= 32'b00000000011100010010000000100011;
ROM[14656] <= 32'b00000000010000010000000100010011;
ROM[14657] <= 32'b00000000000000001110001110110111;
ROM[14658] <= 32'b01010101000000111000001110010011;
ROM[14659] <= 32'b00000000111000111000001110110011;
ROM[14660] <= 32'b00000000011100010010000000100011;
ROM[14661] <= 32'b00000000010000010000000100010011;
ROM[14662] <= 32'b00000000001100010010000000100011;
ROM[14663] <= 32'b00000000010000010000000100010011;
ROM[14664] <= 32'b00000000010000010010000000100011;
ROM[14665] <= 32'b00000000010000010000000100010011;
ROM[14666] <= 32'b00000000010100010010000000100011;
ROM[14667] <= 32'b00000000010000010000000100010011;
ROM[14668] <= 32'b00000000011000010010000000100011;
ROM[14669] <= 32'b00000000010000010000000100010011;
ROM[14670] <= 32'b00000001010000000000001110010011;
ROM[14671] <= 32'b00000000100000111000001110010011;
ROM[14672] <= 32'b01000000011100010000001110110011;
ROM[14673] <= 32'b00000000011100000000001000110011;
ROM[14674] <= 32'b00000000001000000000000110110011;
ROM[14675] <= 32'b01100110000000011011000011101111;
ROM[14676] <= 32'b00000010000000000000001110010011;
ROM[14677] <= 32'b00000000011100010010000000100011;
ROM[14678] <= 32'b00000000010000010000000100010011;
ROM[14679] <= 32'b00000000000000001110001110110111;
ROM[14680] <= 32'b01011010100000111000001110010011;
ROM[14681] <= 32'b00000000111000111000001110110011;
ROM[14682] <= 32'b00000000011100010010000000100011;
ROM[14683] <= 32'b00000000010000010000000100010011;
ROM[14684] <= 32'b00000000001100010010000000100011;
ROM[14685] <= 32'b00000000010000010000000100010011;
ROM[14686] <= 32'b00000000010000010010000000100011;
ROM[14687] <= 32'b00000000010000010000000100010011;
ROM[14688] <= 32'b00000000010100010010000000100011;
ROM[14689] <= 32'b00000000010000010000000100010011;
ROM[14690] <= 32'b00000000011000010010000000100011;
ROM[14691] <= 32'b00000000010000010000000100010011;
ROM[14692] <= 32'b00000001010000000000001110010011;
ROM[14693] <= 32'b00000000100000111000001110010011;
ROM[14694] <= 32'b01000000011100010000001110110011;
ROM[14695] <= 32'b00000000011100000000001000110011;
ROM[14696] <= 32'b00000000001000000000000110110011;
ROM[14697] <= 32'b01100000100000011011000011101111;
ROM[14698] <= 32'b11111111110000010000000100010011;
ROM[14699] <= 32'b00000000000000010010001110000011;
ROM[14700] <= 32'b00000000011100011010010000100011;
ROM[14701] <= 32'b00000000111100000000001110010011;
ROM[14702] <= 32'b00000000011100010010000000100011;
ROM[14703] <= 32'b00000000010000010000000100010011;
ROM[14704] <= 32'b00000000000000001110001110110111;
ROM[14705] <= 32'b01100000110000111000001110010011;
ROM[14706] <= 32'b00000000111000111000001110110011;
ROM[14707] <= 32'b00000000011100010010000000100011;
ROM[14708] <= 32'b00000000010000010000000100010011;
ROM[14709] <= 32'b00000000001100010010000000100011;
ROM[14710] <= 32'b00000000010000010000000100010011;
ROM[14711] <= 32'b00000000010000010010000000100011;
ROM[14712] <= 32'b00000000010000010000000100010011;
ROM[14713] <= 32'b00000000010100010010000000100011;
ROM[14714] <= 32'b00000000010000010000000100010011;
ROM[14715] <= 32'b00000000011000010010000000100011;
ROM[14716] <= 32'b00000000010000010000000100010011;
ROM[14717] <= 32'b00000001010000000000001110010011;
ROM[14718] <= 32'b00000000010000111000001110010011;
ROM[14719] <= 32'b01000000011100010000001110110011;
ROM[14720] <= 32'b00000000011100000000001000110011;
ROM[14721] <= 32'b00000000001000000000000110110011;
ROM[14722] <= 32'b00010011010000011011000011101111;
ROM[14723] <= 32'b00000110100100000000001110010011;
ROM[14724] <= 32'b00000000011100010010000000100011;
ROM[14725] <= 32'b00000000010000010000000100010011;
ROM[14726] <= 32'b00000000000000001110001110110111;
ROM[14727] <= 32'b01100110010000111000001110010011;
ROM[14728] <= 32'b00000000111000111000001110110011;
ROM[14729] <= 32'b00000000011100010010000000100011;
ROM[14730] <= 32'b00000000010000010000000100010011;
ROM[14731] <= 32'b00000000001100010010000000100011;
ROM[14732] <= 32'b00000000010000010000000100010011;
ROM[14733] <= 32'b00000000010000010010000000100011;
ROM[14734] <= 32'b00000000010000010000000100010011;
ROM[14735] <= 32'b00000000010100010010000000100011;
ROM[14736] <= 32'b00000000010000010000000100010011;
ROM[14737] <= 32'b00000000011000010010000000100011;
ROM[14738] <= 32'b00000000010000010000000100010011;
ROM[14739] <= 32'b00000001010000000000001110010011;
ROM[14740] <= 32'b00000000100000111000001110010011;
ROM[14741] <= 32'b01000000011100010000001110110011;
ROM[14742] <= 32'b00000000011100000000001000110011;
ROM[14743] <= 32'b00000000001000000000000110110011;
ROM[14744] <= 32'b01010100110000011011000011101111;
ROM[14745] <= 32'b00000110111000000000001110010011;
ROM[14746] <= 32'b00000000011100010010000000100011;
ROM[14747] <= 32'b00000000010000010000000100010011;
ROM[14748] <= 32'b00000000000000001110001110110111;
ROM[14749] <= 32'b01101011110000111000001110010011;
ROM[14750] <= 32'b00000000111000111000001110110011;
ROM[14751] <= 32'b00000000011100010010000000100011;
ROM[14752] <= 32'b00000000010000010000000100010011;
ROM[14753] <= 32'b00000000001100010010000000100011;
ROM[14754] <= 32'b00000000010000010000000100010011;
ROM[14755] <= 32'b00000000010000010010000000100011;
ROM[14756] <= 32'b00000000010000010000000100010011;
ROM[14757] <= 32'b00000000010100010010000000100011;
ROM[14758] <= 32'b00000000010000010000000100010011;
ROM[14759] <= 32'b00000000011000010010000000100011;
ROM[14760] <= 32'b00000000010000010000000100010011;
ROM[14761] <= 32'b00000001010000000000001110010011;
ROM[14762] <= 32'b00000000100000111000001110010011;
ROM[14763] <= 32'b01000000011100010000001110110011;
ROM[14764] <= 32'b00000000011100000000001000110011;
ROM[14765] <= 32'b00000000001000000000000110110011;
ROM[14766] <= 32'b01001111010000011011000011101111;
ROM[14767] <= 32'b00000111011000000000001110010011;
ROM[14768] <= 32'b00000000011100010010000000100011;
ROM[14769] <= 32'b00000000010000010000000100010011;
ROM[14770] <= 32'b00000000000000001110001110110111;
ROM[14771] <= 32'b01110001010000111000001110010011;
ROM[14772] <= 32'b00000000111000111000001110110011;
ROM[14773] <= 32'b00000000011100010010000000100011;
ROM[14774] <= 32'b00000000010000010000000100010011;
ROM[14775] <= 32'b00000000001100010010000000100011;
ROM[14776] <= 32'b00000000010000010000000100010011;
ROM[14777] <= 32'b00000000010000010010000000100011;
ROM[14778] <= 32'b00000000010000010000000100010011;
ROM[14779] <= 32'b00000000010100010010000000100011;
ROM[14780] <= 32'b00000000010000010000000100010011;
ROM[14781] <= 32'b00000000011000010010000000100011;
ROM[14782] <= 32'b00000000010000010000000100010011;
ROM[14783] <= 32'b00000001010000000000001110010011;
ROM[14784] <= 32'b00000000100000111000001110010011;
ROM[14785] <= 32'b01000000011100010000001110110011;
ROM[14786] <= 32'b00000000011100000000001000110011;
ROM[14787] <= 32'b00000000001000000000000110110011;
ROM[14788] <= 32'b01001001110000011011000011101111;
ROM[14789] <= 32'b00000110000100000000001110010011;
ROM[14790] <= 32'b00000000011100010010000000100011;
ROM[14791] <= 32'b00000000010000010000000100010011;
ROM[14792] <= 32'b00000000000000001110001110110111;
ROM[14793] <= 32'b01110110110000111000001110010011;
ROM[14794] <= 32'b00000000111000111000001110110011;
ROM[14795] <= 32'b00000000011100010010000000100011;
ROM[14796] <= 32'b00000000010000010000000100010011;
ROM[14797] <= 32'b00000000001100010010000000100011;
ROM[14798] <= 32'b00000000010000010000000100010011;
ROM[14799] <= 32'b00000000010000010010000000100011;
ROM[14800] <= 32'b00000000010000010000000100010011;
ROM[14801] <= 32'b00000000010100010010000000100011;
ROM[14802] <= 32'b00000000010000010000000100010011;
ROM[14803] <= 32'b00000000011000010010000000100011;
ROM[14804] <= 32'b00000000010000010000000100010011;
ROM[14805] <= 32'b00000001010000000000001110010011;
ROM[14806] <= 32'b00000000100000111000001110010011;
ROM[14807] <= 32'b01000000011100010000001110110011;
ROM[14808] <= 32'b00000000011100000000001000110011;
ROM[14809] <= 32'b00000000001000000000000110110011;
ROM[14810] <= 32'b01000100010000011011000011101111;
ROM[14811] <= 32'b00000110110000000000001110010011;
ROM[14812] <= 32'b00000000011100010010000000100011;
ROM[14813] <= 32'b00000000010000010000000100010011;
ROM[14814] <= 32'b00000000000000001110001110110111;
ROM[14815] <= 32'b01111100010000111000001110010011;
ROM[14816] <= 32'b00000000111000111000001110110011;
ROM[14817] <= 32'b00000000011100010010000000100011;
ROM[14818] <= 32'b00000000010000010000000100010011;
ROM[14819] <= 32'b00000000001100010010000000100011;
ROM[14820] <= 32'b00000000010000010000000100010011;
ROM[14821] <= 32'b00000000010000010010000000100011;
ROM[14822] <= 32'b00000000010000010000000100010011;
ROM[14823] <= 32'b00000000010100010010000000100011;
ROM[14824] <= 32'b00000000010000010000000100010011;
ROM[14825] <= 32'b00000000011000010010000000100011;
ROM[14826] <= 32'b00000000010000010000000100010011;
ROM[14827] <= 32'b00000001010000000000001110010011;
ROM[14828] <= 32'b00000000100000111000001110010011;
ROM[14829] <= 32'b01000000011100010000001110110011;
ROM[14830] <= 32'b00000000011100000000001000110011;
ROM[14831] <= 32'b00000000001000000000000110110011;
ROM[14832] <= 32'b00111110110000011011000011101111;
ROM[14833] <= 32'b00000110100100000000001110010011;
ROM[14834] <= 32'b00000000011100010010000000100011;
ROM[14835] <= 32'b00000000010000010000000100010011;
ROM[14836] <= 32'b00000000000000001111001110110111;
ROM[14837] <= 32'b10000001110000111000001110010011;
ROM[14838] <= 32'b00000000111000111000001110110011;
ROM[14839] <= 32'b00000000011100010010000000100011;
ROM[14840] <= 32'b00000000010000010000000100010011;
ROM[14841] <= 32'b00000000001100010010000000100011;
ROM[14842] <= 32'b00000000010000010000000100010011;
ROM[14843] <= 32'b00000000010000010010000000100011;
ROM[14844] <= 32'b00000000010000010000000100010011;
ROM[14845] <= 32'b00000000010100010010000000100011;
ROM[14846] <= 32'b00000000010000010000000100010011;
ROM[14847] <= 32'b00000000011000010010000000100011;
ROM[14848] <= 32'b00000000010000010000000100010011;
ROM[14849] <= 32'b00000001010000000000001110010011;
ROM[14850] <= 32'b00000000100000111000001110010011;
ROM[14851] <= 32'b01000000011100010000001110110011;
ROM[14852] <= 32'b00000000011100000000001000110011;
ROM[14853] <= 32'b00000000001000000000000110110011;
ROM[14854] <= 32'b00111001010000011011000011101111;
ROM[14855] <= 32'b00000110010000000000001110010011;
ROM[14856] <= 32'b00000000011100010010000000100011;
ROM[14857] <= 32'b00000000010000010000000100010011;
ROM[14858] <= 32'b00000000000000001111001110110111;
ROM[14859] <= 32'b10000111010000111000001110010011;
ROM[14860] <= 32'b00000000111000111000001110110011;
ROM[14861] <= 32'b00000000011100010010000000100011;
ROM[14862] <= 32'b00000000010000010000000100010011;
ROM[14863] <= 32'b00000000001100010010000000100011;
ROM[14864] <= 32'b00000000010000010000000100010011;
ROM[14865] <= 32'b00000000010000010010000000100011;
ROM[14866] <= 32'b00000000010000010000000100010011;
ROM[14867] <= 32'b00000000010100010010000000100011;
ROM[14868] <= 32'b00000000010000010000000100010011;
ROM[14869] <= 32'b00000000011000010010000000100011;
ROM[14870] <= 32'b00000000010000010000000100010011;
ROM[14871] <= 32'b00000001010000000000001110010011;
ROM[14872] <= 32'b00000000100000111000001110010011;
ROM[14873] <= 32'b01000000011100010000001110110011;
ROM[14874] <= 32'b00000000011100000000001000110011;
ROM[14875] <= 32'b00000000001000000000000110110011;
ROM[14876] <= 32'b00110011110000011011000011101111;
ROM[14877] <= 32'b00000010000000000000001110010011;
ROM[14878] <= 32'b00000000011100010010000000100011;
ROM[14879] <= 32'b00000000010000010000000100010011;
ROM[14880] <= 32'b00000000000000001111001110110111;
ROM[14881] <= 32'b10001100110000111000001110010011;
ROM[14882] <= 32'b00000000111000111000001110110011;
ROM[14883] <= 32'b00000000011100010010000000100011;
ROM[14884] <= 32'b00000000010000010000000100010011;
ROM[14885] <= 32'b00000000001100010010000000100011;
ROM[14886] <= 32'b00000000010000010000000100010011;
ROM[14887] <= 32'b00000000010000010010000000100011;
ROM[14888] <= 32'b00000000010000010000000100010011;
ROM[14889] <= 32'b00000000010100010010000000100011;
ROM[14890] <= 32'b00000000010000010000000100010011;
ROM[14891] <= 32'b00000000011000010010000000100011;
ROM[14892] <= 32'b00000000010000010000000100010011;
ROM[14893] <= 32'b00000001010000000000001110010011;
ROM[14894] <= 32'b00000000100000111000001110010011;
ROM[14895] <= 32'b01000000011100010000001110110011;
ROM[14896] <= 32'b00000000011100000000001000110011;
ROM[14897] <= 32'b00000000001000000000000110110011;
ROM[14898] <= 32'b00101110010000011011000011101111;
ROM[14899] <= 32'b00000110001100000000001110010011;
ROM[14900] <= 32'b00000000011100010010000000100011;
ROM[14901] <= 32'b00000000010000010000000100010011;
ROM[14902] <= 32'b00000000000000001111001110110111;
ROM[14903] <= 32'b10010010010000111000001110010011;
ROM[14904] <= 32'b00000000111000111000001110110011;
ROM[14905] <= 32'b00000000011100010010000000100011;
ROM[14906] <= 32'b00000000010000010000000100010011;
ROM[14907] <= 32'b00000000001100010010000000100011;
ROM[14908] <= 32'b00000000010000010000000100010011;
ROM[14909] <= 32'b00000000010000010010000000100011;
ROM[14910] <= 32'b00000000010000010000000100010011;
ROM[14911] <= 32'b00000000010100010010000000100011;
ROM[14912] <= 32'b00000000010000010000000100010011;
ROM[14913] <= 32'b00000000011000010010000000100011;
ROM[14914] <= 32'b00000000010000010000000100010011;
ROM[14915] <= 32'b00000001010000000000001110010011;
ROM[14916] <= 32'b00000000100000111000001110010011;
ROM[14917] <= 32'b01000000011100010000001110110011;
ROM[14918] <= 32'b00000000011100000000001000110011;
ROM[14919] <= 32'b00000000001000000000000110110011;
ROM[14920] <= 32'b00101000110000011011000011101111;
ROM[14921] <= 32'b00000110111100000000001110010011;
ROM[14922] <= 32'b00000000011100010010000000100011;
ROM[14923] <= 32'b00000000010000010000000100010011;
ROM[14924] <= 32'b00000000000000001111001110110111;
ROM[14925] <= 32'b10010111110000111000001110010011;
ROM[14926] <= 32'b00000000111000111000001110110011;
ROM[14927] <= 32'b00000000011100010010000000100011;
ROM[14928] <= 32'b00000000010000010000000100010011;
ROM[14929] <= 32'b00000000001100010010000000100011;
ROM[14930] <= 32'b00000000010000010000000100010011;
ROM[14931] <= 32'b00000000010000010010000000100011;
ROM[14932] <= 32'b00000000010000010000000100010011;
ROM[14933] <= 32'b00000000010100010010000000100011;
ROM[14934] <= 32'b00000000010000010000000100010011;
ROM[14935] <= 32'b00000000011000010010000000100011;
ROM[14936] <= 32'b00000000010000010000000100010011;
ROM[14937] <= 32'b00000001010000000000001110010011;
ROM[14938] <= 32'b00000000100000111000001110010011;
ROM[14939] <= 32'b01000000011100010000001110110011;
ROM[14940] <= 32'b00000000011100000000001000110011;
ROM[14941] <= 32'b00000000001000000000000110110011;
ROM[14942] <= 32'b00100011010000011011000011101111;
ROM[14943] <= 32'b00000110110100000000001110010011;
ROM[14944] <= 32'b00000000011100010010000000100011;
ROM[14945] <= 32'b00000000010000010000000100010011;
ROM[14946] <= 32'b00000000000000001111001110110111;
ROM[14947] <= 32'b10011101010000111000001110010011;
ROM[14948] <= 32'b00000000111000111000001110110011;
ROM[14949] <= 32'b00000000011100010010000000100011;
ROM[14950] <= 32'b00000000010000010000000100010011;
ROM[14951] <= 32'b00000000001100010010000000100011;
ROM[14952] <= 32'b00000000010000010000000100010011;
ROM[14953] <= 32'b00000000010000010010000000100011;
ROM[14954] <= 32'b00000000010000010000000100010011;
ROM[14955] <= 32'b00000000010100010010000000100011;
ROM[14956] <= 32'b00000000010000010000000100010011;
ROM[14957] <= 32'b00000000011000010010000000100011;
ROM[14958] <= 32'b00000000010000010000000100010011;
ROM[14959] <= 32'b00000001010000000000001110010011;
ROM[14960] <= 32'b00000000100000111000001110010011;
ROM[14961] <= 32'b01000000011100010000001110110011;
ROM[14962] <= 32'b00000000011100000000001000110011;
ROM[14963] <= 32'b00000000001000000000000110110011;
ROM[14964] <= 32'b00011101110000011011000011101111;
ROM[14965] <= 32'b00000110110100000000001110010011;
ROM[14966] <= 32'b00000000011100010010000000100011;
ROM[14967] <= 32'b00000000010000010000000100010011;
ROM[14968] <= 32'b00000000000000001111001110110111;
ROM[14969] <= 32'b10100010110000111000001110010011;
ROM[14970] <= 32'b00000000111000111000001110110011;
ROM[14971] <= 32'b00000000011100010010000000100011;
ROM[14972] <= 32'b00000000010000010000000100010011;
ROM[14973] <= 32'b00000000001100010010000000100011;
ROM[14974] <= 32'b00000000010000010000000100010011;
ROM[14975] <= 32'b00000000010000010010000000100011;
ROM[14976] <= 32'b00000000010000010000000100010011;
ROM[14977] <= 32'b00000000010100010010000000100011;
ROM[14978] <= 32'b00000000010000010000000100010011;
ROM[14979] <= 32'b00000000011000010010000000100011;
ROM[14980] <= 32'b00000000010000010000000100010011;
ROM[14981] <= 32'b00000001010000000000001110010011;
ROM[14982] <= 32'b00000000100000111000001110010011;
ROM[14983] <= 32'b01000000011100010000001110110011;
ROM[14984] <= 32'b00000000011100000000001000110011;
ROM[14985] <= 32'b00000000001000000000000110110011;
ROM[14986] <= 32'b00011000010000011011000011101111;
ROM[14987] <= 32'b00000110000100000000001110010011;
ROM[14988] <= 32'b00000000011100010010000000100011;
ROM[14989] <= 32'b00000000010000010000000100010011;
ROM[14990] <= 32'b00000000000000001111001110110111;
ROM[14991] <= 32'b10101000010000111000001110010011;
ROM[14992] <= 32'b00000000111000111000001110110011;
ROM[14993] <= 32'b00000000011100010010000000100011;
ROM[14994] <= 32'b00000000010000010000000100010011;
ROM[14995] <= 32'b00000000001100010010000000100011;
ROM[14996] <= 32'b00000000010000010000000100010011;
ROM[14997] <= 32'b00000000010000010010000000100011;
ROM[14998] <= 32'b00000000010000010000000100010011;
ROM[14999] <= 32'b00000000010100010010000000100011;
ROM[15000] <= 32'b00000000010000010000000100010011;
ROM[15001] <= 32'b00000000011000010010000000100011;
ROM[15002] <= 32'b00000000010000010000000100010011;
ROM[15003] <= 32'b00000001010000000000001110010011;
ROM[15004] <= 32'b00000000100000111000001110010011;
ROM[15005] <= 32'b01000000011100010000001110110011;
ROM[15006] <= 32'b00000000011100000000001000110011;
ROM[15007] <= 32'b00000000001000000000000110110011;
ROM[15008] <= 32'b00010010110000011011000011101111;
ROM[15009] <= 32'b00000110111000000000001110010011;
ROM[15010] <= 32'b00000000011100010010000000100011;
ROM[15011] <= 32'b00000000010000010000000100010011;
ROM[15012] <= 32'b00000000000000001111001110110111;
ROM[15013] <= 32'b10101101110000111000001110010011;
ROM[15014] <= 32'b00000000111000111000001110110011;
ROM[15015] <= 32'b00000000011100010010000000100011;
ROM[15016] <= 32'b00000000010000010000000100010011;
ROM[15017] <= 32'b00000000001100010010000000100011;
ROM[15018] <= 32'b00000000010000010000000100010011;
ROM[15019] <= 32'b00000000010000010010000000100011;
ROM[15020] <= 32'b00000000010000010000000100010011;
ROM[15021] <= 32'b00000000010100010010000000100011;
ROM[15022] <= 32'b00000000010000010000000100010011;
ROM[15023] <= 32'b00000000011000010010000000100011;
ROM[15024] <= 32'b00000000010000010000000100010011;
ROM[15025] <= 32'b00000001010000000000001110010011;
ROM[15026] <= 32'b00000000100000111000001110010011;
ROM[15027] <= 32'b01000000011100010000001110110011;
ROM[15028] <= 32'b00000000011100000000001000110011;
ROM[15029] <= 32'b00000000001000000000000110110011;
ROM[15030] <= 32'b00001101010000011011000011101111;
ROM[15031] <= 32'b00000110010000000000001110010011;
ROM[15032] <= 32'b00000000011100010010000000100011;
ROM[15033] <= 32'b00000000010000010000000100010011;
ROM[15034] <= 32'b00000000000000001111001110110111;
ROM[15035] <= 32'b10110011010000111000001110010011;
ROM[15036] <= 32'b00000000111000111000001110110011;
ROM[15037] <= 32'b00000000011100010010000000100011;
ROM[15038] <= 32'b00000000010000010000000100010011;
ROM[15039] <= 32'b00000000001100010010000000100011;
ROM[15040] <= 32'b00000000010000010000000100010011;
ROM[15041] <= 32'b00000000010000010010000000100011;
ROM[15042] <= 32'b00000000010000010000000100010011;
ROM[15043] <= 32'b00000000010100010010000000100011;
ROM[15044] <= 32'b00000000010000010000000100010011;
ROM[15045] <= 32'b00000000011000010010000000100011;
ROM[15046] <= 32'b00000000010000010000000100010011;
ROM[15047] <= 32'b00000001010000000000001110010011;
ROM[15048] <= 32'b00000000100000111000001110010011;
ROM[15049] <= 32'b01000000011100010000001110110011;
ROM[15050] <= 32'b00000000011100000000001000110011;
ROM[15051] <= 32'b00000000001000000000000110110011;
ROM[15052] <= 32'b00000111110000011011000011101111;
ROM[15053] <= 32'b11111111110000010000000100010011;
ROM[15054] <= 32'b00000000000000010010001110000011;
ROM[15055] <= 32'b00000000011100011010100000100011;
ROM[15056] <= 32'b00000000000000000000001110010011;
ROM[15057] <= 32'b00000000011100010010000000100011;
ROM[15058] <= 32'b00000000010000010000000100010011;
ROM[15059] <= 32'b11111111110000010000000100010011;
ROM[15060] <= 32'b00000000000000010010001110000011;
ROM[15061] <= 32'b00000000011100011010000000100011;
ROM[15062] <= 32'b00000000000100000000001110010011;
ROM[15063] <= 32'b00000000011100010010000000100011;
ROM[15064] <= 32'b00000000010000010000000100010011;
ROM[15065] <= 32'b11111111110000010000000100010011;
ROM[15066] <= 32'b00000000000000010010001110000011;
ROM[15067] <= 32'b00000000011100011010001000100011;
ROM[15068] <= 32'b00000000000000011010001110000011;
ROM[15069] <= 32'b00000000011100010010000000100011;
ROM[15070] <= 32'b00000000010000010000000100010011;
ROM[15071] <= 32'b00000000010000011010001110000011;
ROM[15072] <= 32'b00000000011100010010000000100011;
ROM[15073] <= 32'b00000000010000010000000100010011;
ROM[15074] <= 32'b11111111110000010000000100010011;
ROM[15075] <= 32'b00000000000000010010001110000011;
ROM[15076] <= 32'b11111111110000010000000100010011;
ROM[15077] <= 32'b00000000000000010010010000000011;
ROM[15078] <= 32'b00000000011101000010001110110011;
ROM[15079] <= 32'b00000000011100010010000000100011;
ROM[15080] <= 32'b00000000010000010000000100010011;
ROM[15081] <= 32'b11111111110000010000000100010011;
ROM[15082] <= 32'b00000000000000010010001110000011;
ROM[15083] <= 32'b01000000011100000000001110110011;
ROM[15084] <= 32'b00000000000100111000001110010011;
ROM[15085] <= 32'b00000000011100010010000000100011;
ROM[15086] <= 32'b00000000010000010000000100010011;
ROM[15087] <= 32'b11111111110000010000000100010011;
ROM[15088] <= 32'b00000000000000010010001110000011;
ROM[15089] <= 32'b00000000000000111000101001100011;
ROM[15090] <= 32'b00000000000000010000001110110111;
ROM[15091] <= 32'b00001000000000111000001110010011;
ROM[15092] <= 32'b00000000111000111000001110110011;
ROM[15093] <= 32'b00000000000000111000000011100111;
ROM[15094] <= 32'b00000000100000011010001110000011;
ROM[15095] <= 32'b00000000011100010010000000100011;
ROM[15096] <= 32'b00000000010000010000000100010011;
ROM[15097] <= 32'b00000000000000001111001110110111;
ROM[15098] <= 32'b11000011000000111000001110010011;
ROM[15099] <= 32'b00000000111000111000001110110011;
ROM[15100] <= 32'b00000000011100010010000000100011;
ROM[15101] <= 32'b00000000010000010000000100010011;
ROM[15102] <= 32'b00000000001100010010000000100011;
ROM[15103] <= 32'b00000000010000010000000100010011;
ROM[15104] <= 32'b00000000010000010010000000100011;
ROM[15105] <= 32'b00000000010000010000000100010011;
ROM[15106] <= 32'b00000000010100010010000000100011;
ROM[15107] <= 32'b00000000010000010000000100010011;
ROM[15108] <= 32'b00000000011000010010000000100011;
ROM[15109] <= 32'b00000000010000010000000100010011;
ROM[15110] <= 32'b00000001010000000000001110010011;
ROM[15111] <= 32'b00000000010000111000001110010011;
ROM[15112] <= 32'b01000000011100010000001110110011;
ROM[15113] <= 32'b00000000011100000000001000110011;
ROM[15114] <= 32'b00000000001000000000000110110011;
ROM[15115] <= 32'b11111011110111111110000011101111;
ROM[15116] <= 32'b11111111110000010000000100010011;
ROM[15117] <= 32'b00000000000000010010001110000011;
ROM[15118] <= 32'b00000000011100011010101000100011;
ROM[15119] <= 32'b00000001010000011010001110000011;
ROM[15120] <= 32'b00000000011100010010000000100011;
ROM[15121] <= 32'b00000000010000010000000100010011;
ROM[15122] <= 32'b00000000000000000000001110010011;
ROM[15123] <= 32'b00000000011100010010000000100011;
ROM[15124] <= 32'b00000000010000010000000100010011;
ROM[15125] <= 32'b00000000000000001111001110110111;
ROM[15126] <= 32'b11001010000000111000001110010011;
ROM[15127] <= 32'b00000000111000111000001110110011;
ROM[15128] <= 32'b00000000011100010010000000100011;
ROM[15129] <= 32'b00000000010000010000000100010011;
ROM[15130] <= 32'b00000000001100010010000000100011;
ROM[15131] <= 32'b00000000010000010000000100010011;
ROM[15132] <= 32'b00000000010000010010000000100011;
ROM[15133] <= 32'b00000000010000010000000100010011;
ROM[15134] <= 32'b00000000010100010010000000100011;
ROM[15135] <= 32'b00000000010000010000000100010011;
ROM[15136] <= 32'b00000000011000010010000000100011;
ROM[15137] <= 32'b00000000010000010000000100010011;
ROM[15138] <= 32'b00000001010000000000001110010011;
ROM[15139] <= 32'b00000000100000111000001110010011;
ROM[15140] <= 32'b01000000011100010000001110110011;
ROM[15141] <= 32'b00000000011100000000001000110011;
ROM[15142] <= 32'b00000000001000000000000110110011;
ROM[15143] <= 32'b01001100000100011010000011101111;
ROM[15144] <= 32'b11111111110000010000000100010011;
ROM[15145] <= 32'b00000000000000010010001110000011;
ROM[15146] <= 32'b00000000011100011010110000100011;
ROM[15147] <= 32'b00000001100000011010001110000011;
ROM[15148] <= 32'b00000000011100010010000000100011;
ROM[15149] <= 32'b00000000010000010000000100010011;
ROM[15150] <= 32'b00000001110000011010001110000011;
ROM[15151] <= 32'b00000000011100010010000000100011;
ROM[15152] <= 32'b00000000010000010000000100010011;
ROM[15153] <= 32'b11111111110000010000000100010011;
ROM[15154] <= 32'b00000000000000010010001110000011;
ROM[15155] <= 32'b11111111110000010000000100010011;
ROM[15156] <= 32'b00000000000000010010010000000011;
ROM[15157] <= 32'b00000000011101000010010010110011;
ROM[15158] <= 32'b00000000100000111010010100110011;
ROM[15159] <= 32'b00000000101001001000001110110011;
ROM[15160] <= 32'b00000000000100111000001110010011;
ROM[15161] <= 32'b00000000000100111111001110010011;
ROM[15162] <= 32'b00000000011100010010000000100011;
ROM[15163] <= 32'b00000000010000010000000100010011;
ROM[15164] <= 32'b11111111110000010000000100010011;
ROM[15165] <= 32'b00000000000000010010001110000011;
ROM[15166] <= 32'b00000000000000111000101001100011;
ROM[15167] <= 32'b00000000000000001111001110110111;
ROM[15168] <= 32'b00100000110000111000001110010011;
ROM[15169] <= 32'b00000000111000111000001110110011;
ROM[15170] <= 32'b00000000000000111000000011100111;
ROM[15171] <= 32'b00000001100000011010001110000011;
ROM[15172] <= 32'b00000000011100010010000000100011;
ROM[15173] <= 32'b00000000010000010000000100010011;
ROM[15174] <= 32'b00000010000000011010001110000011;
ROM[15175] <= 32'b00000000011100010010000000100011;
ROM[15176] <= 32'b00000000010000010000000100010011;
ROM[15177] <= 32'b11111111110000010000000100010011;
ROM[15178] <= 32'b00000000000000010010001110000011;
ROM[15179] <= 32'b11111111110000010000000100010011;
ROM[15180] <= 32'b00000000000000010010010000000011;
ROM[15181] <= 32'b00000000011101000010010010110011;
ROM[15182] <= 32'b00000000100000111010010100110011;
ROM[15183] <= 32'b00000000101001001000001110110011;
ROM[15184] <= 32'b00000000000100111000001110010011;
ROM[15185] <= 32'b00000000000100111111001110010011;
ROM[15186] <= 32'b00000000011100010010000000100011;
ROM[15187] <= 32'b00000000010000010000000100010011;
ROM[15188] <= 32'b11111111110000010000000100010011;
ROM[15189] <= 32'b00000000000000010010001110000011;
ROM[15190] <= 32'b00000000000000111000101001100011;
ROM[15191] <= 32'b00000000000000001111001110110111;
ROM[15192] <= 32'b00010100000000111000001110010011;
ROM[15193] <= 32'b00000000111000111000001110110011;
ROM[15194] <= 32'b00000000000000111000000011100111;
ROM[15195] <= 32'b00000001100000011010001110000011;
ROM[15196] <= 32'b00000000011100010010000000100011;
ROM[15197] <= 32'b00000000010000010000000100010011;
ROM[15198] <= 32'b00000010010000011010001110000011;
ROM[15199] <= 32'b00000000011100010010000000100011;
ROM[15200] <= 32'b00000000010000010000000100010011;
ROM[15201] <= 32'b11111111110000010000000100010011;
ROM[15202] <= 32'b00000000000000010010001110000011;
ROM[15203] <= 32'b11111111110000010000000100010011;
ROM[15204] <= 32'b00000000000000010010010000000011;
ROM[15205] <= 32'b00000000011101000010010010110011;
ROM[15206] <= 32'b00000000100000111010010100110011;
ROM[15207] <= 32'b00000000101001001000001110110011;
ROM[15208] <= 32'b00000000000100111000001110010011;
ROM[15209] <= 32'b00000000000100111111001110010011;
ROM[15210] <= 32'b00000000011100010010000000100011;
ROM[15211] <= 32'b00000000010000010000000100010011;
ROM[15212] <= 32'b11111111110000010000000100010011;
ROM[15213] <= 32'b00000000000000010010001110000011;
ROM[15214] <= 32'b00000000000000111000101001100011;
ROM[15215] <= 32'b00000000000000001111001110110111;
ROM[15216] <= 32'b00010010010000111000001110010011;
ROM[15217] <= 32'b00000000111000111000001110110011;
ROM[15218] <= 32'b00000000000000111000000011100111;
ROM[15219] <= 32'b00000001100000011010001110000011;
ROM[15220] <= 32'b00000000011100010010000000100011;
ROM[15221] <= 32'b00000000010000010000000100010011;
ROM[15222] <= 32'b00000010100000011010001110000011;
ROM[15223] <= 32'b00000000011100010010000000100011;
ROM[15224] <= 32'b00000000010000010000000100010011;
ROM[15225] <= 32'b11111111110000010000000100010011;
ROM[15226] <= 32'b00000000000000010010001110000011;
ROM[15227] <= 32'b11111111110000010000000100010011;
ROM[15228] <= 32'b00000000000000010010010000000011;
ROM[15229] <= 32'b00000000011101000010010010110011;
ROM[15230] <= 32'b00000000100000111010010100110011;
ROM[15231] <= 32'b00000000101001001000001110110011;
ROM[15232] <= 32'b00000000000100111000001110010011;
ROM[15233] <= 32'b00000000000100111111001110010011;
ROM[15234] <= 32'b00000000011100010010000000100011;
ROM[15235] <= 32'b00000000010000010000000100010011;
ROM[15236] <= 32'b11111111110000010000000100010011;
ROM[15237] <= 32'b00000000000000010010001110000011;
ROM[15238] <= 32'b00000000000000111000101001100011;
ROM[15239] <= 32'b00000000000000001111001110110111;
ROM[15240] <= 32'b00001100100000111000001110010011;
ROM[15241] <= 32'b00000000111000111000001110110011;
ROM[15242] <= 32'b00000000000000111000000011100111;
ROM[15243] <= 32'b00000001100000011010001110000011;
ROM[15244] <= 32'b00000000011100010010000000100011;
ROM[15245] <= 32'b00000000010000010000000100010011;
ROM[15246] <= 32'b00000010110000011010001110000011;
ROM[15247] <= 32'b00000000011100010010000000100011;
ROM[15248] <= 32'b00000000010000010000000100010011;
ROM[15249] <= 32'b11111111110000010000000100010011;
ROM[15250] <= 32'b00000000000000010010001110000011;
ROM[15251] <= 32'b11111111110000010000000100010011;
ROM[15252] <= 32'b00000000000000010010010000000011;
ROM[15253] <= 32'b00000000011101000010010010110011;
ROM[15254] <= 32'b00000000100000111010010100110011;
ROM[15255] <= 32'b00000000101001001000001110110011;
ROM[15256] <= 32'b00000000000100111000001110010011;
ROM[15257] <= 32'b00000000000100111111001110010011;
ROM[15258] <= 32'b00000000011100010010000000100011;
ROM[15259] <= 32'b00000000010000010000000100010011;
ROM[15260] <= 32'b11111111110000010000000100010011;
ROM[15261] <= 32'b00000000000000010010001110000011;
ROM[15262] <= 32'b00000000000000111000101001100011;
ROM[15263] <= 32'b00000000000000001111001110110111;
ROM[15264] <= 32'b00000110110000111000001110010011;
ROM[15265] <= 32'b00000000111000111000001110110011;
ROM[15266] <= 32'b00000000000000111000000011100111;
ROM[15267] <= 32'b00000001100000011010001110000011;
ROM[15268] <= 32'b00000000011100010010000000100011;
ROM[15269] <= 32'b00000000010000010000000100010011;
ROM[15270] <= 32'b00000011010000011010001110000011;
ROM[15271] <= 32'b00000000011100010010000000100011;
ROM[15272] <= 32'b00000000010000010000000100010011;
ROM[15273] <= 32'b11111111110000010000000100010011;
ROM[15274] <= 32'b00000000000000010010001110000011;
ROM[15275] <= 32'b11111111110000010000000100010011;
ROM[15276] <= 32'b00000000000000010010010000000011;
ROM[15277] <= 32'b00000000011101000010010010110011;
ROM[15278] <= 32'b00000000100000111010010100110011;
ROM[15279] <= 32'b00000000101001001000001110110011;
ROM[15280] <= 32'b00000000000100111000001110010011;
ROM[15281] <= 32'b00000000000100111111001110010011;
ROM[15282] <= 32'b00000000011100010010000000100011;
ROM[15283] <= 32'b00000000010000010000000100010011;
ROM[15284] <= 32'b11111111110000010000000100010011;
ROM[15285] <= 32'b00000000000000010010001110000011;
ROM[15286] <= 32'b00000000000000111000101001100011;
ROM[15287] <= 32'b00000000000000001111001110110111;
ROM[15288] <= 32'b00000001000000111000001110010011;
ROM[15289] <= 32'b00000000111000111000001110110011;
ROM[15290] <= 32'b00000000000000111000000011100111;
ROM[15291] <= 32'b00000001100000011010001110000011;
ROM[15292] <= 32'b00000000011100010010000000100011;
ROM[15293] <= 32'b00000000010000010000000100010011;
ROM[15294] <= 32'b00000011000000011010001110000011;
ROM[15295] <= 32'b00000000011100010010000000100011;
ROM[15296] <= 32'b00000000010000010000000100010011;
ROM[15297] <= 32'b11111111110000010000000100010011;
ROM[15298] <= 32'b00000000000000010010001110000011;
ROM[15299] <= 32'b11111111110000010000000100010011;
ROM[15300] <= 32'b00000000000000010010010000000011;
ROM[15301] <= 32'b00000000011101000010010010110011;
ROM[15302] <= 32'b00000000100000111010010100110011;
ROM[15303] <= 32'b00000000101001001000001110110011;
ROM[15304] <= 32'b00000000000100111000001110010011;
ROM[15305] <= 32'b00000000000100111111001110010011;
ROM[15306] <= 32'b00000000011100010010000000100011;
ROM[15307] <= 32'b00000000010000010000000100010011;
ROM[15308] <= 32'b11111111110000010000000100010011;
ROM[15309] <= 32'b00000000000000010010001110000011;
ROM[15310] <= 32'b00000000000000111000101001100011;
ROM[15311] <= 32'b00000000000000001111001110110111;
ROM[15312] <= 32'b11111011010000111000001110010011;
ROM[15313] <= 32'b00000000111000111000001110110011;
ROM[15314] <= 32'b00000000000000111000000011100111;
ROM[15315] <= 32'b00000001000000011010001110000011;
ROM[15316] <= 32'b00000000011100010010000000100011;
ROM[15317] <= 32'b00000000010000010000000100010011;
ROM[15318] <= 32'b00000000000000001111001110110111;
ROM[15319] <= 32'b11111010010000111000001110010011;
ROM[15320] <= 32'b00000000111000111000001110110011;
ROM[15321] <= 32'b00000000011100010010000000100011;
ROM[15322] <= 32'b00000000010000010000000100010011;
ROM[15323] <= 32'b00000000001100010010000000100011;
ROM[15324] <= 32'b00000000010000010000000100010011;
ROM[15325] <= 32'b00000000010000010010000000100011;
ROM[15326] <= 32'b00000000010000010000000100010011;
ROM[15327] <= 32'b00000000010100010010000000100011;
ROM[15328] <= 32'b00000000010000010000000100010011;
ROM[15329] <= 32'b00000000011000010010000000100011;
ROM[15330] <= 32'b00000000010000010000000100010011;
ROM[15331] <= 32'b00000001010000000000001110010011;
ROM[15332] <= 32'b00000000010000111000001110010011;
ROM[15333] <= 32'b01000000011100010000001110110011;
ROM[15334] <= 32'b00000000011100000000001000110011;
ROM[15335] <= 32'b00000000001000000000000110110011;
ROM[15336] <= 32'b01111100100100000111000011101111;
ROM[15337] <= 32'b11111111110000010000000100010011;
ROM[15338] <= 32'b00000000000000010010001110000011;
ROM[15339] <= 32'b00000000011101100010000000100011;
ROM[15340] <= 32'b00000101110000000000000011101111;
ROM[15341] <= 32'b00000000000000001111001110110111;
ROM[15342] <= 32'b00000000000000111000001110010011;
ROM[15343] <= 32'b00000000111000111000001110110011;
ROM[15344] <= 32'b00000000011100010010000000100011;
ROM[15345] <= 32'b00000000010000010000000100010011;
ROM[15346] <= 32'b00000000001100010010000000100011;
ROM[15347] <= 32'b00000000010000010000000100010011;
ROM[15348] <= 32'b00000000010000010010000000100011;
ROM[15349] <= 32'b00000000010000010000000100010011;
ROM[15350] <= 32'b00000000010100010010000000100011;
ROM[15351] <= 32'b00000000010000010000000100010011;
ROM[15352] <= 32'b00000000011000010010000000100011;
ROM[15353] <= 32'b00000000010000010000000100010011;
ROM[15354] <= 32'b00000001010000000000001110010011;
ROM[15355] <= 32'b00000000000000111000001110010011;
ROM[15356] <= 32'b01000000011100010000001110110011;
ROM[15357] <= 32'b00000000011100000000001000110011;
ROM[15358] <= 32'b00000000001000000000000110110011;
ROM[15359] <= 32'b01001010100100010100000011101111;
ROM[15360] <= 32'b11111111110000010000000100010011;
ROM[15361] <= 32'b00000000000000010010001110000011;
ROM[15362] <= 32'b00000000011101100010000000100011;
ROM[15363] <= 32'b00000101110000000000000011101111;
ROM[15364] <= 32'b00000000000000001111001110110111;
ROM[15365] <= 32'b00000101110000111000001110010011;
ROM[15366] <= 32'b00000000111000111000001110110011;
ROM[15367] <= 32'b00000000011100010010000000100011;
ROM[15368] <= 32'b00000000010000010000000100010011;
ROM[15369] <= 32'b00000000001100010010000000100011;
ROM[15370] <= 32'b00000000010000010000000100010011;
ROM[15371] <= 32'b00000000010000010010000000100011;
ROM[15372] <= 32'b00000000010000010000000100010011;
ROM[15373] <= 32'b00000000010100010010000000100011;
ROM[15374] <= 32'b00000000010000010000000100010011;
ROM[15375] <= 32'b00000000011000010010000000100011;
ROM[15376] <= 32'b00000000010000010000000100010011;
ROM[15377] <= 32'b00000001010000000000001110010011;
ROM[15378] <= 32'b00000000000000111000001110010011;
ROM[15379] <= 32'b01000000011100010000001110110011;
ROM[15380] <= 32'b00000000011100000000001000110011;
ROM[15381] <= 32'b00000000001000000000000110110011;
ROM[15382] <= 32'b11100100010111110101000011101111;
ROM[15383] <= 32'b11111111110000010000000100010011;
ROM[15384] <= 32'b00000000000000010010001110000011;
ROM[15385] <= 32'b00000000011101100010000000100011;
ROM[15386] <= 32'b00000101110000000000000011101111;
ROM[15387] <= 32'b00000000000000001111001110110111;
ROM[15388] <= 32'b00001011100000111000001110010011;
ROM[15389] <= 32'b00000000111000111000001110110011;
ROM[15390] <= 32'b00000000011100010010000000100011;
ROM[15391] <= 32'b00000000010000010000000100010011;
ROM[15392] <= 32'b00000000001100010010000000100011;
ROM[15393] <= 32'b00000000010000010000000100010011;
ROM[15394] <= 32'b00000000010000010010000000100011;
ROM[15395] <= 32'b00000000010000010000000100010011;
ROM[15396] <= 32'b00000000010100010010000000100011;
ROM[15397] <= 32'b00000000010000010000000100010011;
ROM[15398] <= 32'b00000000011000010010000000100011;
ROM[15399] <= 32'b00000000010000010000000100010011;
ROM[15400] <= 32'b00000001010000000000001110010011;
ROM[15401] <= 32'b00000000000000111000001110010011;
ROM[15402] <= 32'b01000000011100010000001110110011;
ROM[15403] <= 32'b00000000011100000000001000110011;
ROM[15404] <= 32'b00000000001000000000000110110011;
ROM[15405] <= 32'b01100101110000001100000011101111;
ROM[15406] <= 32'b11111111110000010000000100010011;
ROM[15407] <= 32'b00000000000000010010001110000011;
ROM[15408] <= 32'b00000000011101100010000000100011;
ROM[15409] <= 32'b00000101110000000000000011101111;
ROM[15410] <= 32'b00000000000000001111001110110111;
ROM[15411] <= 32'b00010001010000111000001110010011;
ROM[15412] <= 32'b00000000111000111000001110110011;
ROM[15413] <= 32'b00000000011100010010000000100011;
ROM[15414] <= 32'b00000000010000010000000100010011;
ROM[15415] <= 32'b00000000001100010010000000100011;
ROM[15416] <= 32'b00000000010000010000000100010011;
ROM[15417] <= 32'b00000000010000010010000000100011;
ROM[15418] <= 32'b00000000010000010000000100010011;
ROM[15419] <= 32'b00000000010100010010000000100011;
ROM[15420] <= 32'b00000000010000010000000100010011;
ROM[15421] <= 32'b00000000011000010010000000100011;
ROM[15422] <= 32'b00000000010000010000000100010011;
ROM[15423] <= 32'b00000001010000000000001110010011;
ROM[15424] <= 32'b00000000000000111000001110010011;
ROM[15425] <= 32'b01000000011100010000001110110011;
ROM[15426] <= 32'b00000000011100000000001000110011;
ROM[15427] <= 32'b00000000001000000000000110110011;
ROM[15428] <= 32'b11010111000011110011000011101111;
ROM[15429] <= 32'b11111111110000010000000100010011;
ROM[15430] <= 32'b00000000000000010010001110000011;
ROM[15431] <= 32'b00000000011101100010000000100011;
ROM[15432] <= 32'b00000001110000000000000011101111;
ROM[15433] <= 32'b00000000001000000000001110010011;
ROM[15434] <= 32'b00000000011100010010000000100011;
ROM[15435] <= 32'b00000000010000010000000100010011;
ROM[15436] <= 32'b11111111110000010000000100010011;
ROM[15437] <= 32'b00000000000000010010001110000011;
ROM[15438] <= 32'b00000000011100011010000000100011;
ROM[15439] <= 32'b00001100110000000000000011101111;
ROM[15440] <= 32'b00000000000000001111001110110111;
ROM[15441] <= 32'b00011000110000111000001110010011;
ROM[15442] <= 32'b00000000111000111000001110110011;
ROM[15443] <= 32'b00000000011100010010000000100011;
ROM[15444] <= 32'b00000000010000010000000100010011;
ROM[15445] <= 32'b00000000001100010010000000100011;
ROM[15446] <= 32'b00000000010000010000000100010011;
ROM[15447] <= 32'b00000000010000010010000000100011;
ROM[15448] <= 32'b00000000010000010000000100010011;
ROM[15449] <= 32'b00000000010100010010000000100011;
ROM[15450] <= 32'b00000000010000010000000100010011;
ROM[15451] <= 32'b00000000011000010010000000100011;
ROM[15452] <= 32'b00000000010000010000000100010011;
ROM[15453] <= 32'b00000001010000000000001110010011;
ROM[15454] <= 32'b00000000000000111000001110010011;
ROM[15455] <= 32'b01000000011100010000001110110011;
ROM[15456] <= 32'b00000000011100000000001000110011;
ROM[15457] <= 32'b00000000001000000000000110110011;
ROM[15458] <= 32'b01001100000100001110000011101111;
ROM[15459] <= 32'b11111111110000010000000100010011;
ROM[15460] <= 32'b00000000000000010010001110000011;
ROM[15461] <= 32'b00000000011101100010000000100011;
ROM[15462] <= 32'b00000000000000000000001110010011;
ROM[15463] <= 32'b00000000011100010010000000100011;
ROM[15464] <= 32'b00000000010000010000000100010011;
ROM[15465] <= 32'b00000000000000000000001110010011;
ROM[15466] <= 32'b00000000011100010010000000100011;
ROM[15467] <= 32'b00000000010000010000000100010011;
ROM[15468] <= 32'b00000000000000001111001110110111;
ROM[15469] <= 32'b00011111110000111000001110010011;
ROM[15470] <= 32'b00000000111000111000001110110011;
ROM[15471] <= 32'b00000000011100010010000000100011;
ROM[15472] <= 32'b00000000010000010000000100010011;
ROM[15473] <= 32'b00000000001100010010000000100011;
ROM[15474] <= 32'b00000000010000010000000100010011;
ROM[15475] <= 32'b00000000010000010010000000100011;
ROM[15476] <= 32'b00000000010000010000000100010011;
ROM[15477] <= 32'b00000000010100010010000000100011;
ROM[15478] <= 32'b00000000010000010000000100010011;
ROM[15479] <= 32'b00000000011000010010000000100011;
ROM[15480] <= 32'b00000000010000010000000100010011;
ROM[15481] <= 32'b00000001010000000000001110010011;
ROM[15482] <= 32'b00000000100000111000001110010011;
ROM[15483] <= 32'b01000000011100010000001110110011;
ROM[15484] <= 32'b00000000011100000000001000110011;
ROM[15485] <= 32'b00000000001000000000000110110011;
ROM[15486] <= 32'b00100000100100000110000011101111;
ROM[15487] <= 32'b11111111110000010000000100010011;
ROM[15488] <= 32'b00000000000000010010001110000011;
ROM[15489] <= 32'b00000000011101100010000000100011;
ROM[15490] <= 32'b01100001110100000000000011101111;
ROM[15491] <= 32'b00000000011000000000001110010011;
ROM[15492] <= 32'b00000000011100010010000000100011;
ROM[15493] <= 32'b00000000010000010000000100010011;
ROM[15494] <= 32'b00000000000000001111001110110111;
ROM[15495] <= 32'b00100110010000111000001110010011;
ROM[15496] <= 32'b00000000111000111000001110110011;
ROM[15497] <= 32'b00000000011100010010000000100011;
ROM[15498] <= 32'b00000000010000010000000100010011;
ROM[15499] <= 32'b00000000001100010010000000100011;
ROM[15500] <= 32'b00000000010000010000000100010011;
ROM[15501] <= 32'b00000000010000010010000000100011;
ROM[15502] <= 32'b00000000010000010000000100010011;
ROM[15503] <= 32'b00000000010100010010000000100011;
ROM[15504] <= 32'b00000000010000010000000100010011;
ROM[15505] <= 32'b00000000011000010010000000100011;
ROM[15506] <= 32'b00000000010000010000000100010011;
ROM[15507] <= 32'b00000001010000000000001110010011;
ROM[15508] <= 32'b00000000010000111000001110010011;
ROM[15509] <= 32'b01000000011100010000001110110011;
ROM[15510] <= 32'b00000000011100000000001000110011;
ROM[15511] <= 32'b00000000001000000000000110110011;
ROM[15512] <= 32'b01001101110000011010000011101111;
ROM[15513] <= 32'b00000010000000000000001110010011;
ROM[15514] <= 32'b00000000011100010010000000100011;
ROM[15515] <= 32'b00000000010000010000000100010011;
ROM[15516] <= 32'b00000000000000001111001110110111;
ROM[15517] <= 32'b00101011110000111000001110010011;
ROM[15518] <= 32'b00000000111000111000001110110011;
ROM[15519] <= 32'b00000000011100010010000000100011;
ROM[15520] <= 32'b00000000010000010000000100010011;
ROM[15521] <= 32'b00000000001100010010000000100011;
ROM[15522] <= 32'b00000000010000010000000100010011;
ROM[15523] <= 32'b00000000010000010010000000100011;
ROM[15524] <= 32'b00000000010000010000000100010011;
ROM[15525] <= 32'b00000000010100010010000000100011;
ROM[15526] <= 32'b00000000010000010000000100010011;
ROM[15527] <= 32'b00000000011000010010000000100011;
ROM[15528] <= 32'b00000000010000010000000100010011;
ROM[15529] <= 32'b00000001010000000000001110010011;
ROM[15530] <= 32'b00000000100000111000001110010011;
ROM[15531] <= 32'b01000000011100010000001110110011;
ROM[15532] <= 32'b00000000011100000000001000110011;
ROM[15533] <= 32'b00000000001000000000000110110011;
ROM[15534] <= 32'b00001111010100011010000011101111;
ROM[15535] <= 32'b00000110011000000000001110010011;
ROM[15536] <= 32'b00000000011100010010000000100011;
ROM[15537] <= 32'b00000000010000010000000100010011;
ROM[15538] <= 32'b00000000000000001111001110110111;
ROM[15539] <= 32'b00110001010000111000001110010011;
ROM[15540] <= 32'b00000000111000111000001110110011;
ROM[15541] <= 32'b00000000011100010010000000100011;
ROM[15542] <= 32'b00000000010000010000000100010011;
ROM[15543] <= 32'b00000000001100010010000000100011;
ROM[15544] <= 32'b00000000010000010000000100010011;
ROM[15545] <= 32'b00000000010000010010000000100011;
ROM[15546] <= 32'b00000000010000010000000100010011;
ROM[15547] <= 32'b00000000010100010010000000100011;
ROM[15548] <= 32'b00000000010000010000000100010011;
ROM[15549] <= 32'b00000000011000010010000000100011;
ROM[15550] <= 32'b00000000010000010000000100010011;
ROM[15551] <= 32'b00000001010000000000001110010011;
ROM[15552] <= 32'b00000000100000111000001110010011;
ROM[15553] <= 32'b01000000011100010000001110110011;
ROM[15554] <= 32'b00000000011100000000001000110011;
ROM[15555] <= 32'b00000000001000000000000110110011;
ROM[15556] <= 32'b00001001110100011010000011101111;
ROM[15557] <= 32'b00000110100100000000001110010011;
ROM[15558] <= 32'b00000000011100010010000000100011;
ROM[15559] <= 32'b00000000010000010000000100010011;
ROM[15560] <= 32'b00000000000000001111001110110111;
ROM[15561] <= 32'b00110110110000111000001110010011;
ROM[15562] <= 32'b00000000111000111000001110110011;
ROM[15563] <= 32'b00000000011100010010000000100011;
ROM[15564] <= 32'b00000000010000010000000100010011;
ROM[15565] <= 32'b00000000001100010010000000100011;
ROM[15566] <= 32'b00000000010000010000000100010011;
ROM[15567] <= 32'b00000000010000010010000000100011;
ROM[15568] <= 32'b00000000010000010000000100010011;
ROM[15569] <= 32'b00000000010100010010000000100011;
ROM[15570] <= 32'b00000000010000010000000100010011;
ROM[15571] <= 32'b00000000011000010010000000100011;
ROM[15572] <= 32'b00000000010000010000000100010011;
ROM[15573] <= 32'b00000001010000000000001110010011;
ROM[15574] <= 32'b00000000100000111000001110010011;
ROM[15575] <= 32'b01000000011100010000001110110011;
ROM[15576] <= 32'b00000000011100000000001000110011;
ROM[15577] <= 32'b00000000001000000000000110110011;
ROM[15578] <= 32'b00000100010100011010000011101111;
ROM[15579] <= 32'b00000110001000000000001110010011;
ROM[15580] <= 32'b00000000011100010010000000100011;
ROM[15581] <= 32'b00000000010000010000000100010011;
ROM[15582] <= 32'b00000000000000001111001110110111;
ROM[15583] <= 32'b00111100010000111000001110010011;
ROM[15584] <= 32'b00000000111000111000001110110011;
ROM[15585] <= 32'b00000000011100010010000000100011;
ROM[15586] <= 32'b00000000010000010000000100010011;
ROM[15587] <= 32'b00000000001100010010000000100011;
ROM[15588] <= 32'b00000000010000010000000100010011;
ROM[15589] <= 32'b00000000010000010010000000100011;
ROM[15590] <= 32'b00000000010000010000000100010011;
ROM[15591] <= 32'b00000000010100010010000000100011;
ROM[15592] <= 32'b00000000010000010000000100010011;
ROM[15593] <= 32'b00000000011000010010000000100011;
ROM[15594] <= 32'b00000000010000010000000100010011;
ROM[15595] <= 32'b00000001010000000000001110010011;
ROM[15596] <= 32'b00000000100000111000001110010011;
ROM[15597] <= 32'b01000000011100010000001110110011;
ROM[15598] <= 32'b00000000011100000000001000110011;
ROM[15599] <= 32'b00000000001000000000000110110011;
ROM[15600] <= 32'b01111110110000011010000011101111;
ROM[15601] <= 32'b00000110111100000000001110010011;
ROM[15602] <= 32'b00000000011100010010000000100011;
ROM[15603] <= 32'b00000000010000010000000100010011;
ROM[15604] <= 32'b00000000000000001111001110110111;
ROM[15605] <= 32'b01000001110000111000001110010011;
ROM[15606] <= 32'b00000000111000111000001110110011;
ROM[15607] <= 32'b00000000011100010010000000100011;
ROM[15608] <= 32'b00000000010000010000000100010011;
ROM[15609] <= 32'b00000000001100010010000000100011;
ROM[15610] <= 32'b00000000010000010000000100010011;
ROM[15611] <= 32'b00000000010000010010000000100011;
ROM[15612] <= 32'b00000000010000010000000100010011;
ROM[15613] <= 32'b00000000010100010010000000100011;
ROM[15614] <= 32'b00000000010000010000000100010011;
ROM[15615] <= 32'b00000000011000010010000000100011;
ROM[15616] <= 32'b00000000010000010000000100010011;
ROM[15617] <= 32'b00000001010000000000001110010011;
ROM[15618] <= 32'b00000000100000111000001110010011;
ROM[15619] <= 32'b01000000011100010000001110110011;
ROM[15620] <= 32'b00000000011100000000001000110011;
ROM[15621] <= 32'b00000000001000000000000110110011;
ROM[15622] <= 32'b01111001010000011010000011101111;
ROM[15623] <= 32'b00000010000000000000001110010011;
ROM[15624] <= 32'b00000000011100010010000000100011;
ROM[15625] <= 32'b00000000010000010000000100010011;
ROM[15626] <= 32'b00000000000000001111001110110111;
ROM[15627] <= 32'b01000111010000111000001110010011;
ROM[15628] <= 32'b00000000111000111000001110110011;
ROM[15629] <= 32'b00000000011100010010000000100011;
ROM[15630] <= 32'b00000000010000010000000100010011;
ROM[15631] <= 32'b00000000001100010010000000100011;
ROM[15632] <= 32'b00000000010000010000000100010011;
ROM[15633] <= 32'b00000000010000010010000000100011;
ROM[15634] <= 32'b00000000010000010000000100010011;
ROM[15635] <= 32'b00000000010100010010000000100011;
ROM[15636] <= 32'b00000000010000010000000100010011;
ROM[15637] <= 32'b00000000011000010010000000100011;
ROM[15638] <= 32'b00000000010000010000000100010011;
ROM[15639] <= 32'b00000001010000000000001110010011;
ROM[15640] <= 32'b00000000100000111000001110010011;
ROM[15641] <= 32'b01000000011100010000001110110011;
ROM[15642] <= 32'b00000000011100000000001000110011;
ROM[15643] <= 32'b00000000001000000000000110110011;
ROM[15644] <= 32'b01110011110000011010000011101111;
ROM[15645] <= 32'b00000000000000001111001110110111;
ROM[15646] <= 32'b01001100000000111000001110010011;
ROM[15647] <= 32'b00000000111000111000001110110011;
ROM[15648] <= 32'b00000000011100010010000000100011;
ROM[15649] <= 32'b00000000010000010000000100010011;
ROM[15650] <= 32'b00000000001100010010000000100011;
ROM[15651] <= 32'b00000000010000010000000100010011;
ROM[15652] <= 32'b00000000010000010010000000100011;
ROM[15653] <= 32'b00000000010000010000000100010011;
ROM[15654] <= 32'b00000000010100010010000000100011;
ROM[15655] <= 32'b00000000010000010000000100010011;
ROM[15656] <= 32'b00000000011000010010000000100011;
ROM[15657] <= 32'b00000000010000010000000100010011;
ROM[15658] <= 32'b00000001010000000000001110010011;
ROM[15659] <= 32'b00000000010000111000001110010011;
ROM[15660] <= 32'b01000000011100010000001110110011;
ROM[15661] <= 32'b00000000011100000000001000110011;
ROM[15662] <= 32'b00000000001000000000000110110011;
ROM[15663] <= 32'b00101010110100000111000011101111;
ROM[15664] <= 32'b11111111110000010000000100010011;
ROM[15665] <= 32'b00000000000000010010001110000011;
ROM[15666] <= 32'b00000000011101100010000000100011;
ROM[15667] <= 32'b00000000101100000000001110010011;
ROM[15668] <= 32'b00000000011100010010000000100011;
ROM[15669] <= 32'b00000000010000010000000100010011;
ROM[15670] <= 32'b00000000000000001111001110110111;
ROM[15671] <= 32'b01010010010000111000001110010011;
ROM[15672] <= 32'b00000000111000111000001110110011;
ROM[15673] <= 32'b00000000011100010010000000100011;
ROM[15674] <= 32'b00000000010000010000000100010011;
ROM[15675] <= 32'b00000000001100010010000000100011;
ROM[15676] <= 32'b00000000010000010000000100010011;
ROM[15677] <= 32'b00000000010000010010000000100011;
ROM[15678] <= 32'b00000000010000010000000100010011;
ROM[15679] <= 32'b00000000010100010010000000100011;
ROM[15680] <= 32'b00000000010000010000000100010011;
ROM[15681] <= 32'b00000000011000010010000000100011;
ROM[15682] <= 32'b00000000010000010000000100010011;
ROM[15683] <= 32'b00000001010000000000001110010011;
ROM[15684] <= 32'b00000000010000111000001110010011;
ROM[15685] <= 32'b01000000011100010000001110110011;
ROM[15686] <= 32'b00000000011100000000001000110011;
ROM[15687] <= 32'b00000000001000000000000110110011;
ROM[15688] <= 32'b00100001110000011010000011101111;
ROM[15689] <= 32'b00000010000000000000001110010011;
ROM[15690] <= 32'b00000000011100010010000000100011;
ROM[15691] <= 32'b00000000010000010000000100010011;
ROM[15692] <= 32'b00000000000000001111001110110111;
ROM[15693] <= 32'b01010111110000111000001110010011;
ROM[15694] <= 32'b00000000111000111000001110110011;
ROM[15695] <= 32'b00000000011100010010000000100011;
ROM[15696] <= 32'b00000000010000010000000100010011;
ROM[15697] <= 32'b00000000001100010010000000100011;
ROM[15698] <= 32'b00000000010000010000000100010011;
ROM[15699] <= 32'b00000000010000010010000000100011;
ROM[15700] <= 32'b00000000010000010000000100010011;
ROM[15701] <= 32'b00000000010100010010000000100011;
ROM[15702] <= 32'b00000000010000010000000100010011;
ROM[15703] <= 32'b00000000011000010010000000100011;
ROM[15704] <= 32'b00000000010000010000000100010011;
ROM[15705] <= 32'b00000001010000000000001110010011;
ROM[15706] <= 32'b00000000100000111000001110010011;
ROM[15707] <= 32'b01000000011100010000001110110011;
ROM[15708] <= 32'b00000000011100000000001000110011;
ROM[15709] <= 32'b00000000001000000000000110110011;
ROM[15710] <= 32'b01100011010000011010000011101111;
ROM[15711] <= 32'b00000111001100000000001110010011;
ROM[15712] <= 32'b00000000011100010010000000100011;
ROM[15713] <= 32'b00000000010000010000000100010011;
ROM[15714] <= 32'b00000000000000001111001110110111;
ROM[15715] <= 32'b01011101010000111000001110010011;
ROM[15716] <= 32'b00000000111000111000001110110011;
ROM[15717] <= 32'b00000000011100010010000000100011;
ROM[15718] <= 32'b00000000010000010000000100010011;
ROM[15719] <= 32'b00000000001100010010000000100011;
ROM[15720] <= 32'b00000000010000010000000100010011;
ROM[15721] <= 32'b00000000010000010010000000100011;
ROM[15722] <= 32'b00000000010000010000000100010011;
ROM[15723] <= 32'b00000000010100010010000000100011;
ROM[15724] <= 32'b00000000010000010000000100010011;
ROM[15725] <= 32'b00000000011000010010000000100011;
ROM[15726] <= 32'b00000000010000010000000100010011;
ROM[15727] <= 32'b00000001010000000000001110010011;
ROM[15728] <= 32'b00000000100000111000001110010011;
ROM[15729] <= 32'b01000000011100010000001110110011;
ROM[15730] <= 32'b00000000011100000000001000110011;
ROM[15731] <= 32'b00000000001000000000000110110011;
ROM[15732] <= 32'b01011101110000011010000011101111;
ROM[15733] <= 32'b00000110111000000000001110010011;
ROM[15734] <= 32'b00000000011100010010000000100011;
ROM[15735] <= 32'b00000000010000010000000100010011;
ROM[15736] <= 32'b00000000000000001111001110110111;
ROM[15737] <= 32'b01100010110000111000001110010011;
ROM[15738] <= 32'b00000000111000111000001110110011;
ROM[15739] <= 32'b00000000011100010010000000100011;
ROM[15740] <= 32'b00000000010000010000000100010011;
ROM[15741] <= 32'b00000000001100010010000000100011;
ROM[15742] <= 32'b00000000010000010000000100010011;
ROM[15743] <= 32'b00000000010000010010000000100011;
ROM[15744] <= 32'b00000000010000010000000100010011;
ROM[15745] <= 32'b00000000010100010010000000100011;
ROM[15746] <= 32'b00000000010000010000000100010011;
ROM[15747] <= 32'b00000000011000010010000000100011;
ROM[15748] <= 32'b00000000010000010000000100010011;
ROM[15749] <= 32'b00000001010000000000001110010011;
ROM[15750] <= 32'b00000000100000111000001110010011;
ROM[15751] <= 32'b01000000011100010000001110110011;
ROM[15752] <= 32'b00000000011100000000001000110011;
ROM[15753] <= 32'b00000000001000000000000110110011;
ROM[15754] <= 32'b01011000010000011010000011101111;
ROM[15755] <= 32'b00000110000100000000001110010011;
ROM[15756] <= 32'b00000000011100010010000000100011;
ROM[15757] <= 32'b00000000010000010000000100010011;
ROM[15758] <= 32'b00000000000000001111001110110111;
ROM[15759] <= 32'b01101000010000111000001110010011;
ROM[15760] <= 32'b00000000111000111000001110110011;
ROM[15761] <= 32'b00000000011100010010000000100011;
ROM[15762] <= 32'b00000000010000010000000100010011;
ROM[15763] <= 32'b00000000001100010010000000100011;
ROM[15764] <= 32'b00000000010000010000000100010011;
ROM[15765] <= 32'b00000000010000010010000000100011;
ROM[15766] <= 32'b00000000010000010000000100010011;
ROM[15767] <= 32'b00000000010100010010000000100011;
ROM[15768] <= 32'b00000000010000010000000100010011;
ROM[15769] <= 32'b00000000011000010010000000100011;
ROM[15770] <= 32'b00000000010000010000000100010011;
ROM[15771] <= 32'b00000001010000000000001110010011;
ROM[15772] <= 32'b00000000100000111000001110010011;
ROM[15773] <= 32'b01000000011100010000001110110011;
ROM[15774] <= 32'b00000000011100000000001000110011;
ROM[15775] <= 32'b00000000001000000000000110110011;
ROM[15776] <= 32'b01010010110000011010000011101111;
ROM[15777] <= 32'b00000110101100000000001110010011;
ROM[15778] <= 32'b00000000011100010010000000100011;
ROM[15779] <= 32'b00000000010000010000000100010011;
ROM[15780] <= 32'b00000000000000001111001110110111;
ROM[15781] <= 32'b01101101110000111000001110010011;
ROM[15782] <= 32'b00000000111000111000001110110011;
ROM[15783] <= 32'b00000000011100010010000000100011;
ROM[15784] <= 32'b00000000010000010000000100010011;
ROM[15785] <= 32'b00000000001100010010000000100011;
ROM[15786] <= 32'b00000000010000010000000100010011;
ROM[15787] <= 32'b00000000010000010010000000100011;
ROM[15788] <= 32'b00000000010000010000000100010011;
ROM[15789] <= 32'b00000000010100010010000000100011;
ROM[15790] <= 32'b00000000010000010000000100010011;
ROM[15791] <= 32'b00000000011000010010000000100011;
ROM[15792] <= 32'b00000000010000010000000100010011;
ROM[15793] <= 32'b00000001010000000000001110010011;
ROM[15794] <= 32'b00000000100000111000001110010011;
ROM[15795] <= 32'b01000000011100010000001110110011;
ROM[15796] <= 32'b00000000011100000000001000110011;
ROM[15797] <= 32'b00000000001000000000000110110011;
ROM[15798] <= 32'b01001101010000011010000011101111;
ROM[15799] <= 32'b00000110010100000000001110010011;
ROM[15800] <= 32'b00000000011100010010000000100011;
ROM[15801] <= 32'b00000000010000010000000100010011;
ROM[15802] <= 32'b00000000000000001111001110110111;
ROM[15803] <= 32'b01110011010000111000001110010011;
ROM[15804] <= 32'b00000000111000111000001110110011;
ROM[15805] <= 32'b00000000011100010010000000100011;
ROM[15806] <= 32'b00000000010000010000000100010011;
ROM[15807] <= 32'b00000000001100010010000000100011;
ROM[15808] <= 32'b00000000010000010000000100010011;
ROM[15809] <= 32'b00000000010000010010000000100011;
ROM[15810] <= 32'b00000000010000010000000100010011;
ROM[15811] <= 32'b00000000010100010010000000100011;
ROM[15812] <= 32'b00000000010000010000000100010011;
ROM[15813] <= 32'b00000000011000010010000000100011;
ROM[15814] <= 32'b00000000010000010000000100010011;
ROM[15815] <= 32'b00000001010000000000001110010011;
ROM[15816] <= 32'b00000000100000111000001110010011;
ROM[15817] <= 32'b01000000011100010000001110110011;
ROM[15818] <= 32'b00000000011100000000001000110011;
ROM[15819] <= 32'b00000000001000000000000110110011;
ROM[15820] <= 32'b01000111110000011010000011101111;
ROM[15821] <= 32'b00000110011100000000001110010011;
ROM[15822] <= 32'b00000000011100010010000000100011;
ROM[15823] <= 32'b00000000010000010000000100010011;
ROM[15824] <= 32'b00000000000000001111001110110111;
ROM[15825] <= 32'b01111000110000111000001110010011;
ROM[15826] <= 32'b00000000111000111000001110110011;
ROM[15827] <= 32'b00000000011100010010000000100011;
ROM[15828] <= 32'b00000000010000010000000100010011;
ROM[15829] <= 32'b00000000001100010010000000100011;
ROM[15830] <= 32'b00000000010000010000000100010011;
ROM[15831] <= 32'b00000000010000010010000000100011;
ROM[15832] <= 32'b00000000010000010000000100010011;
ROM[15833] <= 32'b00000000010100010010000000100011;
ROM[15834] <= 32'b00000000010000010000000100010011;
ROM[15835] <= 32'b00000000011000010010000000100011;
ROM[15836] <= 32'b00000000010000010000000100010011;
ROM[15837] <= 32'b00000001010000000000001110010011;
ROM[15838] <= 32'b00000000100000111000001110010011;
ROM[15839] <= 32'b01000000011100010000001110110011;
ROM[15840] <= 32'b00000000011100000000001000110011;
ROM[15841] <= 32'b00000000001000000000000110110011;
ROM[15842] <= 32'b01000010010000011010000011101111;
ROM[15843] <= 32'b00000110000100000000001110010011;
ROM[15844] <= 32'b00000000011100010010000000100011;
ROM[15845] <= 32'b00000000010000010000000100010011;
ROM[15846] <= 32'b00000000000000001111001110110111;
ROM[15847] <= 32'b01111110010000111000001110010011;
ROM[15848] <= 32'b00000000111000111000001110110011;
ROM[15849] <= 32'b00000000011100010010000000100011;
ROM[15850] <= 32'b00000000010000010000000100010011;
ROM[15851] <= 32'b00000000001100010010000000100011;
ROM[15852] <= 32'b00000000010000010000000100010011;
ROM[15853] <= 32'b00000000010000010010000000100011;
ROM[15854] <= 32'b00000000010000010000000100010011;
ROM[15855] <= 32'b00000000010100010010000000100011;
ROM[15856] <= 32'b00000000010000010000000100010011;
ROM[15857] <= 32'b00000000011000010010000000100011;
ROM[15858] <= 32'b00000000010000010000000100010011;
ROM[15859] <= 32'b00000001010000000000001110010011;
ROM[15860] <= 32'b00000000100000111000001110010011;
ROM[15861] <= 32'b01000000011100010000001110110011;
ROM[15862] <= 32'b00000000011100000000001000110011;
ROM[15863] <= 32'b00000000001000000000000110110011;
ROM[15864] <= 32'b00111100110000011010000011101111;
ROM[15865] <= 32'b00000110110100000000001110010011;
ROM[15866] <= 32'b00000000011100010010000000100011;
ROM[15867] <= 32'b00000000010000010000000100010011;
ROM[15868] <= 32'b00000000000000010000001110110111;
ROM[15869] <= 32'b10000011110000111000001110010011;
ROM[15870] <= 32'b00000000111000111000001110110011;
ROM[15871] <= 32'b00000000011100010010000000100011;
ROM[15872] <= 32'b00000000010000010000000100010011;
ROM[15873] <= 32'b00000000001100010010000000100011;
ROM[15874] <= 32'b00000000010000010000000100010011;
ROM[15875] <= 32'b00000000010000010010000000100011;
ROM[15876] <= 32'b00000000010000010000000100010011;
ROM[15877] <= 32'b00000000010100010010000000100011;
ROM[15878] <= 32'b00000000010000010000000100010011;
ROM[15879] <= 32'b00000000011000010010000000100011;
ROM[15880] <= 32'b00000000010000010000000100010011;
ROM[15881] <= 32'b00000001010000000000001110010011;
ROM[15882] <= 32'b00000000100000111000001110010011;
ROM[15883] <= 32'b01000000011100010000001110110011;
ROM[15884] <= 32'b00000000011100000000001000110011;
ROM[15885] <= 32'b00000000001000000000000110110011;
ROM[15886] <= 32'b00110111010000011010000011101111;
ROM[15887] <= 32'b00000110010100000000001110010011;
ROM[15888] <= 32'b00000000011100010010000000100011;
ROM[15889] <= 32'b00000000010000010000000100010011;
ROM[15890] <= 32'b00000000000000010000001110110111;
ROM[15891] <= 32'b10001001010000111000001110010011;
ROM[15892] <= 32'b00000000111000111000001110110011;
ROM[15893] <= 32'b00000000011100010010000000100011;
ROM[15894] <= 32'b00000000010000010000000100010011;
ROM[15895] <= 32'b00000000001100010010000000100011;
ROM[15896] <= 32'b00000000010000010000000100010011;
ROM[15897] <= 32'b00000000010000010010000000100011;
ROM[15898] <= 32'b00000000010000010000000100010011;
ROM[15899] <= 32'b00000000010100010010000000100011;
ROM[15900] <= 32'b00000000010000010000000100010011;
ROM[15901] <= 32'b00000000011000010010000000100011;
ROM[15902] <= 32'b00000000010000010000000100010011;
ROM[15903] <= 32'b00000001010000000000001110010011;
ROM[15904] <= 32'b00000000100000111000001110010011;
ROM[15905] <= 32'b01000000011100010000001110110011;
ROM[15906] <= 32'b00000000011100000000001000110011;
ROM[15907] <= 32'b00000000001000000000000110110011;
ROM[15908] <= 32'b00110001110000011010000011101111;
ROM[15909] <= 32'b00000010000000000000001110010011;
ROM[15910] <= 32'b00000000011100010010000000100011;
ROM[15911] <= 32'b00000000010000010000000100010011;
ROM[15912] <= 32'b00000000000000010000001110110111;
ROM[15913] <= 32'b10001110110000111000001110010011;
ROM[15914] <= 32'b00000000111000111000001110110011;
ROM[15915] <= 32'b00000000011100010010000000100011;
ROM[15916] <= 32'b00000000010000010000000100010011;
ROM[15917] <= 32'b00000000001100010010000000100011;
ROM[15918] <= 32'b00000000010000010000000100010011;
ROM[15919] <= 32'b00000000010000010010000000100011;
ROM[15920] <= 32'b00000000010000010000000100010011;
ROM[15921] <= 32'b00000000010100010010000000100011;
ROM[15922] <= 32'b00000000010000010000000100010011;
ROM[15923] <= 32'b00000000011000010010000000100011;
ROM[15924] <= 32'b00000000010000010000000100010011;
ROM[15925] <= 32'b00000001010000000000001110010011;
ROM[15926] <= 32'b00000000100000111000001110010011;
ROM[15927] <= 32'b01000000011100010000001110110011;
ROM[15928] <= 32'b00000000011100000000001000110011;
ROM[15929] <= 32'b00000000001000000000000110110011;
ROM[15930] <= 32'b00101100010000011010000011101111;
ROM[15931] <= 32'b00000000000000010000001110110111;
ROM[15932] <= 32'b10010011100000111000001110010011;
ROM[15933] <= 32'b00000000111000111000001110110011;
ROM[15934] <= 32'b00000000011100010010000000100011;
ROM[15935] <= 32'b00000000010000010000000100010011;
ROM[15936] <= 32'b00000000001100010010000000100011;
ROM[15937] <= 32'b00000000010000010000000100010011;
ROM[15938] <= 32'b00000000010000010010000000100011;
ROM[15939] <= 32'b00000000010000010000000100010011;
ROM[15940] <= 32'b00000000010100010010000000100011;
ROM[15941] <= 32'b00000000010000010000000100010011;
ROM[15942] <= 32'b00000000011000010010000000100011;
ROM[15943] <= 32'b00000000010000010000000100010011;
ROM[15944] <= 32'b00000001010000000000001110010011;
ROM[15945] <= 32'b00000000010000111000001110010011;
ROM[15946] <= 32'b01000000011100010000001110110011;
ROM[15947] <= 32'b00000000011100000000001000110011;
ROM[15948] <= 32'b00000000001000000000000110110011;
ROM[15949] <= 32'b01100011010000000111000011101111;
ROM[15950] <= 32'b11111111110000010000000100010011;
ROM[15951] <= 32'b00000000000000010010001110000011;
ROM[15952] <= 32'b00000000011101100010000000100011;
ROM[15953] <= 32'b00000000011100000000001110010011;
ROM[15954] <= 32'b00000000011100010010000000100011;
ROM[15955] <= 32'b00000000010000010000000100010011;
ROM[15956] <= 32'b00000000000000010000001110110111;
ROM[15957] <= 32'b10011001110000111000001110010011;
ROM[15958] <= 32'b00000000111000111000001110110011;
ROM[15959] <= 32'b00000000011100010010000000100011;
ROM[15960] <= 32'b00000000010000010000000100010011;
ROM[15961] <= 32'b00000000001100010010000000100011;
ROM[15962] <= 32'b00000000010000010000000100010011;
ROM[15963] <= 32'b00000000010000010010000000100011;
ROM[15964] <= 32'b00000000010000010000000100010011;
ROM[15965] <= 32'b00000000010100010010000000100011;
ROM[15966] <= 32'b00000000010000010000000100010011;
ROM[15967] <= 32'b00000000011000010010000000100011;
ROM[15968] <= 32'b00000000010000010000000100010011;
ROM[15969] <= 32'b00000001010000000000001110010011;
ROM[15970] <= 32'b00000000010000111000001110010011;
ROM[15971] <= 32'b01000000011100010000001110110011;
ROM[15972] <= 32'b00000000011100000000001000110011;
ROM[15973] <= 32'b00000000001000000000000110110011;
ROM[15974] <= 32'b01011010010100011001000011101111;
ROM[15975] <= 32'b00000010000000000000001110010011;
ROM[15976] <= 32'b00000000011100010010000000100011;
ROM[15977] <= 32'b00000000010000010000000100010011;
ROM[15978] <= 32'b00000000000000010000001110110111;
ROM[15979] <= 32'b10011111010000111000001110010011;
ROM[15980] <= 32'b00000000111000111000001110110011;
ROM[15981] <= 32'b00000000011100010010000000100011;
ROM[15982] <= 32'b00000000010000010000000100010011;
ROM[15983] <= 32'b00000000001100010010000000100011;
ROM[15984] <= 32'b00000000010000010000000100010011;
ROM[15985] <= 32'b00000000010000010010000000100011;
ROM[15986] <= 32'b00000000010000010000000100010011;
ROM[15987] <= 32'b00000000010100010010000000100011;
ROM[15988] <= 32'b00000000010000010000000100010011;
ROM[15989] <= 32'b00000000011000010010000000100011;
ROM[15990] <= 32'b00000000010000010000000100010011;
ROM[15991] <= 32'b00000001010000000000001110010011;
ROM[15992] <= 32'b00000000100000111000001110010011;
ROM[15993] <= 32'b01000000011100010000001110110011;
ROM[15994] <= 32'b00000000011100000000001000110011;
ROM[15995] <= 32'b00000000001000000000000110110011;
ROM[15996] <= 32'b00011011110000011010000011101111;
ROM[15997] <= 32'b00000111000100000000001110010011;
ROM[15998] <= 32'b00000000011100010010000000100011;
ROM[15999] <= 32'b00000000010000010000000100010011;
ROM[16000] <= 32'b00000000000000010000001110110111;
ROM[16001] <= 32'b10100100110000111000001110010011;
ROM[16002] <= 32'b00000000111000111000001110110011;
ROM[16003] <= 32'b00000000011100010010000000100011;
ROM[16004] <= 32'b00000000010000010000000100010011;
ROM[16005] <= 32'b00000000001100010010000000100011;
ROM[16006] <= 32'b00000000010000010000000100010011;
ROM[16007] <= 32'b00000000010000010010000000100011;
ROM[16008] <= 32'b00000000010000010000000100010011;
ROM[16009] <= 32'b00000000010100010010000000100011;
ROM[16010] <= 32'b00000000010000010000000100010011;
ROM[16011] <= 32'b00000000011000010010000000100011;
ROM[16012] <= 32'b00000000010000010000000100010011;
ROM[16013] <= 32'b00000001010000000000001110010011;
ROM[16014] <= 32'b00000000100000111000001110010011;
ROM[16015] <= 32'b01000000011100010000001110110011;
ROM[16016] <= 32'b00000000011100000000001000110011;
ROM[16017] <= 32'b00000000001000000000000110110011;
ROM[16018] <= 32'b00010110010000011010000011101111;
ROM[16019] <= 32'b00000111001100000000001110010011;
ROM[16020] <= 32'b00000000011100010010000000100011;
ROM[16021] <= 32'b00000000010000010000000100010011;
ROM[16022] <= 32'b00000000000000010000001110110111;
ROM[16023] <= 32'b10101010010000111000001110010011;
ROM[16024] <= 32'b00000000111000111000001110110011;
ROM[16025] <= 32'b00000000011100010010000000100011;
ROM[16026] <= 32'b00000000010000010000000100010011;
ROM[16027] <= 32'b00000000001100010010000000100011;
ROM[16028] <= 32'b00000000010000010000000100010011;
ROM[16029] <= 32'b00000000010000010010000000100011;
ROM[16030] <= 32'b00000000010000010000000100010011;
ROM[16031] <= 32'b00000000010100010010000000100011;
ROM[16032] <= 32'b00000000010000010000000100010011;
ROM[16033] <= 32'b00000000011000010010000000100011;
ROM[16034] <= 32'b00000000010000010000000100010011;
ROM[16035] <= 32'b00000001010000000000001110010011;
ROM[16036] <= 32'b00000000100000111000001110010011;
ROM[16037] <= 32'b01000000011100010000001110110011;
ROM[16038] <= 32'b00000000011100000000001000110011;
ROM[16039] <= 32'b00000000001000000000000110110011;
ROM[16040] <= 32'b00010000110000011010000011101111;
ROM[16041] <= 32'b00000110111100000000001110010011;
ROM[16042] <= 32'b00000000011100010010000000100011;
ROM[16043] <= 32'b00000000010000010000000100010011;
ROM[16044] <= 32'b00000000000000010000001110110111;
ROM[16045] <= 32'b10101111110000111000001110010011;
ROM[16046] <= 32'b00000000111000111000001110110011;
ROM[16047] <= 32'b00000000011100010010000000100011;
ROM[16048] <= 32'b00000000010000010000000100010011;
ROM[16049] <= 32'b00000000001100010010000000100011;
ROM[16050] <= 32'b00000000010000010000000100010011;
ROM[16051] <= 32'b00000000010000010010000000100011;
ROM[16052] <= 32'b00000000010000010000000100010011;
ROM[16053] <= 32'b00000000010100010010000000100011;
ROM[16054] <= 32'b00000000010000010000000100010011;
ROM[16055] <= 32'b00000000011000010010000000100011;
ROM[16056] <= 32'b00000000010000010000000100010011;
ROM[16057] <= 32'b00000001010000000000001110010011;
ROM[16058] <= 32'b00000000100000111000001110010011;
ROM[16059] <= 32'b01000000011100010000001110110011;
ROM[16060] <= 32'b00000000011100000000001000110011;
ROM[16061] <= 32'b00000000001000000000000110110011;
ROM[16062] <= 32'b00001011010000011010000011101111;
ROM[16063] <= 32'b00000111001000000000001110010011;
ROM[16064] <= 32'b00000000011100010010000000100011;
ROM[16065] <= 32'b00000000010000010000000100010011;
ROM[16066] <= 32'b00000000000000010000001110110111;
ROM[16067] <= 32'b10110101010000111000001110010011;
ROM[16068] <= 32'b00000000111000111000001110110011;
ROM[16069] <= 32'b00000000011100010010000000100011;
ROM[16070] <= 32'b00000000010000010000000100010011;
ROM[16071] <= 32'b00000000001100010010000000100011;
ROM[16072] <= 32'b00000000010000010000000100010011;
ROM[16073] <= 32'b00000000010000010010000000100011;
ROM[16074] <= 32'b00000000010000010000000100010011;
ROM[16075] <= 32'b00000000010100010010000000100011;
ROM[16076] <= 32'b00000000010000010000000100010011;
ROM[16077] <= 32'b00000000011000010010000000100011;
ROM[16078] <= 32'b00000000010000010000000100010011;
ROM[16079] <= 32'b00000001010000000000001110010011;
ROM[16080] <= 32'b00000000100000111000001110010011;
ROM[16081] <= 32'b01000000011100010000001110110011;
ROM[16082] <= 32'b00000000011100000000001000110011;
ROM[16083] <= 32'b00000000001000000000000110110011;
ROM[16084] <= 32'b00000101110000011010000011101111;
ROM[16085] <= 32'b00000111010000000000001110010011;
ROM[16086] <= 32'b00000000011100010010000000100011;
ROM[16087] <= 32'b00000000010000010000000100010011;
ROM[16088] <= 32'b00000000000000010000001110110111;
ROM[16089] <= 32'b10111010110000111000001110010011;
ROM[16090] <= 32'b00000000111000111000001110110011;
ROM[16091] <= 32'b00000000011100010010000000100011;
ROM[16092] <= 32'b00000000010000010000000100010011;
ROM[16093] <= 32'b00000000001100010010000000100011;
ROM[16094] <= 32'b00000000010000010000000100010011;
ROM[16095] <= 32'b00000000010000010010000000100011;
ROM[16096] <= 32'b00000000010000010000000100010011;
ROM[16097] <= 32'b00000000010100010010000000100011;
ROM[16098] <= 32'b00000000010000010000000100010011;
ROM[16099] <= 32'b00000000011000010010000000100011;
ROM[16100] <= 32'b00000000010000010000000100010011;
ROM[16101] <= 32'b00000001010000000000001110010011;
ROM[16102] <= 32'b00000000100000111000001110010011;
ROM[16103] <= 32'b01000000011100010000001110110011;
ROM[16104] <= 32'b00000000011100000000001000110011;
ROM[16105] <= 32'b00000000001000000000000110110011;
ROM[16106] <= 32'b00000000010000011010000011101111;
ROM[16107] <= 32'b00000010000000000000001110010011;
ROM[16108] <= 32'b00000000011100010010000000100011;
ROM[16109] <= 32'b00000000010000010000000100010011;
ROM[16110] <= 32'b00000000000000010000001110110111;
ROM[16111] <= 32'b11000000010000111000001110010011;
ROM[16112] <= 32'b00000000111000111000001110110011;
ROM[16113] <= 32'b00000000011100010010000000100011;
ROM[16114] <= 32'b00000000010000010000000100010011;
ROM[16115] <= 32'b00000000001100010010000000100011;
ROM[16116] <= 32'b00000000010000010000000100010011;
ROM[16117] <= 32'b00000000010000010010000000100011;
ROM[16118] <= 32'b00000000010000010000000100010011;
ROM[16119] <= 32'b00000000010100010010000000100011;
ROM[16120] <= 32'b00000000010000010000000100010011;
ROM[16121] <= 32'b00000000011000010010000000100011;
ROM[16122] <= 32'b00000000010000010000000100010011;
ROM[16123] <= 32'b00000001010000000000001110010011;
ROM[16124] <= 32'b00000000100000111000001110010011;
ROM[16125] <= 32'b01000000011100010000001110110011;
ROM[16126] <= 32'b00000000011100000000001000110011;
ROM[16127] <= 32'b00000000001000000000000110110011;
ROM[16128] <= 32'b01111010110100011001000011101111;
ROM[16129] <= 32'b00000000000000010000001110110111;
ROM[16130] <= 32'b11000101000000111000001110010011;
ROM[16131] <= 32'b00000000111000111000001110110011;
ROM[16132] <= 32'b00000000011100010010000000100011;
ROM[16133] <= 32'b00000000010000010000000100010011;
ROM[16134] <= 32'b00000000001100010010000000100011;
ROM[16135] <= 32'b00000000010000010000000100010011;
ROM[16136] <= 32'b00000000010000010010000000100011;
ROM[16137] <= 32'b00000000010000010000000100010011;
ROM[16138] <= 32'b00000000010100010010000000100011;
ROM[16139] <= 32'b00000000010000010000000100010011;
ROM[16140] <= 32'b00000000011000010010000000100011;
ROM[16141] <= 32'b00000000010000010000000100010011;
ROM[16142] <= 32'b00000001010000000000001110010011;
ROM[16143] <= 32'b00000000010000111000001110010011;
ROM[16144] <= 32'b01000000011100010000001110110011;
ROM[16145] <= 32'b00000000011100000000001000110011;
ROM[16146] <= 32'b00000000001000000000000110110011;
ROM[16147] <= 32'b00110001110000000111000011101111;
ROM[16148] <= 32'b11111111110000010000000100010011;
ROM[16149] <= 32'b00000000000000010010001110000011;
ROM[16150] <= 32'b00000000011101100010000000100011;
ROM[16151] <= 32'b00000000100100000000001110010011;
ROM[16152] <= 32'b00000000011100010010000000100011;
ROM[16153] <= 32'b00000000010000010000000100010011;
ROM[16154] <= 32'b00000000000000010000001110110111;
ROM[16155] <= 32'b11001011010000111000001110010011;
ROM[16156] <= 32'b00000000111000111000001110110011;
ROM[16157] <= 32'b00000000011100010010000000100011;
ROM[16158] <= 32'b00000000010000010000000100010011;
ROM[16159] <= 32'b00000000001100010010000000100011;
ROM[16160] <= 32'b00000000010000010000000100010011;
ROM[16161] <= 32'b00000000010000010010000000100011;
ROM[16162] <= 32'b00000000010000010000000100010011;
ROM[16163] <= 32'b00000000010100010010000000100011;
ROM[16164] <= 32'b00000000010000010000000100010011;
ROM[16165] <= 32'b00000000011000010010000000100011;
ROM[16166] <= 32'b00000000010000010000000100010011;
ROM[16167] <= 32'b00000001010000000000001110010011;
ROM[16168] <= 32'b00000000010000111000001110010011;
ROM[16169] <= 32'b01000000011100010000001110110011;
ROM[16170] <= 32'b00000000011100000000001000110011;
ROM[16171] <= 32'b00000000001000000000000110110011;
ROM[16172] <= 32'b00101000110100011001000011101111;
ROM[16173] <= 32'b00000010000000000000001110010011;
ROM[16174] <= 32'b00000000011100010010000000100011;
ROM[16175] <= 32'b00000000010000010000000100010011;
ROM[16176] <= 32'b00000000000000010000001110110111;
ROM[16177] <= 32'b11010000110000111000001110010011;
ROM[16178] <= 32'b00000000111000111000001110110011;
ROM[16179] <= 32'b00000000011100010010000000100011;
ROM[16180] <= 32'b00000000010000010000000100010011;
ROM[16181] <= 32'b00000000001100010010000000100011;
ROM[16182] <= 32'b00000000010000010000000100010011;
ROM[16183] <= 32'b00000000010000010010000000100011;
ROM[16184] <= 32'b00000000010000010000000100010011;
ROM[16185] <= 32'b00000000010100010010000000100011;
ROM[16186] <= 32'b00000000010000010000000100010011;
ROM[16187] <= 32'b00000000011000010010000000100011;
ROM[16188] <= 32'b00000000010000010000000100010011;
ROM[16189] <= 32'b00000001010000000000001110010011;
ROM[16190] <= 32'b00000000100000111000001110010011;
ROM[16191] <= 32'b01000000011100010000001110110011;
ROM[16192] <= 32'b00000000011100000000001000110011;
ROM[16193] <= 32'b00000000001000000000000110110011;
ROM[16194] <= 32'b01101010010100011001000011101111;
ROM[16195] <= 32'b00000110100000000000001110010011;
ROM[16196] <= 32'b00000000011100010010000000100011;
ROM[16197] <= 32'b00000000010000010000000100010011;
ROM[16198] <= 32'b00000000000000010000001110110111;
ROM[16199] <= 32'b11010110010000111000001110010011;
ROM[16200] <= 32'b00000000111000111000001110110011;
ROM[16201] <= 32'b00000000011100010010000000100011;
ROM[16202] <= 32'b00000000010000010000000100010011;
ROM[16203] <= 32'b00000000001100010010000000100011;
ROM[16204] <= 32'b00000000010000010000000100010011;
ROM[16205] <= 32'b00000000010000010010000000100011;
ROM[16206] <= 32'b00000000010000010000000100010011;
ROM[16207] <= 32'b00000000010100010010000000100011;
ROM[16208] <= 32'b00000000010000010000000100010011;
ROM[16209] <= 32'b00000000011000010010000000100011;
ROM[16210] <= 32'b00000000010000010000000100010011;
ROM[16211] <= 32'b00000001010000000000001110010011;
ROM[16212] <= 32'b00000000100000111000001110010011;
ROM[16213] <= 32'b01000000011100010000001110110011;
ROM[16214] <= 32'b00000000011100000000001000110011;
ROM[16215] <= 32'b00000000001000000000000110110011;
ROM[16216] <= 32'b01100100110100011001000011101111;
ROM[16217] <= 32'b00000110000100000000001110010011;
ROM[16218] <= 32'b00000000011100010010000000100011;
ROM[16219] <= 32'b00000000010000010000000100010011;
ROM[16220] <= 32'b00000000000000010000001110110111;
ROM[16221] <= 32'b11011011110000111000001110010011;
ROM[16222] <= 32'b00000000111000111000001110110011;
ROM[16223] <= 32'b00000000011100010010000000100011;
ROM[16224] <= 32'b00000000010000010000000100010011;
ROM[16225] <= 32'b00000000001100010010000000100011;
ROM[16226] <= 32'b00000000010000010000000100010011;
ROM[16227] <= 32'b00000000010000010010000000100011;
ROM[16228] <= 32'b00000000010000010000000100010011;
ROM[16229] <= 32'b00000000010100010010000000100011;
ROM[16230] <= 32'b00000000010000010000000100010011;
ROM[16231] <= 32'b00000000011000010010000000100011;
ROM[16232] <= 32'b00000000010000010000000100010011;
ROM[16233] <= 32'b00000001010000000000001110010011;
ROM[16234] <= 32'b00000000100000111000001110010011;
ROM[16235] <= 32'b01000000011100010000001110110011;
ROM[16236] <= 32'b00000000011100000000001000110011;
ROM[16237] <= 32'b00000000001000000000000110110011;
ROM[16238] <= 32'b01011111010100011001000011101111;
ROM[16239] <= 32'b00000110111000000000001110010011;
ROM[16240] <= 32'b00000000011100010010000000100011;
ROM[16241] <= 32'b00000000010000010000000100010011;
ROM[16242] <= 32'b00000000000000010000001110110111;
ROM[16243] <= 32'b11100001010000111000001110010011;
ROM[16244] <= 32'b00000000111000111000001110110011;
ROM[16245] <= 32'b00000000011100010010000000100011;
ROM[16246] <= 32'b00000000010000010000000100010011;
ROM[16247] <= 32'b00000000001100010010000000100011;
ROM[16248] <= 32'b00000000010000010000000100010011;
ROM[16249] <= 32'b00000000010000010010000000100011;
ROM[16250] <= 32'b00000000010000010000000100010011;
ROM[16251] <= 32'b00000000010100010010000000100011;
ROM[16252] <= 32'b00000000010000010000000100010011;
ROM[16253] <= 32'b00000000011000010010000000100011;
ROM[16254] <= 32'b00000000010000010000000100010011;
ROM[16255] <= 32'b00000001010000000000001110010011;
ROM[16256] <= 32'b00000000100000111000001110010011;
ROM[16257] <= 32'b01000000011100010000001110110011;
ROM[16258] <= 32'b00000000011100000000001000110011;
ROM[16259] <= 32'b00000000001000000000000110110011;
ROM[16260] <= 32'b01011001110100011001000011101111;
ROM[16261] <= 32'b00000110011100000000001110010011;
ROM[16262] <= 32'b00000000011100010010000000100011;
ROM[16263] <= 32'b00000000010000010000000100010011;
ROM[16264] <= 32'b00000000000000010000001110110111;
ROM[16265] <= 32'b11100110110000111000001110010011;
ROM[16266] <= 32'b00000000111000111000001110110011;
ROM[16267] <= 32'b00000000011100010010000000100011;
ROM[16268] <= 32'b00000000010000010000000100010011;
ROM[16269] <= 32'b00000000001100010010000000100011;
ROM[16270] <= 32'b00000000010000010000000100010011;
ROM[16271] <= 32'b00000000010000010010000000100011;
ROM[16272] <= 32'b00000000010000010000000100010011;
ROM[16273] <= 32'b00000000010100010010000000100011;
ROM[16274] <= 32'b00000000010000010000000100010011;
ROM[16275] <= 32'b00000000011000010010000000100011;
ROM[16276] <= 32'b00000000010000010000000100010011;
ROM[16277] <= 32'b00000001010000000000001110010011;
ROM[16278] <= 32'b00000000100000111000001110010011;
ROM[16279] <= 32'b01000000011100010000001110110011;
ROM[16280] <= 32'b00000000011100000000001000110011;
ROM[16281] <= 32'b00000000001000000000000110110011;
ROM[16282] <= 32'b01010100010100011001000011101111;
ROM[16283] <= 32'b00000110110100000000001110010011;
ROM[16284] <= 32'b00000000011100010010000000100011;
ROM[16285] <= 32'b00000000010000010000000100010011;
ROM[16286] <= 32'b00000000000000010000001110110111;
ROM[16287] <= 32'b11101100010000111000001110010011;
ROM[16288] <= 32'b00000000111000111000001110110011;
ROM[16289] <= 32'b00000000011100010010000000100011;
ROM[16290] <= 32'b00000000010000010000000100010011;
ROM[16291] <= 32'b00000000001100010010000000100011;
ROM[16292] <= 32'b00000000010000010000000100010011;
ROM[16293] <= 32'b00000000010000010010000000100011;
ROM[16294] <= 32'b00000000010000010000000100010011;
ROM[16295] <= 32'b00000000010100010010000000100011;
ROM[16296] <= 32'b00000000010000010000000100010011;
ROM[16297] <= 32'b00000000011000010010000000100011;
ROM[16298] <= 32'b00000000010000010000000100010011;
ROM[16299] <= 32'b00000001010000000000001110010011;
ROM[16300] <= 32'b00000000100000111000001110010011;
ROM[16301] <= 32'b01000000011100010000001110110011;
ROM[16302] <= 32'b00000000011100000000001000110011;
ROM[16303] <= 32'b00000000001000000000000110110011;
ROM[16304] <= 32'b01001110110100011001000011101111;
ROM[16305] <= 32'b00000110000100000000001110010011;
ROM[16306] <= 32'b00000000011100010010000000100011;
ROM[16307] <= 32'b00000000010000010000000100010011;
ROM[16308] <= 32'b00000000000000010000001110110111;
ROM[16309] <= 32'b11110001110000111000001110010011;
ROM[16310] <= 32'b00000000111000111000001110110011;
ROM[16311] <= 32'b00000000011100010010000000100011;
ROM[16312] <= 32'b00000000010000010000000100010011;
ROM[16313] <= 32'b00000000001100010010000000100011;
ROM[16314] <= 32'b00000000010000010000000100010011;
ROM[16315] <= 32'b00000000010000010010000000100011;
ROM[16316] <= 32'b00000000010000010000000100010011;
ROM[16317] <= 32'b00000000010100010010000000100011;
ROM[16318] <= 32'b00000000010000010000000100010011;
ROM[16319] <= 32'b00000000011000010010000000100011;
ROM[16320] <= 32'b00000000010000010000000100010011;
ROM[16321] <= 32'b00000001010000000000001110010011;
ROM[16322] <= 32'b00000000100000111000001110010011;
ROM[16323] <= 32'b01000000011100010000001110110011;
ROM[16324] <= 32'b00000000011100000000001000110011;
ROM[16325] <= 32'b00000000001000000000000110110011;
ROM[16326] <= 32'b01001001010100011001000011101111;
ROM[16327] <= 32'b00000110111000000000001110010011;
ROM[16328] <= 32'b00000000011100010010000000100011;
ROM[16329] <= 32'b00000000010000010000000100010011;
ROM[16330] <= 32'b00000000000000010000001110110111;
ROM[16331] <= 32'b11110111010000111000001110010011;
ROM[16332] <= 32'b00000000111000111000001110110011;
ROM[16333] <= 32'b00000000011100010010000000100011;
ROM[16334] <= 32'b00000000010000010000000100010011;
ROM[16335] <= 32'b00000000001100010010000000100011;
ROM[16336] <= 32'b00000000010000010000000100010011;
ROM[16337] <= 32'b00000000010000010010000000100011;
ROM[16338] <= 32'b00000000010000010000000100010011;
ROM[16339] <= 32'b00000000010100010010000000100011;
ROM[16340] <= 32'b00000000010000010000000100010011;
ROM[16341] <= 32'b00000000011000010010000000100011;
ROM[16342] <= 32'b00000000010000010000000100010011;
ROM[16343] <= 32'b00000001010000000000001110010011;
ROM[16344] <= 32'b00000000100000111000001110010011;
ROM[16345] <= 32'b01000000011100010000001110110011;
ROM[16346] <= 32'b00000000011100000000001000110011;
ROM[16347] <= 32'b00000000001000000000000110110011;
ROM[16348] <= 32'b01000011110100011001000011101111;
ROM[16349] <= 32'b00000010000000000000001110010011;
ROM[16350] <= 32'b00000000011100010010000000100011;
ROM[16351] <= 32'b00000000010000010000000100010011;
ROM[16352] <= 32'b00000000000000010000001110110111;
ROM[16353] <= 32'b11111100110000111000001110010011;
ROM[16354] <= 32'b00000000111000111000001110110011;
ROM[16355] <= 32'b00000000011100010010000000100011;
ROM[16356] <= 32'b00000000010000010000000100010011;
ROM[16357] <= 32'b00000000001100010010000000100011;
ROM[16358] <= 32'b00000000010000010000000100010011;
ROM[16359] <= 32'b00000000010000010010000000100011;
ROM[16360] <= 32'b00000000010000010000000100010011;
ROM[16361] <= 32'b00000000010100010010000000100011;
ROM[16362] <= 32'b00000000010000010000000100010011;
ROM[16363] <= 32'b00000000011000010010000000100011;
ROM[16364] <= 32'b00000000010000010000000100010011;
ROM[16365] <= 32'b00000001010000000000001110010011;
ROM[16366] <= 32'b00000000100000111000001110010011;
ROM[16367] <= 32'b01000000011100010000001110110011;
ROM[16368] <= 32'b00000000011100000000001000110011;
ROM[16369] <= 32'b00000000001000000000000110110011;
ROM[16370] <= 32'b00111110010100011001000011101111;
ROM[16371] <= 32'b00000000000000010000001110110111;
ROM[16372] <= 32'b00000001100000111000001110010011;
ROM[16373] <= 32'b00000000111000111000001110110011;
ROM[16374] <= 32'b00000000011100010010000000100011;
ROM[16375] <= 32'b00000000010000010000000100010011;
ROM[16376] <= 32'b00000000001100010010000000100011;
ROM[16377] <= 32'b00000000010000010000000100010011;
ROM[16378] <= 32'b00000000010000010010000000100011;
ROM[16379] <= 32'b00000000010000010000000100010011;
ROM[16380] <= 32'b00000000010100010010000000100011;
ROM[16381] <= 32'b00000000010000010000000100010011;
ROM[16382] <= 32'b00000000011000010010000000100011;
ROM[16383] <= 32'b00000000010000010000000100010011;
ROM[16384] <= 32'b00000001010000000000001110010011;
ROM[16385] <= 32'b00000000010000111000001110010011;
ROM[16386] <= 32'b01000000011100010000001110110011;
ROM[16387] <= 32'b00000000011100000000001000110011;
ROM[16388] <= 32'b00000000001000000000000110110011;
ROM[16389] <= 32'b01110101010100000110000011101111;
ROM[16390] <= 32'b11111111110000010000000100010011;
ROM[16391] <= 32'b00000000000000010010001110000011;
ROM[16392] <= 32'b00000000011101100010000000100011;
ROM[16393] <= 32'b00000000000000010000001110110111;
ROM[16394] <= 32'b00000111000000111000001110010011;
ROM[16395] <= 32'b00000000111000111000001110110011;
ROM[16396] <= 32'b00000000011100010010000000100011;
ROM[16397] <= 32'b00000000010000010000000100010011;
ROM[16398] <= 32'b00000000001100010010000000100011;
ROM[16399] <= 32'b00000000010000010000000100010011;
ROM[16400] <= 32'b00000000010000010010000000100011;
ROM[16401] <= 32'b00000000010000010000000100010011;
ROM[16402] <= 32'b00000000010100010010000000100011;
ROM[16403] <= 32'b00000000010000010000000100010011;
ROM[16404] <= 32'b00000000011000010010000000100011;
ROM[16405] <= 32'b00000000010000010000000100010011;
ROM[16406] <= 32'b00000001010000000000001110010011;
ROM[16407] <= 32'b00000000000000111000001110010011;
ROM[16408] <= 32'b01000000011100010000001110110011;
ROM[16409] <= 32'b00000000011100000000001000110011;
ROM[16410] <= 32'b00000000001000000000000110110011;
ROM[16411] <= 32'b00101111110000000111000011101111;
ROM[16412] <= 32'b11111111110000010000000100010011;
ROM[16413] <= 32'b00000000000000010010001110000011;
ROM[16414] <= 32'b00000000011101100010000000100011;
ROM[16415] <= 32'b10101111010111111110000011101111;
ROM[16416] <= 32'b00000000000000000000001110010011;
ROM[16417] <= 32'b00000000011100010010000000100011;
ROM[16418] <= 32'b00000000010000010000000100010011;
ROM[16419] <= 32'b00000001010000000000001110010011;
ROM[16420] <= 32'b01000000011100011000001110110011;
ROM[16421] <= 32'b00000000000000111010000010000011;
ROM[16422] <= 32'b11111111110000010000000100010011;
ROM[16423] <= 32'b00000000000000010010001110000011;
ROM[16424] <= 32'b00000000011100100010000000100011;
ROM[16425] <= 32'b00000000010000100000000100010011;
ROM[16426] <= 32'b00000001010000000000001110010011;
ROM[16427] <= 32'b01000000011100011000001110110011;
ROM[16428] <= 32'b00000000010000111010000110000011;
ROM[16429] <= 32'b00000000100000111010001000000011;
ROM[16430] <= 32'b00000000110000111010001010000011;
ROM[16431] <= 32'b00000001000000111010001100000011;
ROM[16432] <= 32'b00000000000000001000000011100111;
ROM[16433] <= 32'b00000010000000000000001110010011;
ROM[16434] <= 32'b00000000011100010010000000100011;
ROM[16435] <= 32'b00000000010000010000000100010011;
ROM[16436] <= 32'b00000000000000010000001110110111;
ROM[16437] <= 32'b00010001110000111000001110010011;
ROM[16438] <= 32'b00000000111000111000001110110011;
ROM[16439] <= 32'b00000000011100010010000000100011;
ROM[16440] <= 32'b00000000010000010000000100010011;
ROM[16441] <= 32'b00000000001100010010000000100011;
ROM[16442] <= 32'b00000000010000010000000100010011;
ROM[16443] <= 32'b00000000010000010010000000100011;
ROM[16444] <= 32'b00000000010000010000000100010011;
ROM[16445] <= 32'b00000000010100010010000000100011;
ROM[16446] <= 32'b00000000010000010000000100010011;
ROM[16447] <= 32'b00000000011000010010000000100011;
ROM[16448] <= 32'b00000000010000010000000100010011;
ROM[16449] <= 32'b00000001010000000000001110010011;
ROM[16450] <= 32'b00000000010000111000001110010011;
ROM[16451] <= 32'b01000000011100010000001110110011;
ROM[16452] <= 32'b00000000011100000000001000110011;
ROM[16453] <= 32'b00000000001000000000000110110011;
ROM[16454] <= 32'b11110110100111101111000011101111;
ROM[16455] <= 32'b11111111110000010000000100010011;
ROM[16456] <= 32'b00000000000000010010001110000011;
ROM[16457] <= 32'b00000100011101101010001000100011;
ROM[16458] <= 32'b00000000000100000000001110010011;
ROM[16459] <= 32'b00000000011100010010000000100011;
ROM[16460] <= 32'b00000000010000010000000100010011;
ROM[16461] <= 32'b00000100010001101010001110000011;
ROM[16462] <= 32'b00000000011100010010000000100011;
ROM[16463] <= 32'b00000000010000010000000100010011;
ROM[16464] <= 32'b00000000000000000000001110010011;
ROM[16465] <= 32'b00000000011100010010000000100011;
ROM[16466] <= 32'b00000000010000010000000100010011;
ROM[16467] <= 32'b11111111110000010000000100010011;
ROM[16468] <= 32'b00000000000000010010001110000011;
ROM[16469] <= 32'b11111111110000010000000100010011;
ROM[16470] <= 32'b00000000000000010010010000000011;
ROM[16471] <= 32'b00000000011101000000001110110011;
ROM[16472] <= 32'b00000000011100010010000000100011;
ROM[16473] <= 32'b00000000010000010000000100010011;
ROM[16474] <= 32'b11111111110000010000000100010011;
ROM[16475] <= 32'b00000000000000010010001110000011;
ROM[16476] <= 32'b00000000000000111000001100010011;
ROM[16477] <= 32'b11111111110000010000000100010011;
ROM[16478] <= 32'b00000000000000010010001110000011;
ROM[16479] <= 32'b00000000110100110000010000110011;
ROM[16480] <= 32'b00000000011101000010000000100011;
ROM[16481] <= 32'b00000000001000000000001110010011;
ROM[16482] <= 32'b00000000011100010010000000100011;
ROM[16483] <= 32'b00000000010000010000000100010011;
ROM[16484] <= 32'b00000100010001101010001110000011;
ROM[16485] <= 32'b00000000011100010010000000100011;
ROM[16486] <= 32'b00000000010000010000000100010011;
ROM[16487] <= 32'b00000000010000000000001110010011;
ROM[16488] <= 32'b00000000011100010010000000100011;
ROM[16489] <= 32'b00000000010000010000000100010011;
ROM[16490] <= 32'b11111111110000010000000100010011;
ROM[16491] <= 32'b00000000000000010010001110000011;
ROM[16492] <= 32'b11111111110000010000000100010011;
ROM[16493] <= 32'b00000000000000010010010000000011;
ROM[16494] <= 32'b00000000011101000000001110110011;
ROM[16495] <= 32'b00000000011100010010000000100011;
ROM[16496] <= 32'b00000000010000010000000100010011;
ROM[16497] <= 32'b11111111110000010000000100010011;
ROM[16498] <= 32'b00000000000000010010001110000011;
ROM[16499] <= 32'b00000000000000111000001100010011;
ROM[16500] <= 32'b11111111110000010000000100010011;
ROM[16501] <= 32'b00000000000000010010001110000011;
ROM[16502] <= 32'b00000000110100110000010000110011;
ROM[16503] <= 32'b00000000011101000010000000100011;
ROM[16504] <= 32'b00000000010000000000001110010011;
ROM[16505] <= 32'b00000000011100010010000000100011;
ROM[16506] <= 32'b00000000010000010000000100010011;
ROM[16507] <= 32'b00000100010001101010001110000011;
ROM[16508] <= 32'b00000000011100010010000000100011;
ROM[16509] <= 32'b00000000010000010000000100010011;
ROM[16510] <= 32'b00000000100000000000001110010011;
ROM[16511] <= 32'b00000000011100010010000000100011;
ROM[16512] <= 32'b00000000010000010000000100010011;
ROM[16513] <= 32'b11111111110000010000000100010011;
ROM[16514] <= 32'b00000000000000010010001110000011;
ROM[16515] <= 32'b11111111110000010000000100010011;
ROM[16516] <= 32'b00000000000000010010010000000011;
ROM[16517] <= 32'b00000000011101000000001110110011;
ROM[16518] <= 32'b00000000011100010010000000100011;
ROM[16519] <= 32'b00000000010000010000000100010011;
ROM[16520] <= 32'b11111111110000010000000100010011;
ROM[16521] <= 32'b00000000000000010010001110000011;
ROM[16522] <= 32'b00000000000000111000001100010011;
ROM[16523] <= 32'b11111111110000010000000100010011;
ROM[16524] <= 32'b00000000000000010010001110000011;
ROM[16525] <= 32'b00000000110100110000010000110011;
ROM[16526] <= 32'b00000000011101000010000000100011;
ROM[16527] <= 32'b00000000100000000000001110010011;
ROM[16528] <= 32'b00000000011100010010000000100011;
ROM[16529] <= 32'b00000000010000010000000100010011;
ROM[16530] <= 32'b00000100010001101010001110000011;
ROM[16531] <= 32'b00000000011100010010000000100011;
ROM[16532] <= 32'b00000000010000010000000100010011;
ROM[16533] <= 32'b00000000110000000000001110010011;
ROM[16534] <= 32'b00000000011100010010000000100011;
ROM[16535] <= 32'b00000000010000010000000100010011;
ROM[16536] <= 32'b11111111110000010000000100010011;
ROM[16537] <= 32'b00000000000000010010001110000011;
ROM[16538] <= 32'b11111111110000010000000100010011;
ROM[16539] <= 32'b00000000000000010010010000000011;
ROM[16540] <= 32'b00000000011101000000001110110011;
ROM[16541] <= 32'b00000000011100010010000000100011;
ROM[16542] <= 32'b00000000010000010000000100010011;
ROM[16543] <= 32'b11111111110000010000000100010011;
ROM[16544] <= 32'b00000000000000010010001110000011;
ROM[16545] <= 32'b00000000000000111000001100010011;
ROM[16546] <= 32'b11111111110000010000000100010011;
ROM[16547] <= 32'b00000000000000010010001110000011;
ROM[16548] <= 32'b00000000110100110000010000110011;
ROM[16549] <= 32'b00000000011101000010000000100011;
ROM[16550] <= 32'b00000001000000000000001110010011;
ROM[16551] <= 32'b00000000011100010010000000100011;
ROM[16552] <= 32'b00000000010000010000000100010011;
ROM[16553] <= 32'b00000100010001101010001110000011;
ROM[16554] <= 32'b00000000011100010010000000100011;
ROM[16555] <= 32'b00000000010000010000000100010011;
ROM[16556] <= 32'b00000001000000000000001110010011;
ROM[16557] <= 32'b00000000011100010010000000100011;
ROM[16558] <= 32'b00000000010000010000000100010011;
ROM[16559] <= 32'b11111111110000010000000100010011;
ROM[16560] <= 32'b00000000000000010010001110000011;
ROM[16561] <= 32'b11111111110000010000000100010011;
ROM[16562] <= 32'b00000000000000010010010000000011;
ROM[16563] <= 32'b00000000011101000000001110110011;
ROM[16564] <= 32'b00000000011100010010000000100011;
ROM[16565] <= 32'b00000000010000010000000100010011;
ROM[16566] <= 32'b11111111110000010000000100010011;
ROM[16567] <= 32'b00000000000000010010001110000011;
ROM[16568] <= 32'b00000000000000111000001100010011;
ROM[16569] <= 32'b11111111110000010000000100010011;
ROM[16570] <= 32'b00000000000000010010001110000011;
ROM[16571] <= 32'b00000000110100110000010000110011;
ROM[16572] <= 32'b00000000011101000010000000100011;
ROM[16573] <= 32'b00000010000000000000001110010011;
ROM[16574] <= 32'b00000000011100010010000000100011;
ROM[16575] <= 32'b00000000010000010000000100010011;
ROM[16576] <= 32'b00000100010001101010001110000011;
ROM[16577] <= 32'b00000000011100010010000000100011;
ROM[16578] <= 32'b00000000010000010000000100010011;
ROM[16579] <= 32'b00000001010000000000001110010011;
ROM[16580] <= 32'b00000000011100010010000000100011;
ROM[16581] <= 32'b00000000010000010000000100010011;
ROM[16582] <= 32'b11111111110000010000000100010011;
ROM[16583] <= 32'b00000000000000010010001110000011;
ROM[16584] <= 32'b11111111110000010000000100010011;
ROM[16585] <= 32'b00000000000000010010010000000011;
ROM[16586] <= 32'b00000000011101000000001110110011;
ROM[16587] <= 32'b00000000011100010010000000100011;
ROM[16588] <= 32'b00000000010000010000000100010011;
ROM[16589] <= 32'b11111111110000010000000100010011;
ROM[16590] <= 32'b00000000000000010010001110000011;
ROM[16591] <= 32'b00000000000000111000001100010011;
ROM[16592] <= 32'b11111111110000010000000100010011;
ROM[16593] <= 32'b00000000000000010010001110000011;
ROM[16594] <= 32'b00000000110100110000010000110011;
ROM[16595] <= 32'b00000000011101000010000000100011;
ROM[16596] <= 32'b00000100000000000000001110010011;
ROM[16597] <= 32'b00000000011100010010000000100011;
ROM[16598] <= 32'b00000000010000010000000100010011;
ROM[16599] <= 32'b00000100010001101010001110000011;
ROM[16600] <= 32'b00000000011100010010000000100011;
ROM[16601] <= 32'b00000000010000010000000100010011;
ROM[16602] <= 32'b00000001100000000000001110010011;
ROM[16603] <= 32'b00000000011100010010000000100011;
ROM[16604] <= 32'b00000000010000010000000100010011;
ROM[16605] <= 32'b11111111110000010000000100010011;
ROM[16606] <= 32'b00000000000000010010001110000011;
ROM[16607] <= 32'b11111111110000010000000100010011;
ROM[16608] <= 32'b00000000000000010010010000000011;
ROM[16609] <= 32'b00000000011101000000001110110011;
ROM[16610] <= 32'b00000000011100010010000000100011;
ROM[16611] <= 32'b00000000010000010000000100010011;
ROM[16612] <= 32'b11111111110000010000000100010011;
ROM[16613] <= 32'b00000000000000010010001110000011;
ROM[16614] <= 32'b00000000000000111000001100010011;
ROM[16615] <= 32'b11111111110000010000000100010011;
ROM[16616] <= 32'b00000000000000010010001110000011;
ROM[16617] <= 32'b00000000110100110000010000110011;
ROM[16618] <= 32'b00000000011101000010000000100011;
ROM[16619] <= 32'b00001000000000000000001110010011;
ROM[16620] <= 32'b00000000011100010010000000100011;
ROM[16621] <= 32'b00000000010000010000000100010011;
ROM[16622] <= 32'b00000100010001101010001110000011;
ROM[16623] <= 32'b00000000011100010010000000100011;
ROM[16624] <= 32'b00000000010000010000000100010011;
ROM[16625] <= 32'b00000001110000000000001110010011;
ROM[16626] <= 32'b00000000011100010010000000100011;
ROM[16627] <= 32'b00000000010000010000000100010011;
ROM[16628] <= 32'b11111111110000010000000100010011;
ROM[16629] <= 32'b00000000000000010010001110000011;
ROM[16630] <= 32'b11111111110000010000000100010011;
ROM[16631] <= 32'b00000000000000010010010000000011;
ROM[16632] <= 32'b00000000011101000000001110110011;
ROM[16633] <= 32'b00000000011100010010000000100011;
ROM[16634] <= 32'b00000000010000010000000100010011;
ROM[16635] <= 32'b11111111110000010000000100010011;
ROM[16636] <= 32'b00000000000000010010001110000011;
ROM[16637] <= 32'b00000000000000111000001100010011;
ROM[16638] <= 32'b11111111110000010000000100010011;
ROM[16639] <= 32'b00000000000000010010001110000011;
ROM[16640] <= 32'b00000000110100110000010000110011;
ROM[16641] <= 32'b00000000011101000010000000100011;
ROM[16642] <= 32'b00010000000000000000001110010011;
ROM[16643] <= 32'b00000000011100010010000000100011;
ROM[16644] <= 32'b00000000010000010000000100010011;
ROM[16645] <= 32'b00000100010001101010001110000011;
ROM[16646] <= 32'b00000000011100010010000000100011;
ROM[16647] <= 32'b00000000010000010000000100010011;
ROM[16648] <= 32'b00000010000000000000001110010011;
ROM[16649] <= 32'b00000000011100010010000000100011;
ROM[16650] <= 32'b00000000010000010000000100010011;
ROM[16651] <= 32'b11111111110000010000000100010011;
ROM[16652] <= 32'b00000000000000010010001110000011;
ROM[16653] <= 32'b11111111110000010000000100010011;
ROM[16654] <= 32'b00000000000000010010010000000011;
ROM[16655] <= 32'b00000000011101000000001110110011;
ROM[16656] <= 32'b00000000011100010010000000100011;
ROM[16657] <= 32'b00000000010000010000000100010011;
ROM[16658] <= 32'b11111111110000010000000100010011;
ROM[16659] <= 32'b00000000000000010010001110000011;
ROM[16660] <= 32'b00000000000000111000001100010011;
ROM[16661] <= 32'b11111111110000010000000100010011;
ROM[16662] <= 32'b00000000000000010010001110000011;
ROM[16663] <= 32'b00000000110100110000010000110011;
ROM[16664] <= 32'b00000000011101000010000000100011;
ROM[16665] <= 32'b00100000000000000000001110010011;
ROM[16666] <= 32'b00000000011100010010000000100011;
ROM[16667] <= 32'b00000000010000010000000100010011;
ROM[16668] <= 32'b00000100010001101010001110000011;
ROM[16669] <= 32'b00000000011100010010000000100011;
ROM[16670] <= 32'b00000000010000010000000100010011;
ROM[16671] <= 32'b00000010010000000000001110010011;
ROM[16672] <= 32'b00000000011100010010000000100011;
ROM[16673] <= 32'b00000000010000010000000100010011;
ROM[16674] <= 32'b11111111110000010000000100010011;
ROM[16675] <= 32'b00000000000000010010001110000011;
ROM[16676] <= 32'b11111111110000010000000100010011;
ROM[16677] <= 32'b00000000000000010010010000000011;
ROM[16678] <= 32'b00000000011101000000001110110011;
ROM[16679] <= 32'b00000000011100010010000000100011;
ROM[16680] <= 32'b00000000010000010000000100010011;
ROM[16681] <= 32'b11111111110000010000000100010011;
ROM[16682] <= 32'b00000000000000010010001110000011;
ROM[16683] <= 32'b00000000000000111000001100010011;
ROM[16684] <= 32'b11111111110000010000000100010011;
ROM[16685] <= 32'b00000000000000010010001110000011;
ROM[16686] <= 32'b00000000110100110000010000110011;
ROM[16687] <= 32'b00000000011101000010000000100011;
ROM[16688] <= 32'b01000000000000000000001110010011;
ROM[16689] <= 32'b00000000011100010010000000100011;
ROM[16690] <= 32'b00000000010000010000000100010011;
ROM[16691] <= 32'b00000100010001101010001110000011;
ROM[16692] <= 32'b00000000011100010010000000100011;
ROM[16693] <= 32'b00000000010000010000000100010011;
ROM[16694] <= 32'b00000010100000000000001110010011;
ROM[16695] <= 32'b00000000011100010010000000100011;
ROM[16696] <= 32'b00000000010000010000000100010011;
ROM[16697] <= 32'b11111111110000010000000100010011;
ROM[16698] <= 32'b00000000000000010010001110000011;
ROM[16699] <= 32'b11111111110000010000000100010011;
ROM[16700] <= 32'b00000000000000010010010000000011;
ROM[16701] <= 32'b00000000011101000000001110110011;
ROM[16702] <= 32'b00000000011100010010000000100011;
ROM[16703] <= 32'b00000000010000010000000100010011;
ROM[16704] <= 32'b11111111110000010000000100010011;
ROM[16705] <= 32'b00000000000000010010001110000011;
ROM[16706] <= 32'b00000000000000111000001100010011;
ROM[16707] <= 32'b11111111110000010000000100010011;
ROM[16708] <= 32'b00000000000000010010001110000011;
ROM[16709] <= 32'b00000000110100110000010000110011;
ROM[16710] <= 32'b00000000011101000010000000100011;
ROM[16711] <= 32'b00000000000000000001001110110111;
ROM[16712] <= 32'b10000000000000111000001110010011;
ROM[16713] <= 32'b00000000011100010010000000100011;
ROM[16714] <= 32'b00000000010000010000000100010011;
ROM[16715] <= 32'b00000100010001101010001110000011;
ROM[16716] <= 32'b00000000011100010010000000100011;
ROM[16717] <= 32'b00000000010000010000000100010011;
ROM[16718] <= 32'b00000010110000000000001110010011;
ROM[16719] <= 32'b00000000011100010010000000100011;
ROM[16720] <= 32'b00000000010000010000000100010011;
ROM[16721] <= 32'b11111111110000010000000100010011;
ROM[16722] <= 32'b00000000000000010010001110000011;
ROM[16723] <= 32'b11111111110000010000000100010011;
ROM[16724] <= 32'b00000000000000010010010000000011;
ROM[16725] <= 32'b00000000011101000000001110110011;
ROM[16726] <= 32'b00000000011100010010000000100011;
ROM[16727] <= 32'b00000000010000010000000100010011;
ROM[16728] <= 32'b11111111110000010000000100010011;
ROM[16729] <= 32'b00000000000000010010001110000011;
ROM[16730] <= 32'b00000000000000111000001100010011;
ROM[16731] <= 32'b11111111110000010000000100010011;
ROM[16732] <= 32'b00000000000000010010001110000011;
ROM[16733] <= 32'b00000000110100110000010000110011;
ROM[16734] <= 32'b00000000011101000010000000100011;
ROM[16735] <= 32'b00000000000000000001001110110111;
ROM[16736] <= 32'b00000000000000111000001110010011;
ROM[16737] <= 32'b00000000011100010010000000100011;
ROM[16738] <= 32'b00000000010000010000000100010011;
ROM[16739] <= 32'b00000100010001101010001110000011;
ROM[16740] <= 32'b00000000011100010010000000100011;
ROM[16741] <= 32'b00000000010000010000000100010011;
ROM[16742] <= 32'b00000011000000000000001110010011;
ROM[16743] <= 32'b00000000011100010010000000100011;
ROM[16744] <= 32'b00000000010000010000000100010011;
ROM[16745] <= 32'b11111111110000010000000100010011;
ROM[16746] <= 32'b00000000000000010010001110000011;
ROM[16747] <= 32'b11111111110000010000000100010011;
ROM[16748] <= 32'b00000000000000010010010000000011;
ROM[16749] <= 32'b00000000011101000000001110110011;
ROM[16750] <= 32'b00000000011100010010000000100011;
ROM[16751] <= 32'b00000000010000010000000100010011;
ROM[16752] <= 32'b11111111110000010000000100010011;
ROM[16753] <= 32'b00000000000000010010001110000011;
ROM[16754] <= 32'b00000000000000111000001100010011;
ROM[16755] <= 32'b11111111110000010000000100010011;
ROM[16756] <= 32'b00000000000000010010001110000011;
ROM[16757] <= 32'b00000000110100110000010000110011;
ROM[16758] <= 32'b00000000011101000010000000100011;
ROM[16759] <= 32'b00000000000000000010001110110111;
ROM[16760] <= 32'b00000000000000111000001110010011;
ROM[16761] <= 32'b00000000011100010010000000100011;
ROM[16762] <= 32'b00000000010000010000000100010011;
ROM[16763] <= 32'b00000100010001101010001110000011;
ROM[16764] <= 32'b00000000011100010010000000100011;
ROM[16765] <= 32'b00000000010000010000000100010011;
ROM[16766] <= 32'b00000011010000000000001110010011;
ROM[16767] <= 32'b00000000011100010010000000100011;
ROM[16768] <= 32'b00000000010000010000000100010011;
ROM[16769] <= 32'b11111111110000010000000100010011;
ROM[16770] <= 32'b00000000000000010010001110000011;
ROM[16771] <= 32'b11111111110000010000000100010011;
ROM[16772] <= 32'b00000000000000010010010000000011;
ROM[16773] <= 32'b00000000011101000000001110110011;
ROM[16774] <= 32'b00000000011100010010000000100011;
ROM[16775] <= 32'b00000000010000010000000100010011;
ROM[16776] <= 32'b11111111110000010000000100010011;
ROM[16777] <= 32'b00000000000000010010001110000011;
ROM[16778] <= 32'b00000000000000111000001100010011;
ROM[16779] <= 32'b11111111110000010000000100010011;
ROM[16780] <= 32'b00000000000000010010001110000011;
ROM[16781] <= 32'b00000000110100110000010000110011;
ROM[16782] <= 32'b00000000011101000010000000100011;
ROM[16783] <= 32'b00000000000000000100001110110111;
ROM[16784] <= 32'b00000000000000111000001110010011;
ROM[16785] <= 32'b00000000011100010010000000100011;
ROM[16786] <= 32'b00000000010000010000000100010011;
ROM[16787] <= 32'b00000100010001101010001110000011;
ROM[16788] <= 32'b00000000011100010010000000100011;
ROM[16789] <= 32'b00000000010000010000000100010011;
ROM[16790] <= 32'b00000011100000000000001110010011;
ROM[16791] <= 32'b00000000011100010010000000100011;
ROM[16792] <= 32'b00000000010000010000000100010011;
ROM[16793] <= 32'b11111111110000010000000100010011;
ROM[16794] <= 32'b00000000000000010010001110000011;
ROM[16795] <= 32'b11111111110000010000000100010011;
ROM[16796] <= 32'b00000000000000010010010000000011;
ROM[16797] <= 32'b00000000011101000000001110110011;
ROM[16798] <= 32'b00000000011100010010000000100011;
ROM[16799] <= 32'b00000000010000010000000100010011;
ROM[16800] <= 32'b11111111110000010000000100010011;
ROM[16801] <= 32'b00000000000000010010001110000011;
ROM[16802] <= 32'b00000000000000111000001100010011;
ROM[16803] <= 32'b11111111110000010000000100010011;
ROM[16804] <= 32'b00000000000000010010001110000011;
ROM[16805] <= 32'b00000000110100110000010000110011;
ROM[16806] <= 32'b00000000011101000010000000100011;
ROM[16807] <= 32'b00000000000000000100001110110111;
ROM[16808] <= 32'b00000000000000111000001110010011;
ROM[16809] <= 32'b00000000011100010010000000100011;
ROM[16810] <= 32'b00000000010000010000000100010011;
ROM[16811] <= 32'b00000000000000000100001110110111;
ROM[16812] <= 32'b00000000000000111000001110010011;
ROM[16813] <= 32'b00000000011100010010000000100011;
ROM[16814] <= 32'b00000000010000010000000100010011;
ROM[16815] <= 32'b11111111110000010000000100010011;
ROM[16816] <= 32'b00000000000000010010001110000011;
ROM[16817] <= 32'b11111111110000010000000100010011;
ROM[16818] <= 32'b00000000000000010010010000000011;
ROM[16819] <= 32'b00000000011101000000001110110011;
ROM[16820] <= 32'b00000000011100010010000000100011;
ROM[16821] <= 32'b00000000010000010000000100010011;
ROM[16822] <= 32'b00000100010001101010001110000011;
ROM[16823] <= 32'b00000000011100010010000000100011;
ROM[16824] <= 32'b00000000010000010000000100010011;
ROM[16825] <= 32'b00000011110000000000001110010011;
ROM[16826] <= 32'b00000000011100010010000000100011;
ROM[16827] <= 32'b00000000010000010000000100010011;
ROM[16828] <= 32'b11111111110000010000000100010011;
ROM[16829] <= 32'b00000000000000010010001110000011;
ROM[16830] <= 32'b11111111110000010000000100010011;
ROM[16831] <= 32'b00000000000000010010010000000011;
ROM[16832] <= 32'b00000000011101000000001110110011;
ROM[16833] <= 32'b00000000011100010010000000100011;
ROM[16834] <= 32'b00000000010000010000000100010011;
ROM[16835] <= 32'b11111111110000010000000100010011;
ROM[16836] <= 32'b00000000000000010010001110000011;
ROM[16837] <= 32'b00000000000000111000001100010011;
ROM[16838] <= 32'b11111111110000010000000100010011;
ROM[16839] <= 32'b00000000000000010010001110000011;
ROM[16840] <= 32'b00000000110100110000010000110011;
ROM[16841] <= 32'b00000000011101000010000000100011;
ROM[16842] <= 32'b00000100010001101010001110000011;
ROM[16843] <= 32'b00000000011100010010000000100011;
ROM[16844] <= 32'b00000000010000010000000100010011;
ROM[16845] <= 32'b00000011110000000000001110010011;
ROM[16846] <= 32'b00000000011100010010000000100011;
ROM[16847] <= 32'b00000000010000010000000100010011;
ROM[16848] <= 32'b11111111110000010000000100010011;
ROM[16849] <= 32'b00000000000000010010001110000011;
ROM[16850] <= 32'b11111111110000010000000100010011;
ROM[16851] <= 32'b00000000000000010010010000000011;
ROM[16852] <= 32'b00000000011101000000001110110011;
ROM[16853] <= 32'b00000000011100010010000000100011;
ROM[16854] <= 32'b00000000010000010000000100010011;
ROM[16855] <= 32'b11111111110000010000000100010011;
ROM[16856] <= 32'b00000000000000010010001110000011;
ROM[16857] <= 32'b00000000000000111000001100010011;
ROM[16858] <= 32'b00000000110100110000010000110011;
ROM[16859] <= 32'b00000000000001000010001110000011;
ROM[16860] <= 32'b00000000011100010010000000100011;
ROM[16861] <= 32'b00000000010000010000000100010011;
ROM[16862] <= 32'b00000100010001101010001110000011;
ROM[16863] <= 32'b00000000011100010010000000100011;
ROM[16864] <= 32'b00000000010000010000000100010011;
ROM[16865] <= 32'b00000011110000000000001110010011;
ROM[16866] <= 32'b00000000011100010010000000100011;
ROM[16867] <= 32'b00000000010000010000000100010011;
ROM[16868] <= 32'b11111111110000010000000100010011;
ROM[16869] <= 32'b00000000000000010010001110000011;
ROM[16870] <= 32'b11111111110000010000000100010011;
ROM[16871] <= 32'b00000000000000010010010000000011;
ROM[16872] <= 32'b00000000011101000000001110110011;
ROM[16873] <= 32'b00000000011100010010000000100011;
ROM[16874] <= 32'b00000000010000010000000100010011;
ROM[16875] <= 32'b11111111110000010000000100010011;
ROM[16876] <= 32'b00000000000000010010001110000011;
ROM[16877] <= 32'b00000000000000111000001100010011;
ROM[16878] <= 32'b00000000110100110000010000110011;
ROM[16879] <= 32'b00000000000001000010001110000011;
ROM[16880] <= 32'b00000000011100010010000000100011;
ROM[16881] <= 32'b00000000010000010000000100010011;
ROM[16882] <= 32'b11111111110000010000000100010011;
ROM[16883] <= 32'b00000000000000010010001110000011;
ROM[16884] <= 32'b11111111110000010000000100010011;
ROM[16885] <= 32'b00000000000000010010010000000011;
ROM[16886] <= 32'b00000000011101000000001110110011;
ROM[16887] <= 32'b00000000011100010010000000100011;
ROM[16888] <= 32'b00000000010000010000000100010011;
ROM[16889] <= 32'b00000100010001101010001110000011;
ROM[16890] <= 32'b00000000011100010010000000100011;
ROM[16891] <= 32'b00000000010000010000000100010011;
ROM[16892] <= 32'b00000100000000000000001110010011;
ROM[16893] <= 32'b00000000011100010010000000100011;
ROM[16894] <= 32'b00000000010000010000000100010011;
ROM[16895] <= 32'b11111111110000010000000100010011;
ROM[16896] <= 32'b00000000000000010010001110000011;
ROM[16897] <= 32'b11111111110000010000000100010011;
ROM[16898] <= 32'b00000000000000010010010000000011;
ROM[16899] <= 32'b00000000011101000000001110110011;
ROM[16900] <= 32'b00000000011100010010000000100011;
ROM[16901] <= 32'b00000000010000010000000100010011;
ROM[16902] <= 32'b11111111110000010000000100010011;
ROM[16903] <= 32'b00000000000000010010001110000011;
ROM[16904] <= 32'b00000000000000111000001100010011;
ROM[16905] <= 32'b11111111110000010000000100010011;
ROM[16906] <= 32'b00000000000000010010001110000011;
ROM[16907] <= 32'b00000000110100110000010000110011;
ROM[16908] <= 32'b00000000011101000010000000100011;
ROM[16909] <= 32'b00000100010001101010001110000011;
ROM[16910] <= 32'b00000000011100010010000000100011;
ROM[16911] <= 32'b00000000010000010000000100010011;
ROM[16912] <= 32'b00000100000000000000001110010011;
ROM[16913] <= 32'b00000000011100010010000000100011;
ROM[16914] <= 32'b00000000010000010000000100010011;
ROM[16915] <= 32'b11111111110000010000000100010011;
ROM[16916] <= 32'b00000000000000010010001110000011;
ROM[16917] <= 32'b11111111110000010000000100010011;
ROM[16918] <= 32'b00000000000000010010010000000011;
ROM[16919] <= 32'b00000000011101000000001110110011;
ROM[16920] <= 32'b00000000011100010010000000100011;
ROM[16921] <= 32'b00000000010000010000000100010011;
ROM[16922] <= 32'b11111111110000010000000100010011;
ROM[16923] <= 32'b00000000000000010010001110000011;
ROM[16924] <= 32'b00000000000000111000001100010011;
ROM[16925] <= 32'b00000000110100110000010000110011;
ROM[16926] <= 32'b00000000000001000010001110000011;
ROM[16927] <= 32'b00000000011100010010000000100011;
ROM[16928] <= 32'b00000000010000010000000100010011;
ROM[16929] <= 32'b00000100010001101010001110000011;
ROM[16930] <= 32'b00000000011100010010000000100011;
ROM[16931] <= 32'b00000000010000010000000100010011;
ROM[16932] <= 32'b00000100000000000000001110010011;
ROM[16933] <= 32'b00000000011100010010000000100011;
ROM[16934] <= 32'b00000000010000010000000100010011;
ROM[16935] <= 32'b11111111110000010000000100010011;
ROM[16936] <= 32'b00000000000000010010001110000011;
ROM[16937] <= 32'b11111111110000010000000100010011;
ROM[16938] <= 32'b00000000000000010010010000000011;
ROM[16939] <= 32'b00000000011101000000001110110011;
ROM[16940] <= 32'b00000000011100010010000000100011;
ROM[16941] <= 32'b00000000010000010000000100010011;
ROM[16942] <= 32'b11111111110000010000000100010011;
ROM[16943] <= 32'b00000000000000010010001110000011;
ROM[16944] <= 32'b00000000000000111000001100010011;
ROM[16945] <= 32'b00000000110100110000010000110011;
ROM[16946] <= 32'b00000000000001000010001110000011;
ROM[16947] <= 32'b00000000011100010010000000100011;
ROM[16948] <= 32'b00000000010000010000000100010011;
ROM[16949] <= 32'b11111111110000010000000100010011;
ROM[16950] <= 32'b00000000000000010010001110000011;
ROM[16951] <= 32'b11111111110000010000000100010011;
ROM[16952] <= 32'b00000000000000010010010000000011;
ROM[16953] <= 32'b00000000011101000000001110110011;
ROM[16954] <= 32'b00000000011100010010000000100011;
ROM[16955] <= 32'b00000000010000010000000100010011;
ROM[16956] <= 32'b00000100010001101010001110000011;
ROM[16957] <= 32'b00000000011100010010000000100011;
ROM[16958] <= 32'b00000000010000010000000100010011;
ROM[16959] <= 32'b00000100010000000000001110010011;
ROM[16960] <= 32'b00000000011100010010000000100011;
ROM[16961] <= 32'b00000000010000010000000100010011;
ROM[16962] <= 32'b11111111110000010000000100010011;
ROM[16963] <= 32'b00000000000000010010001110000011;
ROM[16964] <= 32'b11111111110000010000000100010011;
ROM[16965] <= 32'b00000000000000010010010000000011;
ROM[16966] <= 32'b00000000011101000000001110110011;
ROM[16967] <= 32'b00000000011100010010000000100011;
ROM[16968] <= 32'b00000000010000010000000100010011;
ROM[16969] <= 32'b11111111110000010000000100010011;
ROM[16970] <= 32'b00000000000000010010001110000011;
ROM[16971] <= 32'b00000000000000111000001100010011;
ROM[16972] <= 32'b11111111110000010000000100010011;
ROM[16973] <= 32'b00000000000000010010001110000011;
ROM[16974] <= 32'b00000000110100110000010000110011;
ROM[16975] <= 32'b00000000011101000010000000100011;
ROM[16976] <= 32'b00000100010001101010001110000011;
ROM[16977] <= 32'b00000000011100010010000000100011;
ROM[16978] <= 32'b00000000010000010000000100010011;
ROM[16979] <= 32'b00000100010000000000001110010011;
ROM[16980] <= 32'b00000000011100010010000000100011;
ROM[16981] <= 32'b00000000010000010000000100010011;
ROM[16982] <= 32'b11111111110000010000000100010011;
ROM[16983] <= 32'b00000000000000010010001110000011;
ROM[16984] <= 32'b11111111110000010000000100010011;
ROM[16985] <= 32'b00000000000000010010010000000011;
ROM[16986] <= 32'b00000000011101000000001110110011;
ROM[16987] <= 32'b00000000011100010010000000100011;
ROM[16988] <= 32'b00000000010000010000000100010011;
ROM[16989] <= 32'b11111111110000010000000100010011;
ROM[16990] <= 32'b00000000000000010010001110000011;
ROM[16991] <= 32'b00000000000000111000001100010011;
ROM[16992] <= 32'b00000000110100110000010000110011;
ROM[16993] <= 32'b00000000000001000010001110000011;
ROM[16994] <= 32'b00000000011100010010000000100011;
ROM[16995] <= 32'b00000000010000010000000100010011;
ROM[16996] <= 32'b00000100010001101010001110000011;
ROM[16997] <= 32'b00000000011100010010000000100011;
ROM[16998] <= 32'b00000000010000010000000100010011;
ROM[16999] <= 32'b00000100010000000000001110010011;
ROM[17000] <= 32'b00000000011100010010000000100011;
ROM[17001] <= 32'b00000000010000010000000100010011;
ROM[17002] <= 32'b11111111110000010000000100010011;
ROM[17003] <= 32'b00000000000000010010001110000011;
ROM[17004] <= 32'b11111111110000010000000100010011;
ROM[17005] <= 32'b00000000000000010010010000000011;
ROM[17006] <= 32'b00000000011101000000001110110011;
ROM[17007] <= 32'b00000000011100010010000000100011;
ROM[17008] <= 32'b00000000010000010000000100010011;
ROM[17009] <= 32'b11111111110000010000000100010011;
ROM[17010] <= 32'b00000000000000010010001110000011;
ROM[17011] <= 32'b00000000000000111000001100010011;
ROM[17012] <= 32'b00000000110100110000010000110011;
ROM[17013] <= 32'b00000000000001000010001110000011;
ROM[17014] <= 32'b00000000011100010010000000100011;
ROM[17015] <= 32'b00000000010000010000000100010011;
ROM[17016] <= 32'b11111111110000010000000100010011;
ROM[17017] <= 32'b00000000000000010010001110000011;
ROM[17018] <= 32'b11111111110000010000000100010011;
ROM[17019] <= 32'b00000000000000010010010000000011;
ROM[17020] <= 32'b00000000011101000000001110110011;
ROM[17021] <= 32'b00000000011100010010000000100011;
ROM[17022] <= 32'b00000000010000010000000100010011;
ROM[17023] <= 32'b00000100010001101010001110000011;
ROM[17024] <= 32'b00000000011100010010000000100011;
ROM[17025] <= 32'b00000000010000010000000100010011;
ROM[17026] <= 32'b00000100100000000000001110010011;
ROM[17027] <= 32'b00000000011100010010000000100011;
ROM[17028] <= 32'b00000000010000010000000100010011;
ROM[17029] <= 32'b11111111110000010000000100010011;
ROM[17030] <= 32'b00000000000000010010001110000011;
ROM[17031] <= 32'b11111111110000010000000100010011;
ROM[17032] <= 32'b00000000000000010010010000000011;
ROM[17033] <= 32'b00000000011101000000001110110011;
ROM[17034] <= 32'b00000000011100010010000000100011;
ROM[17035] <= 32'b00000000010000010000000100010011;
ROM[17036] <= 32'b11111111110000010000000100010011;
ROM[17037] <= 32'b00000000000000010010001110000011;
ROM[17038] <= 32'b00000000000000111000001100010011;
ROM[17039] <= 32'b11111111110000010000000100010011;
ROM[17040] <= 32'b00000000000000010010001110000011;
ROM[17041] <= 32'b00000000110100110000010000110011;
ROM[17042] <= 32'b00000000011101000010000000100011;
ROM[17043] <= 32'b00000100010001101010001110000011;
ROM[17044] <= 32'b00000000011100010010000000100011;
ROM[17045] <= 32'b00000000010000010000000100010011;
ROM[17046] <= 32'b00000100100000000000001110010011;
ROM[17047] <= 32'b00000000011100010010000000100011;
ROM[17048] <= 32'b00000000010000010000000100010011;
ROM[17049] <= 32'b11111111110000010000000100010011;
ROM[17050] <= 32'b00000000000000010010001110000011;
ROM[17051] <= 32'b11111111110000010000000100010011;
ROM[17052] <= 32'b00000000000000010010010000000011;
ROM[17053] <= 32'b00000000011101000000001110110011;
ROM[17054] <= 32'b00000000011100010010000000100011;
ROM[17055] <= 32'b00000000010000010000000100010011;
ROM[17056] <= 32'b11111111110000010000000100010011;
ROM[17057] <= 32'b00000000000000010010001110000011;
ROM[17058] <= 32'b00000000000000111000001100010011;
ROM[17059] <= 32'b00000000110100110000010000110011;
ROM[17060] <= 32'b00000000000001000010001110000011;
ROM[17061] <= 32'b00000000011100010010000000100011;
ROM[17062] <= 32'b00000000010000010000000100010011;
ROM[17063] <= 32'b00000100010001101010001110000011;
ROM[17064] <= 32'b00000000011100010010000000100011;
ROM[17065] <= 32'b00000000010000010000000100010011;
ROM[17066] <= 32'b00000100100000000000001110010011;
ROM[17067] <= 32'b00000000011100010010000000100011;
ROM[17068] <= 32'b00000000010000010000000100010011;
ROM[17069] <= 32'b11111111110000010000000100010011;
ROM[17070] <= 32'b00000000000000010010001110000011;
ROM[17071] <= 32'b11111111110000010000000100010011;
ROM[17072] <= 32'b00000000000000010010010000000011;
ROM[17073] <= 32'b00000000011101000000001110110011;
ROM[17074] <= 32'b00000000011100010010000000100011;
ROM[17075] <= 32'b00000000010000010000000100010011;
ROM[17076] <= 32'b11111111110000010000000100010011;
ROM[17077] <= 32'b00000000000000010010001110000011;
ROM[17078] <= 32'b00000000000000111000001100010011;
ROM[17079] <= 32'b00000000110100110000010000110011;
ROM[17080] <= 32'b00000000000001000010001110000011;
ROM[17081] <= 32'b00000000011100010010000000100011;
ROM[17082] <= 32'b00000000010000010000000100010011;
ROM[17083] <= 32'b11111111110000010000000100010011;
ROM[17084] <= 32'b00000000000000010010001110000011;
ROM[17085] <= 32'b11111111110000010000000100010011;
ROM[17086] <= 32'b00000000000000010010010000000011;
ROM[17087] <= 32'b00000000011101000000001110110011;
ROM[17088] <= 32'b00000000011100010010000000100011;
ROM[17089] <= 32'b00000000010000010000000100010011;
ROM[17090] <= 32'b00000100010001101010001110000011;
ROM[17091] <= 32'b00000000011100010010000000100011;
ROM[17092] <= 32'b00000000010000010000000100010011;
ROM[17093] <= 32'b00000100110000000000001110010011;
ROM[17094] <= 32'b00000000011100010010000000100011;
ROM[17095] <= 32'b00000000010000010000000100010011;
ROM[17096] <= 32'b11111111110000010000000100010011;
ROM[17097] <= 32'b00000000000000010010001110000011;
ROM[17098] <= 32'b11111111110000010000000100010011;
ROM[17099] <= 32'b00000000000000010010010000000011;
ROM[17100] <= 32'b00000000011101000000001110110011;
ROM[17101] <= 32'b00000000011100010010000000100011;
ROM[17102] <= 32'b00000000010000010000000100010011;
ROM[17103] <= 32'b11111111110000010000000100010011;
ROM[17104] <= 32'b00000000000000010010001110000011;
ROM[17105] <= 32'b00000000000000111000001100010011;
ROM[17106] <= 32'b11111111110000010000000100010011;
ROM[17107] <= 32'b00000000000000010010001110000011;
ROM[17108] <= 32'b00000000110100110000010000110011;
ROM[17109] <= 32'b00000000011101000010000000100011;
ROM[17110] <= 32'b00000100010001101010001110000011;
ROM[17111] <= 32'b00000000011100010010000000100011;
ROM[17112] <= 32'b00000000010000010000000100010011;
ROM[17113] <= 32'b00000100110000000000001110010011;
ROM[17114] <= 32'b00000000011100010010000000100011;
ROM[17115] <= 32'b00000000010000010000000100010011;
ROM[17116] <= 32'b11111111110000010000000100010011;
ROM[17117] <= 32'b00000000000000010010001110000011;
ROM[17118] <= 32'b11111111110000010000000100010011;
ROM[17119] <= 32'b00000000000000010010010000000011;
ROM[17120] <= 32'b00000000011101000000001110110011;
ROM[17121] <= 32'b00000000011100010010000000100011;
ROM[17122] <= 32'b00000000010000010000000100010011;
ROM[17123] <= 32'b11111111110000010000000100010011;
ROM[17124] <= 32'b00000000000000010010001110000011;
ROM[17125] <= 32'b00000000000000111000001100010011;
ROM[17126] <= 32'b00000000110100110000010000110011;
ROM[17127] <= 32'b00000000000001000010001110000011;
ROM[17128] <= 32'b00000000011100010010000000100011;
ROM[17129] <= 32'b00000000010000010000000100010011;
ROM[17130] <= 32'b00000100010001101010001110000011;
ROM[17131] <= 32'b00000000011100010010000000100011;
ROM[17132] <= 32'b00000000010000010000000100010011;
ROM[17133] <= 32'b00000100110000000000001110010011;
ROM[17134] <= 32'b00000000011100010010000000100011;
ROM[17135] <= 32'b00000000010000010000000100010011;
ROM[17136] <= 32'b11111111110000010000000100010011;
ROM[17137] <= 32'b00000000000000010010001110000011;
ROM[17138] <= 32'b11111111110000010000000100010011;
ROM[17139] <= 32'b00000000000000010010010000000011;
ROM[17140] <= 32'b00000000011101000000001110110011;
ROM[17141] <= 32'b00000000011100010010000000100011;
ROM[17142] <= 32'b00000000010000010000000100010011;
ROM[17143] <= 32'b11111111110000010000000100010011;
ROM[17144] <= 32'b00000000000000010010001110000011;
ROM[17145] <= 32'b00000000000000111000001100010011;
ROM[17146] <= 32'b00000000110100110000010000110011;
ROM[17147] <= 32'b00000000000001000010001110000011;
ROM[17148] <= 32'b00000000011100010010000000100011;
ROM[17149] <= 32'b00000000010000010000000100010011;
ROM[17150] <= 32'b11111111110000010000000100010011;
ROM[17151] <= 32'b00000000000000010010001110000011;
ROM[17152] <= 32'b11111111110000010000000100010011;
ROM[17153] <= 32'b00000000000000010010010000000011;
ROM[17154] <= 32'b00000000011101000000001110110011;
ROM[17155] <= 32'b00000000011100010010000000100011;
ROM[17156] <= 32'b00000000010000010000000100010011;
ROM[17157] <= 32'b00000100010001101010001110000011;
ROM[17158] <= 32'b00000000011100010010000000100011;
ROM[17159] <= 32'b00000000010000010000000100010011;
ROM[17160] <= 32'b00000101000000000000001110010011;
ROM[17161] <= 32'b00000000011100010010000000100011;
ROM[17162] <= 32'b00000000010000010000000100010011;
ROM[17163] <= 32'b11111111110000010000000100010011;
ROM[17164] <= 32'b00000000000000010010001110000011;
ROM[17165] <= 32'b11111111110000010000000100010011;
ROM[17166] <= 32'b00000000000000010010010000000011;
ROM[17167] <= 32'b00000000011101000000001110110011;
ROM[17168] <= 32'b00000000011100010010000000100011;
ROM[17169] <= 32'b00000000010000010000000100010011;
ROM[17170] <= 32'b11111111110000010000000100010011;
ROM[17171] <= 32'b00000000000000010010001110000011;
ROM[17172] <= 32'b00000000000000111000001100010011;
ROM[17173] <= 32'b11111111110000010000000100010011;
ROM[17174] <= 32'b00000000000000010010001110000011;
ROM[17175] <= 32'b00000000110100110000010000110011;
ROM[17176] <= 32'b00000000011101000010000000100011;
ROM[17177] <= 32'b00000100010001101010001110000011;
ROM[17178] <= 32'b00000000011100010010000000100011;
ROM[17179] <= 32'b00000000010000010000000100010011;
ROM[17180] <= 32'b00000101000000000000001110010011;
ROM[17181] <= 32'b00000000011100010010000000100011;
ROM[17182] <= 32'b00000000010000010000000100010011;
ROM[17183] <= 32'b11111111110000010000000100010011;
ROM[17184] <= 32'b00000000000000010010001110000011;
ROM[17185] <= 32'b11111111110000010000000100010011;
ROM[17186] <= 32'b00000000000000010010010000000011;
ROM[17187] <= 32'b00000000011101000000001110110011;
ROM[17188] <= 32'b00000000011100010010000000100011;
ROM[17189] <= 32'b00000000010000010000000100010011;
ROM[17190] <= 32'b11111111110000010000000100010011;
ROM[17191] <= 32'b00000000000000010010001110000011;
ROM[17192] <= 32'b00000000000000111000001100010011;
ROM[17193] <= 32'b00000000110100110000010000110011;
ROM[17194] <= 32'b00000000000001000010001110000011;
ROM[17195] <= 32'b00000000011100010010000000100011;
ROM[17196] <= 32'b00000000010000010000000100010011;
ROM[17197] <= 32'b00000100010001101010001110000011;
ROM[17198] <= 32'b00000000011100010010000000100011;
ROM[17199] <= 32'b00000000010000010000000100010011;
ROM[17200] <= 32'b00000101000000000000001110010011;
ROM[17201] <= 32'b00000000011100010010000000100011;
ROM[17202] <= 32'b00000000010000010000000100010011;
ROM[17203] <= 32'b11111111110000010000000100010011;
ROM[17204] <= 32'b00000000000000010010001110000011;
ROM[17205] <= 32'b11111111110000010000000100010011;
ROM[17206] <= 32'b00000000000000010010010000000011;
ROM[17207] <= 32'b00000000011101000000001110110011;
ROM[17208] <= 32'b00000000011100010010000000100011;
ROM[17209] <= 32'b00000000010000010000000100010011;
ROM[17210] <= 32'b11111111110000010000000100010011;
ROM[17211] <= 32'b00000000000000010010001110000011;
ROM[17212] <= 32'b00000000000000111000001100010011;
ROM[17213] <= 32'b00000000110100110000010000110011;
ROM[17214] <= 32'b00000000000001000010001110000011;
ROM[17215] <= 32'b00000000011100010010000000100011;
ROM[17216] <= 32'b00000000010000010000000100010011;
ROM[17217] <= 32'b11111111110000010000000100010011;
ROM[17218] <= 32'b00000000000000010010001110000011;
ROM[17219] <= 32'b11111111110000010000000100010011;
ROM[17220] <= 32'b00000000000000010010010000000011;
ROM[17221] <= 32'b00000000011101000000001110110011;
ROM[17222] <= 32'b00000000011100010010000000100011;
ROM[17223] <= 32'b00000000010000010000000100010011;
ROM[17224] <= 32'b00000100010001101010001110000011;
ROM[17225] <= 32'b00000000011100010010000000100011;
ROM[17226] <= 32'b00000000010000010000000100010011;
ROM[17227] <= 32'b00000101010000000000001110010011;
ROM[17228] <= 32'b00000000011100010010000000100011;
ROM[17229] <= 32'b00000000010000010000000100010011;
ROM[17230] <= 32'b11111111110000010000000100010011;
ROM[17231] <= 32'b00000000000000010010001110000011;
ROM[17232] <= 32'b11111111110000010000000100010011;
ROM[17233] <= 32'b00000000000000010010010000000011;
ROM[17234] <= 32'b00000000011101000000001110110011;
ROM[17235] <= 32'b00000000011100010010000000100011;
ROM[17236] <= 32'b00000000010000010000000100010011;
ROM[17237] <= 32'b11111111110000010000000100010011;
ROM[17238] <= 32'b00000000000000010010001110000011;
ROM[17239] <= 32'b00000000000000111000001100010011;
ROM[17240] <= 32'b11111111110000010000000100010011;
ROM[17241] <= 32'b00000000000000010010001110000011;
ROM[17242] <= 32'b00000000110100110000010000110011;
ROM[17243] <= 32'b00000000011101000010000000100011;
ROM[17244] <= 32'b00000100010001101010001110000011;
ROM[17245] <= 32'b00000000011100010010000000100011;
ROM[17246] <= 32'b00000000010000010000000100010011;
ROM[17247] <= 32'b00000101010000000000001110010011;
ROM[17248] <= 32'b00000000011100010010000000100011;
ROM[17249] <= 32'b00000000010000010000000100010011;
ROM[17250] <= 32'b11111111110000010000000100010011;
ROM[17251] <= 32'b00000000000000010010001110000011;
ROM[17252] <= 32'b11111111110000010000000100010011;
ROM[17253] <= 32'b00000000000000010010010000000011;
ROM[17254] <= 32'b00000000011101000000001110110011;
ROM[17255] <= 32'b00000000011100010010000000100011;
ROM[17256] <= 32'b00000000010000010000000100010011;
ROM[17257] <= 32'b11111111110000010000000100010011;
ROM[17258] <= 32'b00000000000000010010001110000011;
ROM[17259] <= 32'b00000000000000111000001100010011;
ROM[17260] <= 32'b00000000110100110000010000110011;
ROM[17261] <= 32'b00000000000001000010001110000011;
ROM[17262] <= 32'b00000000011100010010000000100011;
ROM[17263] <= 32'b00000000010000010000000100010011;
ROM[17264] <= 32'b00000100010001101010001110000011;
ROM[17265] <= 32'b00000000011100010010000000100011;
ROM[17266] <= 32'b00000000010000010000000100010011;
ROM[17267] <= 32'b00000101010000000000001110010011;
ROM[17268] <= 32'b00000000011100010010000000100011;
ROM[17269] <= 32'b00000000010000010000000100010011;
ROM[17270] <= 32'b11111111110000010000000100010011;
ROM[17271] <= 32'b00000000000000010010001110000011;
ROM[17272] <= 32'b11111111110000010000000100010011;
ROM[17273] <= 32'b00000000000000010010010000000011;
ROM[17274] <= 32'b00000000011101000000001110110011;
ROM[17275] <= 32'b00000000011100010010000000100011;
ROM[17276] <= 32'b00000000010000010000000100010011;
ROM[17277] <= 32'b11111111110000010000000100010011;
ROM[17278] <= 32'b00000000000000010010001110000011;
ROM[17279] <= 32'b00000000000000111000001100010011;
ROM[17280] <= 32'b00000000110100110000010000110011;
ROM[17281] <= 32'b00000000000001000010001110000011;
ROM[17282] <= 32'b00000000011100010010000000100011;
ROM[17283] <= 32'b00000000010000010000000100010011;
ROM[17284] <= 32'b11111111110000010000000100010011;
ROM[17285] <= 32'b00000000000000010010001110000011;
ROM[17286] <= 32'b11111111110000010000000100010011;
ROM[17287] <= 32'b00000000000000010010010000000011;
ROM[17288] <= 32'b00000000011101000000001110110011;
ROM[17289] <= 32'b00000000011100010010000000100011;
ROM[17290] <= 32'b00000000010000010000000100010011;
ROM[17291] <= 32'b00000100010001101010001110000011;
ROM[17292] <= 32'b00000000011100010010000000100011;
ROM[17293] <= 32'b00000000010000010000000100010011;
ROM[17294] <= 32'b00000101100000000000001110010011;
ROM[17295] <= 32'b00000000011100010010000000100011;
ROM[17296] <= 32'b00000000010000010000000100010011;
ROM[17297] <= 32'b11111111110000010000000100010011;
ROM[17298] <= 32'b00000000000000010010001110000011;
ROM[17299] <= 32'b11111111110000010000000100010011;
ROM[17300] <= 32'b00000000000000010010010000000011;
ROM[17301] <= 32'b00000000011101000000001110110011;
ROM[17302] <= 32'b00000000011100010010000000100011;
ROM[17303] <= 32'b00000000010000010000000100010011;
ROM[17304] <= 32'b11111111110000010000000100010011;
ROM[17305] <= 32'b00000000000000010010001110000011;
ROM[17306] <= 32'b00000000000000111000001100010011;
ROM[17307] <= 32'b11111111110000010000000100010011;
ROM[17308] <= 32'b00000000000000010010001110000011;
ROM[17309] <= 32'b00000000110100110000010000110011;
ROM[17310] <= 32'b00000000011101000010000000100011;
ROM[17311] <= 32'b00000100010001101010001110000011;
ROM[17312] <= 32'b00000000011100010010000000100011;
ROM[17313] <= 32'b00000000010000010000000100010011;
ROM[17314] <= 32'b00000101100000000000001110010011;
ROM[17315] <= 32'b00000000011100010010000000100011;
ROM[17316] <= 32'b00000000010000010000000100010011;
ROM[17317] <= 32'b11111111110000010000000100010011;
ROM[17318] <= 32'b00000000000000010010001110000011;
ROM[17319] <= 32'b11111111110000010000000100010011;
ROM[17320] <= 32'b00000000000000010010010000000011;
ROM[17321] <= 32'b00000000011101000000001110110011;
ROM[17322] <= 32'b00000000011100010010000000100011;
ROM[17323] <= 32'b00000000010000010000000100010011;
ROM[17324] <= 32'b11111111110000010000000100010011;
ROM[17325] <= 32'b00000000000000010010001110000011;
ROM[17326] <= 32'b00000000000000111000001100010011;
ROM[17327] <= 32'b00000000110100110000010000110011;
ROM[17328] <= 32'b00000000000001000010001110000011;
ROM[17329] <= 32'b00000000011100010010000000100011;
ROM[17330] <= 32'b00000000010000010000000100010011;
ROM[17331] <= 32'b00000100010001101010001110000011;
ROM[17332] <= 32'b00000000011100010010000000100011;
ROM[17333] <= 32'b00000000010000010000000100010011;
ROM[17334] <= 32'b00000101100000000000001110010011;
ROM[17335] <= 32'b00000000011100010010000000100011;
ROM[17336] <= 32'b00000000010000010000000100010011;
ROM[17337] <= 32'b11111111110000010000000100010011;
ROM[17338] <= 32'b00000000000000010010001110000011;
ROM[17339] <= 32'b11111111110000010000000100010011;
ROM[17340] <= 32'b00000000000000010010010000000011;
ROM[17341] <= 32'b00000000011101000000001110110011;
ROM[17342] <= 32'b00000000011100010010000000100011;
ROM[17343] <= 32'b00000000010000010000000100010011;
ROM[17344] <= 32'b11111111110000010000000100010011;
ROM[17345] <= 32'b00000000000000010010001110000011;
ROM[17346] <= 32'b00000000000000111000001100010011;
ROM[17347] <= 32'b00000000110100110000010000110011;
ROM[17348] <= 32'b00000000000001000010001110000011;
ROM[17349] <= 32'b00000000011100010010000000100011;
ROM[17350] <= 32'b00000000010000010000000100010011;
ROM[17351] <= 32'b11111111110000010000000100010011;
ROM[17352] <= 32'b00000000000000010010001110000011;
ROM[17353] <= 32'b11111111110000010000000100010011;
ROM[17354] <= 32'b00000000000000010010010000000011;
ROM[17355] <= 32'b00000000011101000000001110110011;
ROM[17356] <= 32'b00000000011100010010000000100011;
ROM[17357] <= 32'b00000000010000010000000100010011;
ROM[17358] <= 32'b00000100010001101010001110000011;
ROM[17359] <= 32'b00000000011100010010000000100011;
ROM[17360] <= 32'b00000000010000010000000100010011;
ROM[17361] <= 32'b00000101110000000000001110010011;
ROM[17362] <= 32'b00000000011100010010000000100011;
ROM[17363] <= 32'b00000000010000010000000100010011;
ROM[17364] <= 32'b11111111110000010000000100010011;
ROM[17365] <= 32'b00000000000000010010001110000011;
ROM[17366] <= 32'b11111111110000010000000100010011;
ROM[17367] <= 32'b00000000000000010010010000000011;
ROM[17368] <= 32'b00000000011101000000001110110011;
ROM[17369] <= 32'b00000000011100010010000000100011;
ROM[17370] <= 32'b00000000010000010000000100010011;
ROM[17371] <= 32'b11111111110000010000000100010011;
ROM[17372] <= 32'b00000000000000010010001110000011;
ROM[17373] <= 32'b00000000000000111000001100010011;
ROM[17374] <= 32'b11111111110000010000000100010011;
ROM[17375] <= 32'b00000000000000010010001110000011;
ROM[17376] <= 32'b00000000110100110000010000110011;
ROM[17377] <= 32'b00000000011101000010000000100011;
ROM[17378] <= 32'b00000100010001101010001110000011;
ROM[17379] <= 32'b00000000011100010010000000100011;
ROM[17380] <= 32'b00000000010000010000000100010011;
ROM[17381] <= 32'b00000101110000000000001110010011;
ROM[17382] <= 32'b00000000011100010010000000100011;
ROM[17383] <= 32'b00000000010000010000000100010011;
ROM[17384] <= 32'b11111111110000010000000100010011;
ROM[17385] <= 32'b00000000000000010010001110000011;
ROM[17386] <= 32'b11111111110000010000000100010011;
ROM[17387] <= 32'b00000000000000010010010000000011;
ROM[17388] <= 32'b00000000011101000000001110110011;
ROM[17389] <= 32'b00000000011100010010000000100011;
ROM[17390] <= 32'b00000000010000010000000100010011;
ROM[17391] <= 32'b11111111110000010000000100010011;
ROM[17392] <= 32'b00000000000000010010001110000011;
ROM[17393] <= 32'b00000000000000111000001100010011;
ROM[17394] <= 32'b00000000110100110000010000110011;
ROM[17395] <= 32'b00000000000001000010001110000011;
ROM[17396] <= 32'b00000000011100010010000000100011;
ROM[17397] <= 32'b00000000010000010000000100010011;
ROM[17398] <= 32'b00000100010001101010001110000011;
ROM[17399] <= 32'b00000000011100010010000000100011;
ROM[17400] <= 32'b00000000010000010000000100010011;
ROM[17401] <= 32'b00000101110000000000001110010011;
ROM[17402] <= 32'b00000000011100010010000000100011;
ROM[17403] <= 32'b00000000010000010000000100010011;
ROM[17404] <= 32'b11111111110000010000000100010011;
ROM[17405] <= 32'b00000000000000010010001110000011;
ROM[17406] <= 32'b11111111110000010000000100010011;
ROM[17407] <= 32'b00000000000000010010010000000011;
ROM[17408] <= 32'b00000000011101000000001110110011;
ROM[17409] <= 32'b00000000011100010010000000100011;
ROM[17410] <= 32'b00000000010000010000000100010011;
ROM[17411] <= 32'b11111111110000010000000100010011;
ROM[17412] <= 32'b00000000000000010010001110000011;
ROM[17413] <= 32'b00000000000000111000001100010011;
ROM[17414] <= 32'b00000000110100110000010000110011;
ROM[17415] <= 32'b00000000000001000010001110000011;
ROM[17416] <= 32'b00000000011100010010000000100011;
ROM[17417] <= 32'b00000000010000010000000100010011;
ROM[17418] <= 32'b11111111110000010000000100010011;
ROM[17419] <= 32'b00000000000000010010001110000011;
ROM[17420] <= 32'b11111111110000010000000100010011;
ROM[17421] <= 32'b00000000000000010010010000000011;
ROM[17422] <= 32'b00000000011101000000001110110011;
ROM[17423] <= 32'b00000000011100010010000000100011;
ROM[17424] <= 32'b00000000010000010000000100010011;
ROM[17425] <= 32'b00000100010001101010001110000011;
ROM[17426] <= 32'b00000000011100010010000000100011;
ROM[17427] <= 32'b00000000010000010000000100010011;
ROM[17428] <= 32'b00000110000000000000001110010011;
ROM[17429] <= 32'b00000000011100010010000000100011;
ROM[17430] <= 32'b00000000010000010000000100010011;
ROM[17431] <= 32'b11111111110000010000000100010011;
ROM[17432] <= 32'b00000000000000010010001110000011;
ROM[17433] <= 32'b11111111110000010000000100010011;
ROM[17434] <= 32'b00000000000000010010010000000011;
ROM[17435] <= 32'b00000000011101000000001110110011;
ROM[17436] <= 32'b00000000011100010010000000100011;
ROM[17437] <= 32'b00000000010000010000000100010011;
ROM[17438] <= 32'b11111111110000010000000100010011;
ROM[17439] <= 32'b00000000000000010010001110000011;
ROM[17440] <= 32'b00000000000000111000001100010011;
ROM[17441] <= 32'b11111111110000010000000100010011;
ROM[17442] <= 32'b00000000000000010010001110000011;
ROM[17443] <= 32'b00000000110100110000010000110011;
ROM[17444] <= 32'b00000000011101000010000000100011;
ROM[17445] <= 32'b00000100010001101010001110000011;
ROM[17446] <= 32'b00000000011100010010000000100011;
ROM[17447] <= 32'b00000000010000010000000100010011;
ROM[17448] <= 32'b00000110000000000000001110010011;
ROM[17449] <= 32'b00000000011100010010000000100011;
ROM[17450] <= 32'b00000000010000010000000100010011;
ROM[17451] <= 32'b11111111110000010000000100010011;
ROM[17452] <= 32'b00000000000000010010001110000011;
ROM[17453] <= 32'b11111111110000010000000100010011;
ROM[17454] <= 32'b00000000000000010010010000000011;
ROM[17455] <= 32'b00000000011101000000001110110011;
ROM[17456] <= 32'b00000000011100010010000000100011;
ROM[17457] <= 32'b00000000010000010000000100010011;
ROM[17458] <= 32'b11111111110000010000000100010011;
ROM[17459] <= 32'b00000000000000010010001110000011;
ROM[17460] <= 32'b00000000000000111000001100010011;
ROM[17461] <= 32'b00000000110100110000010000110011;
ROM[17462] <= 32'b00000000000001000010001110000011;
ROM[17463] <= 32'b00000000011100010010000000100011;
ROM[17464] <= 32'b00000000010000010000000100010011;
ROM[17465] <= 32'b00000100010001101010001110000011;
ROM[17466] <= 32'b00000000011100010010000000100011;
ROM[17467] <= 32'b00000000010000010000000100010011;
ROM[17468] <= 32'b00000110000000000000001110010011;
ROM[17469] <= 32'b00000000011100010010000000100011;
ROM[17470] <= 32'b00000000010000010000000100010011;
ROM[17471] <= 32'b11111111110000010000000100010011;
ROM[17472] <= 32'b00000000000000010010001110000011;
ROM[17473] <= 32'b11111111110000010000000100010011;
ROM[17474] <= 32'b00000000000000010010010000000011;
ROM[17475] <= 32'b00000000011101000000001110110011;
ROM[17476] <= 32'b00000000011100010010000000100011;
ROM[17477] <= 32'b00000000010000010000000100010011;
ROM[17478] <= 32'b11111111110000010000000100010011;
ROM[17479] <= 32'b00000000000000010010001110000011;
ROM[17480] <= 32'b00000000000000111000001100010011;
ROM[17481] <= 32'b00000000110100110000010000110011;
ROM[17482] <= 32'b00000000000001000010001110000011;
ROM[17483] <= 32'b00000000011100010010000000100011;
ROM[17484] <= 32'b00000000010000010000000100010011;
ROM[17485] <= 32'b11111111110000010000000100010011;
ROM[17486] <= 32'b00000000000000010010001110000011;
ROM[17487] <= 32'b11111111110000010000000100010011;
ROM[17488] <= 32'b00000000000000010010010000000011;
ROM[17489] <= 32'b00000000011101000000001110110011;
ROM[17490] <= 32'b00000000011100010010000000100011;
ROM[17491] <= 32'b00000000010000010000000100010011;
ROM[17492] <= 32'b00000100010001101010001110000011;
ROM[17493] <= 32'b00000000011100010010000000100011;
ROM[17494] <= 32'b00000000010000010000000100010011;
ROM[17495] <= 32'b00000110010000000000001110010011;
ROM[17496] <= 32'b00000000011100010010000000100011;
ROM[17497] <= 32'b00000000010000010000000100010011;
ROM[17498] <= 32'b11111111110000010000000100010011;
ROM[17499] <= 32'b00000000000000010010001110000011;
ROM[17500] <= 32'b11111111110000010000000100010011;
ROM[17501] <= 32'b00000000000000010010010000000011;
ROM[17502] <= 32'b00000000011101000000001110110011;
ROM[17503] <= 32'b00000000011100010010000000100011;
ROM[17504] <= 32'b00000000010000010000000100010011;
ROM[17505] <= 32'b11111111110000010000000100010011;
ROM[17506] <= 32'b00000000000000010010001110000011;
ROM[17507] <= 32'b00000000000000111000001100010011;
ROM[17508] <= 32'b11111111110000010000000100010011;
ROM[17509] <= 32'b00000000000000010010001110000011;
ROM[17510] <= 32'b00000000110100110000010000110011;
ROM[17511] <= 32'b00000000011101000010000000100011;
ROM[17512] <= 32'b00000100010001101010001110000011;
ROM[17513] <= 32'b00000000011100010010000000100011;
ROM[17514] <= 32'b00000000010000010000000100010011;
ROM[17515] <= 32'b00000110010000000000001110010011;
ROM[17516] <= 32'b00000000011100010010000000100011;
ROM[17517] <= 32'b00000000010000010000000100010011;
ROM[17518] <= 32'b11111111110000010000000100010011;
ROM[17519] <= 32'b00000000000000010010001110000011;
ROM[17520] <= 32'b11111111110000010000000100010011;
ROM[17521] <= 32'b00000000000000010010010000000011;
ROM[17522] <= 32'b00000000011101000000001110110011;
ROM[17523] <= 32'b00000000011100010010000000100011;
ROM[17524] <= 32'b00000000010000010000000100010011;
ROM[17525] <= 32'b11111111110000010000000100010011;
ROM[17526] <= 32'b00000000000000010010001110000011;
ROM[17527] <= 32'b00000000000000111000001100010011;
ROM[17528] <= 32'b00000000110100110000010000110011;
ROM[17529] <= 32'b00000000000001000010001110000011;
ROM[17530] <= 32'b00000000011100010010000000100011;
ROM[17531] <= 32'b00000000010000010000000100010011;
ROM[17532] <= 32'b00000100010001101010001110000011;
ROM[17533] <= 32'b00000000011100010010000000100011;
ROM[17534] <= 32'b00000000010000010000000100010011;
ROM[17535] <= 32'b00000110010000000000001110010011;
ROM[17536] <= 32'b00000000011100010010000000100011;
ROM[17537] <= 32'b00000000010000010000000100010011;
ROM[17538] <= 32'b11111111110000010000000100010011;
ROM[17539] <= 32'b00000000000000010010001110000011;
ROM[17540] <= 32'b11111111110000010000000100010011;
ROM[17541] <= 32'b00000000000000010010010000000011;
ROM[17542] <= 32'b00000000011101000000001110110011;
ROM[17543] <= 32'b00000000011100010010000000100011;
ROM[17544] <= 32'b00000000010000010000000100010011;
ROM[17545] <= 32'b11111111110000010000000100010011;
ROM[17546] <= 32'b00000000000000010010001110000011;
ROM[17547] <= 32'b00000000000000111000001100010011;
ROM[17548] <= 32'b00000000110100110000010000110011;
ROM[17549] <= 32'b00000000000001000010001110000011;
ROM[17550] <= 32'b00000000011100010010000000100011;
ROM[17551] <= 32'b00000000010000010000000100010011;
ROM[17552] <= 32'b11111111110000010000000100010011;
ROM[17553] <= 32'b00000000000000010010001110000011;
ROM[17554] <= 32'b11111111110000010000000100010011;
ROM[17555] <= 32'b00000000000000010010010000000011;
ROM[17556] <= 32'b00000000011101000000001110110011;
ROM[17557] <= 32'b00000000011100010010000000100011;
ROM[17558] <= 32'b00000000010000010000000100010011;
ROM[17559] <= 32'b00000100010001101010001110000011;
ROM[17560] <= 32'b00000000011100010010000000100011;
ROM[17561] <= 32'b00000000010000010000000100010011;
ROM[17562] <= 32'b00000110100000000000001110010011;
ROM[17563] <= 32'b00000000011100010010000000100011;
ROM[17564] <= 32'b00000000010000010000000100010011;
ROM[17565] <= 32'b11111111110000010000000100010011;
ROM[17566] <= 32'b00000000000000010010001110000011;
ROM[17567] <= 32'b11111111110000010000000100010011;
ROM[17568] <= 32'b00000000000000010010010000000011;
ROM[17569] <= 32'b00000000011101000000001110110011;
ROM[17570] <= 32'b00000000011100010010000000100011;
ROM[17571] <= 32'b00000000010000010000000100010011;
ROM[17572] <= 32'b11111111110000010000000100010011;
ROM[17573] <= 32'b00000000000000010010001110000011;
ROM[17574] <= 32'b00000000000000111000001100010011;
ROM[17575] <= 32'b11111111110000010000000100010011;
ROM[17576] <= 32'b00000000000000010010001110000011;
ROM[17577] <= 32'b00000000110100110000010000110011;
ROM[17578] <= 32'b00000000011101000010000000100011;
ROM[17579] <= 32'b00000100010001101010001110000011;
ROM[17580] <= 32'b00000000011100010010000000100011;
ROM[17581] <= 32'b00000000010000010000000100010011;
ROM[17582] <= 32'b00000110100000000000001110010011;
ROM[17583] <= 32'b00000000011100010010000000100011;
ROM[17584] <= 32'b00000000010000010000000100010011;
ROM[17585] <= 32'b11111111110000010000000100010011;
ROM[17586] <= 32'b00000000000000010010001110000011;
ROM[17587] <= 32'b11111111110000010000000100010011;
ROM[17588] <= 32'b00000000000000010010010000000011;
ROM[17589] <= 32'b00000000011101000000001110110011;
ROM[17590] <= 32'b00000000011100010010000000100011;
ROM[17591] <= 32'b00000000010000010000000100010011;
ROM[17592] <= 32'b11111111110000010000000100010011;
ROM[17593] <= 32'b00000000000000010010001110000011;
ROM[17594] <= 32'b00000000000000111000001100010011;
ROM[17595] <= 32'b00000000110100110000010000110011;
ROM[17596] <= 32'b00000000000001000010001110000011;
ROM[17597] <= 32'b00000000011100010010000000100011;
ROM[17598] <= 32'b00000000010000010000000100010011;
ROM[17599] <= 32'b00000100010001101010001110000011;
ROM[17600] <= 32'b00000000011100010010000000100011;
ROM[17601] <= 32'b00000000010000010000000100010011;
ROM[17602] <= 32'b00000110100000000000001110010011;
ROM[17603] <= 32'b00000000011100010010000000100011;
ROM[17604] <= 32'b00000000010000010000000100010011;
ROM[17605] <= 32'b11111111110000010000000100010011;
ROM[17606] <= 32'b00000000000000010010001110000011;
ROM[17607] <= 32'b11111111110000010000000100010011;
ROM[17608] <= 32'b00000000000000010010010000000011;
ROM[17609] <= 32'b00000000011101000000001110110011;
ROM[17610] <= 32'b00000000011100010010000000100011;
ROM[17611] <= 32'b00000000010000010000000100010011;
ROM[17612] <= 32'b11111111110000010000000100010011;
ROM[17613] <= 32'b00000000000000010010001110000011;
ROM[17614] <= 32'b00000000000000111000001100010011;
ROM[17615] <= 32'b00000000110100110000010000110011;
ROM[17616] <= 32'b00000000000001000010001110000011;
ROM[17617] <= 32'b00000000011100010010000000100011;
ROM[17618] <= 32'b00000000010000010000000100010011;
ROM[17619] <= 32'b11111111110000010000000100010011;
ROM[17620] <= 32'b00000000000000010010001110000011;
ROM[17621] <= 32'b11111111110000010000000100010011;
ROM[17622] <= 32'b00000000000000010010010000000011;
ROM[17623] <= 32'b00000000011101000000001110110011;
ROM[17624] <= 32'b00000000011100010010000000100011;
ROM[17625] <= 32'b00000000010000010000000100010011;
ROM[17626] <= 32'b00000100010001101010001110000011;
ROM[17627] <= 32'b00000000011100010010000000100011;
ROM[17628] <= 32'b00000000010000010000000100010011;
ROM[17629] <= 32'b00000110110000000000001110010011;
ROM[17630] <= 32'b00000000011100010010000000100011;
ROM[17631] <= 32'b00000000010000010000000100010011;
ROM[17632] <= 32'b11111111110000010000000100010011;
ROM[17633] <= 32'b00000000000000010010001110000011;
ROM[17634] <= 32'b11111111110000010000000100010011;
ROM[17635] <= 32'b00000000000000010010010000000011;
ROM[17636] <= 32'b00000000011101000000001110110011;
ROM[17637] <= 32'b00000000011100010010000000100011;
ROM[17638] <= 32'b00000000010000010000000100010011;
ROM[17639] <= 32'b11111111110000010000000100010011;
ROM[17640] <= 32'b00000000000000010010001110000011;
ROM[17641] <= 32'b00000000000000111000001100010011;
ROM[17642] <= 32'b11111111110000010000000100010011;
ROM[17643] <= 32'b00000000000000010010001110000011;
ROM[17644] <= 32'b00000000110100110000010000110011;
ROM[17645] <= 32'b00000000011101000010000000100011;
ROM[17646] <= 32'b00000100010001101010001110000011;
ROM[17647] <= 32'b00000000011100010010000000100011;
ROM[17648] <= 32'b00000000010000010000000100010011;
ROM[17649] <= 32'b00000110110000000000001110010011;
ROM[17650] <= 32'b00000000011100010010000000100011;
ROM[17651] <= 32'b00000000010000010000000100010011;
ROM[17652] <= 32'b11111111110000010000000100010011;
ROM[17653] <= 32'b00000000000000010010001110000011;
ROM[17654] <= 32'b11111111110000010000000100010011;
ROM[17655] <= 32'b00000000000000010010010000000011;
ROM[17656] <= 32'b00000000011101000000001110110011;
ROM[17657] <= 32'b00000000011100010010000000100011;
ROM[17658] <= 32'b00000000010000010000000100010011;
ROM[17659] <= 32'b11111111110000010000000100010011;
ROM[17660] <= 32'b00000000000000010010001110000011;
ROM[17661] <= 32'b00000000000000111000001100010011;
ROM[17662] <= 32'b00000000110100110000010000110011;
ROM[17663] <= 32'b00000000000001000010001110000011;
ROM[17664] <= 32'b00000000011100010010000000100011;
ROM[17665] <= 32'b00000000010000010000000100010011;
ROM[17666] <= 32'b00000100010001101010001110000011;
ROM[17667] <= 32'b00000000011100010010000000100011;
ROM[17668] <= 32'b00000000010000010000000100010011;
ROM[17669] <= 32'b00000110110000000000001110010011;
ROM[17670] <= 32'b00000000011100010010000000100011;
ROM[17671] <= 32'b00000000010000010000000100010011;
ROM[17672] <= 32'b11111111110000010000000100010011;
ROM[17673] <= 32'b00000000000000010010001110000011;
ROM[17674] <= 32'b11111111110000010000000100010011;
ROM[17675] <= 32'b00000000000000010010010000000011;
ROM[17676] <= 32'b00000000011101000000001110110011;
ROM[17677] <= 32'b00000000011100010010000000100011;
ROM[17678] <= 32'b00000000010000010000000100010011;
ROM[17679] <= 32'b11111111110000010000000100010011;
ROM[17680] <= 32'b00000000000000010010001110000011;
ROM[17681] <= 32'b00000000000000111000001100010011;
ROM[17682] <= 32'b00000000110100110000010000110011;
ROM[17683] <= 32'b00000000000001000010001110000011;
ROM[17684] <= 32'b00000000011100010010000000100011;
ROM[17685] <= 32'b00000000010000010000000100010011;
ROM[17686] <= 32'b11111111110000010000000100010011;
ROM[17687] <= 32'b00000000000000010010001110000011;
ROM[17688] <= 32'b11111111110000010000000100010011;
ROM[17689] <= 32'b00000000000000010010010000000011;
ROM[17690] <= 32'b00000000011101000000001110110011;
ROM[17691] <= 32'b00000000011100010010000000100011;
ROM[17692] <= 32'b00000000010000010000000100010011;
ROM[17693] <= 32'b00000100010001101010001110000011;
ROM[17694] <= 32'b00000000011100010010000000100011;
ROM[17695] <= 32'b00000000010000010000000100010011;
ROM[17696] <= 32'b00000111000000000000001110010011;
ROM[17697] <= 32'b00000000011100010010000000100011;
ROM[17698] <= 32'b00000000010000010000000100010011;
ROM[17699] <= 32'b11111111110000010000000100010011;
ROM[17700] <= 32'b00000000000000010010001110000011;
ROM[17701] <= 32'b11111111110000010000000100010011;
ROM[17702] <= 32'b00000000000000010010010000000011;
ROM[17703] <= 32'b00000000011101000000001110110011;
ROM[17704] <= 32'b00000000011100010010000000100011;
ROM[17705] <= 32'b00000000010000010000000100010011;
ROM[17706] <= 32'b11111111110000010000000100010011;
ROM[17707] <= 32'b00000000000000010010001110000011;
ROM[17708] <= 32'b00000000000000111000001100010011;
ROM[17709] <= 32'b11111111110000010000000100010011;
ROM[17710] <= 32'b00000000000000010010001110000011;
ROM[17711] <= 32'b00000000110100110000010000110011;
ROM[17712] <= 32'b00000000011101000010000000100011;
ROM[17713] <= 32'b00000100010001101010001110000011;
ROM[17714] <= 32'b00000000011100010010000000100011;
ROM[17715] <= 32'b00000000010000010000000100010011;
ROM[17716] <= 32'b00000111000000000000001110010011;
ROM[17717] <= 32'b00000000011100010010000000100011;
ROM[17718] <= 32'b00000000010000010000000100010011;
ROM[17719] <= 32'b11111111110000010000000100010011;
ROM[17720] <= 32'b00000000000000010010001110000011;
ROM[17721] <= 32'b11111111110000010000000100010011;
ROM[17722] <= 32'b00000000000000010010010000000011;
ROM[17723] <= 32'b00000000011101000000001110110011;
ROM[17724] <= 32'b00000000011100010010000000100011;
ROM[17725] <= 32'b00000000010000010000000100010011;
ROM[17726] <= 32'b11111111110000010000000100010011;
ROM[17727] <= 32'b00000000000000010010001110000011;
ROM[17728] <= 32'b00000000000000111000001100010011;
ROM[17729] <= 32'b00000000110100110000010000110011;
ROM[17730] <= 32'b00000000000001000010001110000011;
ROM[17731] <= 32'b00000000011100010010000000100011;
ROM[17732] <= 32'b00000000010000010000000100010011;
ROM[17733] <= 32'b00000100010001101010001110000011;
ROM[17734] <= 32'b00000000011100010010000000100011;
ROM[17735] <= 32'b00000000010000010000000100010011;
ROM[17736] <= 32'b00000111000000000000001110010011;
ROM[17737] <= 32'b00000000011100010010000000100011;
ROM[17738] <= 32'b00000000010000010000000100010011;
ROM[17739] <= 32'b11111111110000010000000100010011;
ROM[17740] <= 32'b00000000000000010010001110000011;
ROM[17741] <= 32'b11111111110000010000000100010011;
ROM[17742] <= 32'b00000000000000010010010000000011;
ROM[17743] <= 32'b00000000011101000000001110110011;
ROM[17744] <= 32'b00000000011100010010000000100011;
ROM[17745] <= 32'b00000000010000010000000100010011;
ROM[17746] <= 32'b11111111110000010000000100010011;
ROM[17747] <= 32'b00000000000000010010001110000011;
ROM[17748] <= 32'b00000000000000111000001100010011;
ROM[17749] <= 32'b00000000110100110000010000110011;
ROM[17750] <= 32'b00000000000001000010001110000011;
ROM[17751] <= 32'b00000000011100010010000000100011;
ROM[17752] <= 32'b00000000010000010000000100010011;
ROM[17753] <= 32'b11111111110000010000000100010011;
ROM[17754] <= 32'b00000000000000010010001110000011;
ROM[17755] <= 32'b11111111110000010000000100010011;
ROM[17756] <= 32'b00000000000000010010010000000011;
ROM[17757] <= 32'b00000000011101000000001110110011;
ROM[17758] <= 32'b00000000011100010010000000100011;
ROM[17759] <= 32'b00000000010000010000000100010011;
ROM[17760] <= 32'b00000100010001101010001110000011;
ROM[17761] <= 32'b00000000011100010010000000100011;
ROM[17762] <= 32'b00000000010000010000000100010011;
ROM[17763] <= 32'b00000111010000000000001110010011;
ROM[17764] <= 32'b00000000011100010010000000100011;
ROM[17765] <= 32'b00000000010000010000000100010011;
ROM[17766] <= 32'b11111111110000010000000100010011;
ROM[17767] <= 32'b00000000000000010010001110000011;
ROM[17768] <= 32'b11111111110000010000000100010011;
ROM[17769] <= 32'b00000000000000010010010000000011;
ROM[17770] <= 32'b00000000011101000000001110110011;
ROM[17771] <= 32'b00000000011100010010000000100011;
ROM[17772] <= 32'b00000000010000010000000100010011;
ROM[17773] <= 32'b11111111110000010000000100010011;
ROM[17774] <= 32'b00000000000000010010001110000011;
ROM[17775] <= 32'b00000000000000111000001100010011;
ROM[17776] <= 32'b11111111110000010000000100010011;
ROM[17777] <= 32'b00000000000000010010001110000011;
ROM[17778] <= 32'b00000000110100110000010000110011;
ROM[17779] <= 32'b00000000011101000010000000100011;
ROM[17780] <= 32'b00000100010001101010001110000011;
ROM[17781] <= 32'b00000000011100010010000000100011;
ROM[17782] <= 32'b00000000010000010000000100010011;
ROM[17783] <= 32'b00000111010000000000001110010011;
ROM[17784] <= 32'b00000000011100010010000000100011;
ROM[17785] <= 32'b00000000010000010000000100010011;
ROM[17786] <= 32'b11111111110000010000000100010011;
ROM[17787] <= 32'b00000000000000010010001110000011;
ROM[17788] <= 32'b11111111110000010000000100010011;
ROM[17789] <= 32'b00000000000000010010010000000011;
ROM[17790] <= 32'b00000000011101000000001110110011;
ROM[17791] <= 32'b00000000011100010010000000100011;
ROM[17792] <= 32'b00000000010000010000000100010011;
ROM[17793] <= 32'b11111111110000010000000100010011;
ROM[17794] <= 32'b00000000000000010010001110000011;
ROM[17795] <= 32'b00000000000000111000001100010011;
ROM[17796] <= 32'b00000000110100110000010000110011;
ROM[17797] <= 32'b00000000000001000010001110000011;
ROM[17798] <= 32'b00000000011100010010000000100011;
ROM[17799] <= 32'b00000000010000010000000100010011;
ROM[17800] <= 32'b00000100010001101010001110000011;
ROM[17801] <= 32'b00000000011100010010000000100011;
ROM[17802] <= 32'b00000000010000010000000100010011;
ROM[17803] <= 32'b00000111010000000000001110010011;
ROM[17804] <= 32'b00000000011100010010000000100011;
ROM[17805] <= 32'b00000000010000010000000100010011;
ROM[17806] <= 32'b11111111110000010000000100010011;
ROM[17807] <= 32'b00000000000000010010001110000011;
ROM[17808] <= 32'b11111111110000010000000100010011;
ROM[17809] <= 32'b00000000000000010010010000000011;
ROM[17810] <= 32'b00000000011101000000001110110011;
ROM[17811] <= 32'b00000000011100010010000000100011;
ROM[17812] <= 32'b00000000010000010000000100010011;
ROM[17813] <= 32'b11111111110000010000000100010011;
ROM[17814] <= 32'b00000000000000010010001110000011;
ROM[17815] <= 32'b00000000000000111000001100010011;
ROM[17816] <= 32'b00000000110100110000010000110011;
ROM[17817] <= 32'b00000000000001000010001110000011;
ROM[17818] <= 32'b00000000011100010010000000100011;
ROM[17819] <= 32'b00000000010000010000000100010011;
ROM[17820] <= 32'b11111111110000010000000100010011;
ROM[17821] <= 32'b00000000000000010010001110000011;
ROM[17822] <= 32'b11111111110000010000000100010011;
ROM[17823] <= 32'b00000000000000010010010000000011;
ROM[17824] <= 32'b00000000011101000000001110110011;
ROM[17825] <= 32'b00000000011100010010000000100011;
ROM[17826] <= 32'b00000000010000010000000100010011;
ROM[17827] <= 32'b00000100010001101010001110000011;
ROM[17828] <= 32'b00000000011100010010000000100011;
ROM[17829] <= 32'b00000000010000010000000100010011;
ROM[17830] <= 32'b00000111100000000000001110010011;
ROM[17831] <= 32'b00000000011100010010000000100011;
ROM[17832] <= 32'b00000000010000010000000100010011;
ROM[17833] <= 32'b11111111110000010000000100010011;
ROM[17834] <= 32'b00000000000000010010001110000011;
ROM[17835] <= 32'b11111111110000010000000100010011;
ROM[17836] <= 32'b00000000000000010010010000000011;
ROM[17837] <= 32'b00000000011101000000001110110011;
ROM[17838] <= 32'b00000000011100010010000000100011;
ROM[17839] <= 32'b00000000010000010000000100010011;
ROM[17840] <= 32'b11111111110000010000000100010011;
ROM[17841] <= 32'b00000000000000010010001110000011;
ROM[17842] <= 32'b00000000000000111000001100010011;
ROM[17843] <= 32'b11111111110000010000000100010011;
ROM[17844] <= 32'b00000000000000010010001110000011;
ROM[17845] <= 32'b00000000110100110000010000110011;
ROM[17846] <= 32'b00000000011101000010000000100011;
ROM[17847] <= 32'b00000100010001101010001110000011;
ROM[17848] <= 32'b00000000011100010010000000100011;
ROM[17849] <= 32'b00000000010000010000000100010011;
ROM[17850] <= 32'b00000111100000000000001110010011;
ROM[17851] <= 32'b00000000011100010010000000100011;
ROM[17852] <= 32'b00000000010000010000000100010011;
ROM[17853] <= 32'b11111111110000010000000100010011;
ROM[17854] <= 32'b00000000000000010010001110000011;
ROM[17855] <= 32'b11111111110000010000000100010011;
ROM[17856] <= 32'b00000000000000010010010000000011;
ROM[17857] <= 32'b00000000011101000000001110110011;
ROM[17858] <= 32'b00000000011100010010000000100011;
ROM[17859] <= 32'b00000000010000010000000100010011;
ROM[17860] <= 32'b11111111110000010000000100010011;
ROM[17861] <= 32'b00000000000000010010001110000011;
ROM[17862] <= 32'b00000000000000111000001100010011;
ROM[17863] <= 32'b00000000110100110000010000110011;
ROM[17864] <= 32'b00000000000001000010001110000011;
ROM[17865] <= 32'b00000000011100010010000000100011;
ROM[17866] <= 32'b00000000010000010000000100010011;
ROM[17867] <= 32'b00000100010001101010001110000011;
ROM[17868] <= 32'b00000000011100010010000000100011;
ROM[17869] <= 32'b00000000010000010000000100010011;
ROM[17870] <= 32'b00000111100000000000001110010011;
ROM[17871] <= 32'b00000000011100010010000000100011;
ROM[17872] <= 32'b00000000010000010000000100010011;
ROM[17873] <= 32'b11111111110000010000000100010011;
ROM[17874] <= 32'b00000000000000010010001110000011;
ROM[17875] <= 32'b11111111110000010000000100010011;
ROM[17876] <= 32'b00000000000000010010010000000011;
ROM[17877] <= 32'b00000000011101000000001110110011;
ROM[17878] <= 32'b00000000011100010010000000100011;
ROM[17879] <= 32'b00000000010000010000000100010011;
ROM[17880] <= 32'b11111111110000010000000100010011;
ROM[17881] <= 32'b00000000000000010010001110000011;
ROM[17882] <= 32'b00000000000000111000001100010011;
ROM[17883] <= 32'b00000000110100110000010000110011;
ROM[17884] <= 32'b00000000000001000010001110000011;
ROM[17885] <= 32'b00000000011100010010000000100011;
ROM[17886] <= 32'b00000000010000010000000100010011;
ROM[17887] <= 32'b11111111110000010000000100010011;
ROM[17888] <= 32'b00000000000000010010001110000011;
ROM[17889] <= 32'b11111111110000010000000100010011;
ROM[17890] <= 32'b00000000000000010010010000000011;
ROM[17891] <= 32'b00000000011101000000001110110011;
ROM[17892] <= 32'b00000000011100010010000000100011;
ROM[17893] <= 32'b00000000010000010000000100010011;
ROM[17894] <= 32'b00000100010001101010001110000011;
ROM[17895] <= 32'b00000000011100010010000000100011;
ROM[17896] <= 32'b00000000010000010000000100010011;
ROM[17897] <= 32'b00000111110000000000001110010011;
ROM[17898] <= 32'b00000000011100010010000000100011;
ROM[17899] <= 32'b00000000010000010000000100010011;
ROM[17900] <= 32'b11111111110000010000000100010011;
ROM[17901] <= 32'b00000000000000010010001110000011;
ROM[17902] <= 32'b11111111110000010000000100010011;
ROM[17903] <= 32'b00000000000000010010010000000011;
ROM[17904] <= 32'b00000000011101000000001110110011;
ROM[17905] <= 32'b00000000011100010010000000100011;
ROM[17906] <= 32'b00000000010000010000000100010011;
ROM[17907] <= 32'b11111111110000010000000100010011;
ROM[17908] <= 32'b00000000000000010010001110000011;
ROM[17909] <= 32'b00000000000000111000001100010011;
ROM[17910] <= 32'b11111111110000010000000100010011;
ROM[17911] <= 32'b00000000000000010010001110000011;
ROM[17912] <= 32'b00000000110100110000010000110011;
ROM[17913] <= 32'b00000000011101000010000000100011;
ROM[17914] <= 32'b00000000000000000000001110010011;
ROM[17915] <= 32'b00000000011100010010000000100011;
ROM[17916] <= 32'b00000000010000010000000100010011;
ROM[17917] <= 32'b00000001010000000000001110010011;
ROM[17918] <= 32'b01000000011100011000001110110011;
ROM[17919] <= 32'b00000000000000111010000010000011;
ROM[17920] <= 32'b11111111110000010000000100010011;
ROM[17921] <= 32'b00000000000000010010001110000011;
ROM[17922] <= 32'b00000000011100100010000000100011;
ROM[17923] <= 32'b00000000010000100000000100010011;
ROM[17924] <= 32'b00000001010000000000001110010011;
ROM[17925] <= 32'b01000000011100011000001110110011;
ROM[17926] <= 32'b00000000010000111010000110000011;
ROM[17927] <= 32'b00000000100000111010001000000011;
ROM[17928] <= 32'b00000000110000111010001010000011;
ROM[17929] <= 32'b00000001000000111010001100000011;
ROM[17930] <= 32'b00000000000000001000000011100111;
ROM[17931] <= 32'b00000000000000010010000000100011;
ROM[17932] <= 32'b00000000010000010000000100010011;
ROM[17933] <= 32'b00000000000000010010000000100011;
ROM[17934] <= 32'b00000000010000010000000100010011;
ROM[17935] <= 32'b00000000000000010010000000100011;
ROM[17936] <= 32'b00000000010000010000000100010011;
ROM[17937] <= 32'b00000000000000000000001110010011;
ROM[17938] <= 32'b00000000011100010010000000100011;
ROM[17939] <= 32'b00000000010000010000000100010011;
ROM[17940] <= 32'b11111111110000010000000100010011;
ROM[17941] <= 32'b00000000000000010010001110000011;
ROM[17942] <= 32'b00000000011100011010000000100011;
ROM[17943] <= 32'b00000000000000100010001110000011;
ROM[17944] <= 32'b00000000011100010010000000100011;
ROM[17945] <= 32'b00000000010000010000000100010011;
ROM[17946] <= 32'b11111111110000010000000100010011;
ROM[17947] <= 32'b00000000000000010010001110000011;
ROM[17948] <= 32'b00000000011100011010001000100011;
ROM[17949] <= 32'b00000000000000000000001110010011;
ROM[17950] <= 32'b00000000011100010010000000100011;
ROM[17951] <= 32'b00000000010000010000000100010011;
ROM[17952] <= 32'b11111111110000010000000100010011;
ROM[17953] <= 32'b00000000000000010010001110000011;
ROM[17954] <= 32'b00000000011100011010010000100011;
ROM[17955] <= 32'b00000000100000011010001110000011;
ROM[17956] <= 32'b00000000011100010010000000100011;
ROM[17957] <= 32'b00000000010000010000000100010011;
ROM[17958] <= 32'b00001000000000000000001110010011;
ROM[17959] <= 32'b00000000011100010010000000100011;
ROM[17960] <= 32'b00000000010000010000000100010011;
ROM[17961] <= 32'b11111111110000010000000100010011;
ROM[17962] <= 32'b00000000000000010010001110000011;
ROM[17963] <= 32'b11111111110000010000000100010011;
ROM[17964] <= 32'b00000000000000010010010000000011;
ROM[17965] <= 32'b00000000011101000010001110110011;
ROM[17966] <= 32'b00000000011100010010000000100011;
ROM[17967] <= 32'b00000000010000010000000100010011;
ROM[17968] <= 32'b11111111110000010000000100010011;
ROM[17969] <= 32'b00000000000000010010001110000011;
ROM[17970] <= 32'b01000000011100000000001110110011;
ROM[17971] <= 32'b00000000000100111000001110010011;
ROM[17972] <= 32'b00000000011100010010000000100011;
ROM[17973] <= 32'b00000000010000010000000100010011;
ROM[17974] <= 32'b11111111110000010000000100010011;
ROM[17975] <= 32'b00000000000000010010001110000011;
ROM[17976] <= 32'b00000000000000111000101001100011;
ROM[17977] <= 32'b00000000000000010010001110110111;
ROM[17978] <= 32'b10101010000000111000001110010011;
ROM[17979] <= 32'b00000000111000111000001110110011;
ROM[17980] <= 32'b00000000000000111000000011100111;
ROM[17981] <= 32'b00000000010000100010001110000011;
ROM[17982] <= 32'b00000000011100010010000000100011;
ROM[17983] <= 32'b00000000010000010000000100010011;
ROM[17984] <= 32'b00000100010001101010001110000011;
ROM[17985] <= 32'b00000000011100010010000000100011;
ROM[17986] <= 32'b00000000010000010000000100010011;
ROM[17987] <= 32'b00000000100000011010001110000011;
ROM[17988] <= 32'b00000000011100010010000000100011;
ROM[17989] <= 32'b00000000010000010000000100010011;
ROM[17990] <= 32'b11111111110000010000000100010011;
ROM[17991] <= 32'b00000000000000010010001110000011;
ROM[17992] <= 32'b11111111110000010000000100010011;
ROM[17993] <= 32'b00000000000000010010010000000011;
ROM[17994] <= 32'b00000000011101000000001110110011;
ROM[17995] <= 32'b00000000011100010010000000100011;
ROM[17996] <= 32'b00000000010000010000000100010011;
ROM[17997] <= 32'b11111111110000010000000100010011;
ROM[17998] <= 32'b00000000000000010010001110000011;
ROM[17999] <= 32'b00000000000000111000001100010011;
ROM[18000] <= 32'b00000000110100110000010000110011;
ROM[18001] <= 32'b00000000000001000010001110000011;
ROM[18002] <= 32'b00000000011100010010000000100011;
ROM[18003] <= 32'b00000000010000010000000100010011;
ROM[18004] <= 32'b11111111110000010000000100010011;
ROM[18005] <= 32'b00000000000000010010001110000011;
ROM[18006] <= 32'b11111111110000010000000100010011;
ROM[18007] <= 32'b00000000000000010010010000000011;
ROM[18008] <= 32'b00000000011101000111001110110011;
ROM[18009] <= 32'b00000000011100010010000000100011;
ROM[18010] <= 32'b00000000010000010000000100010011;
ROM[18011] <= 32'b00000000000000000000001110010011;
ROM[18012] <= 32'b00000000011100010010000000100011;
ROM[18013] <= 32'b00000000010000010000000100010011;
ROM[18014] <= 32'b11111111110000010000000100010011;
ROM[18015] <= 32'b00000000000000010010001110000011;
ROM[18016] <= 32'b11111111110000010000000100010011;
ROM[18017] <= 32'b00000000000000010010010000000011;
ROM[18018] <= 32'b00000000011101000010010010110011;
ROM[18019] <= 32'b00000000100000111010010100110011;
ROM[18020] <= 32'b00000000101001001000001110110011;
ROM[18021] <= 32'b00000000000100111000001110010011;
ROM[18022] <= 32'b00000000000100111111001110010011;
ROM[18023] <= 32'b00000000011100010010000000100011;
ROM[18024] <= 32'b00000000010000010000000100010011;
ROM[18025] <= 32'b11111111110000010000000100010011;
ROM[18026] <= 32'b00000000000000010010001110000011;
ROM[18027] <= 32'b01000000011100000000001110110011;
ROM[18028] <= 32'b00000000000100111000001110010011;
ROM[18029] <= 32'b00000000011100010010000000100011;
ROM[18030] <= 32'b00000000010000010000000100010011;
ROM[18031] <= 32'b11111111110000010000000100010011;
ROM[18032] <= 32'b00000000000000010010001110000011;
ROM[18033] <= 32'b00000000000000111000101001100011;
ROM[18034] <= 32'b00000000000000010010001110110111;
ROM[18035] <= 32'b10011101110000111000001110010011;
ROM[18036] <= 32'b00000000111000111000001110110011;
ROM[18037] <= 32'b00000000000000111000000011100111;
ROM[18038] <= 32'b00000100010000000000000011101111;
ROM[18039] <= 32'b00000000000000011010001110000011;
ROM[18040] <= 32'b00000000011100010010000000100011;
ROM[18041] <= 32'b00000000010000010000000100010011;
ROM[18042] <= 32'b00000000010000011010001110000011;
ROM[18043] <= 32'b00000000011100010010000000100011;
ROM[18044] <= 32'b00000000010000010000000100010011;
ROM[18045] <= 32'b11111111110000010000000100010011;
ROM[18046] <= 32'b00000000000000010010001110000011;
ROM[18047] <= 32'b11111111110000010000000100010011;
ROM[18048] <= 32'b00000000000000010010010000000011;
ROM[18049] <= 32'b00000000011101000000001110110011;
ROM[18050] <= 32'b00000000011100010010000000100011;
ROM[18051] <= 32'b00000000010000010000000100010011;
ROM[18052] <= 32'b11111111110000010000000100010011;
ROM[18053] <= 32'b00000000000000010010001110000011;
ROM[18054] <= 32'b00000000011100011010000000100011;
ROM[18055] <= 32'b00000000010000011010001110000011;
ROM[18056] <= 32'b00000000011100010010000000100011;
ROM[18057] <= 32'b00000000010000010000000100010011;
ROM[18058] <= 32'b00000000010000011010001110000011;
ROM[18059] <= 32'b00000000011100010010000000100011;
ROM[18060] <= 32'b00000000010000010000000100010011;
ROM[18061] <= 32'b11111111110000010000000100010011;
ROM[18062] <= 32'b00000000000000010010001110000011;
ROM[18063] <= 32'b11111111110000010000000100010011;
ROM[18064] <= 32'b00000000000000010010010000000011;
ROM[18065] <= 32'b00000000011101000000001110110011;
ROM[18066] <= 32'b00000000011100010010000000100011;
ROM[18067] <= 32'b00000000010000010000000100010011;
ROM[18068] <= 32'b11111111110000010000000100010011;
ROM[18069] <= 32'b00000000000000010010001110000011;
ROM[18070] <= 32'b00000000011100011010001000100011;
ROM[18071] <= 32'b00000000100000011010001110000011;
ROM[18072] <= 32'b00000000011100010010000000100011;
ROM[18073] <= 32'b00000000010000010000000100010011;
ROM[18074] <= 32'b00000000010000000000001110010011;
ROM[18075] <= 32'b00000000011100010010000000100011;
ROM[18076] <= 32'b00000000010000010000000100010011;
ROM[18077] <= 32'b11111111110000010000000100010011;
ROM[18078] <= 32'b00000000000000010010001110000011;
ROM[18079] <= 32'b11111111110000010000000100010011;
ROM[18080] <= 32'b00000000000000010010010000000011;
ROM[18081] <= 32'b00000000011101000000001110110011;
ROM[18082] <= 32'b00000000011100010010000000100011;
ROM[18083] <= 32'b00000000010000010000000100010011;
ROM[18084] <= 32'b11111111110000010000000100010011;
ROM[18085] <= 32'b00000000000000010010001110000011;
ROM[18086] <= 32'b00000000011100011010010000100011;
ROM[18087] <= 32'b11011111000111111111000011101111;
ROM[18088] <= 32'b00000000000000011010001110000011;
ROM[18089] <= 32'b00000000011100010010000000100011;
ROM[18090] <= 32'b00000000010000010000000100010011;
ROM[18091] <= 32'b00000001010000000000001110010011;
ROM[18092] <= 32'b01000000011100011000001110110011;
ROM[18093] <= 32'b00000000000000111010000010000011;
ROM[18094] <= 32'b11111111110000010000000100010011;
ROM[18095] <= 32'b00000000000000010010001110000011;
ROM[18096] <= 32'b00000000011100100010000000100011;
ROM[18097] <= 32'b00000000010000100000000100010011;
ROM[18098] <= 32'b00000001010000000000001110010011;
ROM[18099] <= 32'b01000000011100011000001110110011;
ROM[18100] <= 32'b00000000010000111010000110000011;
ROM[18101] <= 32'b00000000100000111010001000000011;
ROM[18102] <= 32'b00000000110000111010001010000011;
ROM[18103] <= 32'b00000001000000111010001100000011;
ROM[18104] <= 32'b00000000000000001000000011100111;
ROM[18105] <= 32'b00000000000000100010001110000011;
ROM[18106] <= 32'b00000000011100010010000000100011;
ROM[18107] <= 32'b00000000010000010000000100010011;
ROM[18108] <= 32'b00000000000000000000001110010011;
ROM[18109] <= 32'b00000000011100010010000000100011;
ROM[18110] <= 32'b00000000010000010000000100010011;
ROM[18111] <= 32'b11111111110000010000000100010011;
ROM[18112] <= 32'b00000000000000010010001110000011;
ROM[18113] <= 32'b11111111110000010000000100010011;
ROM[18114] <= 32'b00000000000000010010010000000011;
ROM[18115] <= 32'b00000000011101000010001110110011;
ROM[18116] <= 32'b00000000011100010010000000100011;
ROM[18117] <= 32'b00000000010000010000000100010011;
ROM[18118] <= 32'b11111111110000010000000100010011;
ROM[18119] <= 32'b00000000000000010010001110000011;
ROM[18120] <= 32'b00000000000000111000101001100011;
ROM[18121] <= 32'b00000000000000010010001110110111;
ROM[18122] <= 32'b10110011100000111000001110010011;
ROM[18123] <= 32'b00000000111000111000001110110011;
ROM[18124] <= 32'b00000000000000111000000011100111;
ROM[18125] <= 32'b00000011000000000000000011101111;
ROM[18126] <= 32'b00000000000000100010001110000011;
ROM[18127] <= 32'b00000000011100010010000000100011;
ROM[18128] <= 32'b00000000010000010000000100010011;
ROM[18129] <= 32'b11111111110000010000000100010011;
ROM[18130] <= 32'b00000000000000010010001110000011;
ROM[18131] <= 32'b01000000011100000000001110110011;
ROM[18132] <= 32'b00000000011100010010000000100011;
ROM[18133] <= 32'b00000000010000010000000100010011;
ROM[18134] <= 32'b11111111110000010000000100010011;
ROM[18135] <= 32'b00000000000000010010001110000011;
ROM[18136] <= 32'b00000000011100100010000000100011;
ROM[18137] <= 32'b00000000000000100010001110000011;
ROM[18138] <= 32'b00000000011100010010000000100011;
ROM[18139] <= 32'b00000000010000010000000100010011;
ROM[18140] <= 32'b00000001010000000000001110010011;
ROM[18141] <= 32'b01000000011100011000001110110011;
ROM[18142] <= 32'b00000000000000111010000010000011;
ROM[18143] <= 32'b11111111110000010000000100010011;
ROM[18144] <= 32'b00000000000000010010001110000011;
ROM[18145] <= 32'b00000000011100100010000000100011;
ROM[18146] <= 32'b00000000010000100000000100010011;
ROM[18147] <= 32'b00000001010000000000001110010011;
ROM[18148] <= 32'b01000000011100011000001110110011;
ROM[18149] <= 32'b00000000010000111010000110000011;
ROM[18150] <= 32'b00000000100000111010001000000011;
ROM[18151] <= 32'b00000000110000111010001010000011;
ROM[18152] <= 32'b00000001000000111010001100000011;
ROM[18153] <= 32'b00000000000000001000000011100111;
ROM[18154] <= 32'b00000000000000010010000000100011;
ROM[18155] <= 32'b00000000010000010000000100010011;
ROM[18156] <= 32'b00000000000000010010000000100011;
ROM[18157] <= 32'b00000000010000010000000100010011;
ROM[18158] <= 32'b00000000000000010010000000100011;
ROM[18159] <= 32'b00000000010000010000000100010011;
ROM[18160] <= 32'b00000000010000100010001110000011;
ROM[18161] <= 32'b00000000011100010010000000100011;
ROM[18162] <= 32'b00000000010000010000000100010011;
ROM[18163] <= 32'b00000000000000000000001110010011;
ROM[18164] <= 32'b00000000011100010010000000100011;
ROM[18165] <= 32'b00000000010000010000000100010011;
ROM[18166] <= 32'b11111111110000010000000100010011;
ROM[18167] <= 32'b00000000000000010010001110000011;
ROM[18168] <= 32'b11111111110000010000000100010011;
ROM[18169] <= 32'b00000000000000010010010000000011;
ROM[18170] <= 32'b00000000011101000010010010110011;
ROM[18171] <= 32'b00000000100000111010010100110011;
ROM[18172] <= 32'b00000000101001001000001110110011;
ROM[18173] <= 32'b00000000000100111000001110010011;
ROM[18174] <= 32'b00000000000100111111001110010011;
ROM[18175] <= 32'b00000000011100010010000000100011;
ROM[18176] <= 32'b00000000010000010000000100010011;
ROM[18177] <= 32'b11111111110000010000000100010011;
ROM[18178] <= 32'b00000000000000010010001110000011;
ROM[18179] <= 32'b00000000000000111000101001100011;
ROM[18180] <= 32'b00000000000000010010001110110111;
ROM[18181] <= 32'b11000010010000111000001110010011;
ROM[18182] <= 32'b00000000111000111000001110110011;
ROM[18183] <= 32'b00000000000000111000000011100111;
ROM[18184] <= 32'b00000101110000000000000011101111;
ROM[18185] <= 32'b00000000000100000000001110010011;
ROM[18186] <= 32'b00000000011100010010000000100011;
ROM[18187] <= 32'b00000000010000010000000100010011;
ROM[18188] <= 32'b11111111110000010000000100010011;
ROM[18189] <= 32'b00000000000000010010001110000011;
ROM[18190] <= 32'b01000000011100000000001110110011;
ROM[18191] <= 32'b00000000011100010010000000100011;
ROM[18192] <= 32'b00000000010000010000000100010011;
ROM[18193] <= 32'b00000001010000000000001110010011;
ROM[18194] <= 32'b01000000011100011000001110110011;
ROM[18195] <= 32'b00000000000000111010000010000011;
ROM[18196] <= 32'b11111111110000010000000100010011;
ROM[18197] <= 32'b00000000000000010010001110000011;
ROM[18198] <= 32'b00000000011100100010000000100011;
ROM[18199] <= 32'b00000000010000100000000100010011;
ROM[18200] <= 32'b00000001010000000000001110010011;
ROM[18201] <= 32'b01000000011100011000001110110011;
ROM[18202] <= 32'b00000000010000111010000110000011;
ROM[18203] <= 32'b00000000100000111010001000000011;
ROM[18204] <= 32'b00000000110000111010001010000011;
ROM[18205] <= 32'b00000001000000111010001100000011;
ROM[18206] <= 32'b00000000000000001000000011100111;
ROM[18207] <= 32'b00000000000000100010001110000011;
ROM[18208] <= 32'b00000000011100010010000000100011;
ROM[18209] <= 32'b00000000010000010000000100010011;
ROM[18210] <= 32'b00000000000000000000001110010011;
ROM[18211] <= 32'b00000000011100010010000000100011;
ROM[18212] <= 32'b00000000010000010000000100010011;
ROM[18213] <= 32'b11111111110000010000000100010011;
ROM[18214] <= 32'b00000000000000010010001110000011;
ROM[18215] <= 32'b11111111110000010000000100010011;
ROM[18216] <= 32'b00000000000000010010010000000011;
ROM[18217] <= 32'b00000000011101000010001110110011;
ROM[18218] <= 32'b00000000011100010010000000100011;
ROM[18219] <= 32'b00000000010000010000000100010011;
ROM[18220] <= 32'b00000000010000100010001110000011;
ROM[18221] <= 32'b00000000011100010010000000100011;
ROM[18222] <= 32'b00000000010000010000000100010011;
ROM[18223] <= 32'b00000000000000000000001110010011;
ROM[18224] <= 32'b00000000011100010010000000100011;
ROM[18225] <= 32'b00000000010000010000000100010011;
ROM[18226] <= 32'b11111111110000010000000100010011;
ROM[18227] <= 32'b00000000000000010010001110000011;
ROM[18228] <= 32'b11111111110000010000000100010011;
ROM[18229] <= 32'b00000000000000010010010000000011;
ROM[18230] <= 32'b00000000011101000010001110110011;
ROM[18231] <= 32'b00000000011100010010000000100011;
ROM[18232] <= 32'b00000000010000010000000100010011;
ROM[18233] <= 32'b11111111110000010000000100010011;
ROM[18234] <= 32'b00000000000000010010001110000011;
ROM[18235] <= 32'b11111111110000010000000100010011;
ROM[18236] <= 32'b00000000000000010010010000000011;
ROM[18237] <= 32'b00000000011101000010010010110011;
ROM[18238] <= 32'b00000000100000111010010100110011;
ROM[18239] <= 32'b00000000101001001000001110110011;
ROM[18240] <= 32'b00000000000100111000001110010011;
ROM[18241] <= 32'b00000000000100111111001110010011;
ROM[18242] <= 32'b00000000011100010010000000100011;
ROM[18243] <= 32'b00000000010000010000000100010011;
ROM[18244] <= 32'b11111111110000010000000100010011;
ROM[18245] <= 32'b00000000000000010010001110000011;
ROM[18246] <= 32'b01000000011100000000001110110011;
ROM[18247] <= 32'b00000000000100111000001110010011;
ROM[18248] <= 32'b00000000011100010010000000100011;
ROM[18249] <= 32'b00000000010000010000000100010011;
ROM[18250] <= 32'b11111111110000010000000100010011;
ROM[18251] <= 32'b00000000000000010010001110000011;
ROM[18252] <= 32'b00000000011100011010001000100011;
ROM[18253] <= 32'b00000000000000100010001110000011;
ROM[18254] <= 32'b00000000011100010010000000100011;
ROM[18255] <= 32'b00000000010000010000000100010011;
ROM[18256] <= 32'b00000000000000010010001110110111;
ROM[18257] <= 32'b11011000110000111000001110010011;
ROM[18258] <= 32'b00000000111000111000001110110011;
ROM[18259] <= 32'b00000000011100010010000000100011;
ROM[18260] <= 32'b00000000010000010000000100010011;
ROM[18261] <= 32'b00000000001100010010000000100011;
ROM[18262] <= 32'b00000000010000010000000100010011;
ROM[18263] <= 32'b00000000010000010010000000100011;
ROM[18264] <= 32'b00000000010000010000000100010011;
ROM[18265] <= 32'b00000000010100010010000000100011;
ROM[18266] <= 32'b00000000010000010000000100010011;
ROM[18267] <= 32'b00000000011000010010000000100011;
ROM[18268] <= 32'b00000000010000010000000100010011;
ROM[18269] <= 32'b00000001010000000000001110010011;
ROM[18270] <= 32'b00000000010000111000001110010011;
ROM[18271] <= 32'b01000000011100010000001110110011;
ROM[18272] <= 32'b00000000011100000000001000110011;
ROM[18273] <= 32'b00000000001000000000000110110011;
ROM[18274] <= 32'b11010101110111111111000011101111;
ROM[18275] <= 32'b11111111110000010000000100010011;
ROM[18276] <= 32'b00000000000000010010001110000011;
ROM[18277] <= 32'b00000000011100100010000000100011;
ROM[18278] <= 32'b00000000010000100010001110000011;
ROM[18279] <= 32'b00000000011100010010000000100011;
ROM[18280] <= 32'b00000000010000010000000100010011;
ROM[18281] <= 32'b00000000000000010010001110110111;
ROM[18282] <= 32'b11011111000000111000001110010011;
ROM[18283] <= 32'b00000000111000111000001110110011;
ROM[18284] <= 32'b00000000011100010010000000100011;
ROM[18285] <= 32'b00000000010000010000000100010011;
ROM[18286] <= 32'b00000000001100010010000000100011;
ROM[18287] <= 32'b00000000010000010000000100010011;
ROM[18288] <= 32'b00000000010000010010000000100011;
ROM[18289] <= 32'b00000000010000010000000100010011;
ROM[18290] <= 32'b00000000010100010010000000100011;
ROM[18291] <= 32'b00000000010000010000000100010011;
ROM[18292] <= 32'b00000000011000010010000000100011;
ROM[18293] <= 32'b00000000010000010000000100010011;
ROM[18294] <= 32'b00000001010000000000001110010011;
ROM[18295] <= 32'b00000000010000111000001110010011;
ROM[18296] <= 32'b01000000011100010000001110110011;
ROM[18297] <= 32'b00000000011100000000001000110011;
ROM[18298] <= 32'b00000000001000000000000110110011;
ROM[18299] <= 32'b11001111100111111111000011101111;
ROM[18300] <= 32'b11111111110000010000000100010011;
ROM[18301] <= 32'b00000000000000010010001110000011;
ROM[18302] <= 32'b00000000011100100010001000100011;
ROM[18303] <= 32'b00000000000000000000001110010011;
ROM[18304] <= 32'b00000000011100010010000000100011;
ROM[18305] <= 32'b00000000010000010000000100010011;
ROM[18306] <= 32'b11111111110000010000000100010011;
ROM[18307] <= 32'b00000000000000010010001110000011;
ROM[18308] <= 32'b00000000011100011010000000100011;
ROM[18309] <= 32'b00000000010000100010001110000011;
ROM[18310] <= 32'b00000000011100010010000000100011;
ROM[18311] <= 32'b00000000010000010000000100010011;
ROM[18312] <= 32'b00000000000000100010001110000011;
ROM[18313] <= 32'b00000000011100010010000000100011;
ROM[18314] <= 32'b00000000010000010000000100010011;
ROM[18315] <= 32'b11111111110000010000000100010011;
ROM[18316] <= 32'b00000000000000010010001110000011;
ROM[18317] <= 32'b11111111110000010000000100010011;
ROM[18318] <= 32'b00000000000000010010010000000011;
ROM[18319] <= 32'b00000000100000111010001110110011;
ROM[18320] <= 32'b00000000011100010010000000100011;
ROM[18321] <= 32'b00000000010000010000000100010011;
ROM[18322] <= 32'b11111111110000010000000100010011;
ROM[18323] <= 32'b00000000000000010010001110000011;
ROM[18324] <= 32'b01000000011100000000001110110011;
ROM[18325] <= 32'b00000000000100111000001110010011;
ROM[18326] <= 32'b00000000011100010010000000100011;
ROM[18327] <= 32'b00000000010000010000000100010011;
ROM[18328] <= 32'b11111111110000010000000100010011;
ROM[18329] <= 32'b00000000000000010010001110000011;
ROM[18330] <= 32'b00000000011100011010010000100011;
ROM[18331] <= 32'b00000000100000011010001110000011;
ROM[18332] <= 32'b00000000011100010010000000100011;
ROM[18333] <= 32'b00000000010000010000000100010011;
ROM[18334] <= 32'b11111111110000010000000100010011;
ROM[18335] <= 32'b00000000000000010010001110000011;
ROM[18336] <= 32'b01000000011100000000001110110011;
ROM[18337] <= 32'b00000000000100111000001110010011;
ROM[18338] <= 32'b00000000011100010010000000100011;
ROM[18339] <= 32'b00000000010000010000000100010011;
ROM[18340] <= 32'b11111111110000010000000100010011;
ROM[18341] <= 32'b00000000000000010010001110000011;
ROM[18342] <= 32'b00000000000000111000101001100011;
ROM[18343] <= 32'b00000000000000010010001110110111;
ROM[18344] <= 32'b11111000100000111000001110010011;
ROM[18345] <= 32'b00000000111000111000001110110011;
ROM[18346] <= 32'b00000000000000111000000011100111;
ROM[18347] <= 32'b00000000000000100010001110000011;
ROM[18348] <= 32'b00000000011100010010000000100011;
ROM[18349] <= 32'b00000000010000010000000100010011;
ROM[18350] <= 32'b00000000010000100010001110000011;
ROM[18351] <= 32'b00000000011100010010000000100011;
ROM[18352] <= 32'b00000000010000010000000100010011;
ROM[18353] <= 32'b11111111110000010000000100010011;
ROM[18354] <= 32'b00000000000000010010001110000011;
ROM[18355] <= 32'b11111111110000010000000100010011;
ROM[18356] <= 32'b00000000000000010010010000000011;
ROM[18357] <= 32'b01000000011101000000001110110011;
ROM[18358] <= 32'b00000000011100010010000000100011;
ROM[18359] <= 32'b00000000010000010000000100010011;
ROM[18360] <= 32'b11111111110000010000000100010011;
ROM[18361] <= 32'b00000000000000010010001110000011;
ROM[18362] <= 32'b00000000011100100010000000100011;
ROM[18363] <= 32'b00000000000000011010001110000011;
ROM[18364] <= 32'b00000000011100010010000000100011;
ROM[18365] <= 32'b00000000010000010000000100010011;
ROM[18366] <= 32'b00000000000100000000001110010011;
ROM[18367] <= 32'b00000000011100010010000000100011;
ROM[18368] <= 32'b00000000010000010000000100010011;
ROM[18369] <= 32'b11111111110000010000000100010011;
ROM[18370] <= 32'b00000000000000010010001110000011;
ROM[18371] <= 32'b11111111110000010000000100010011;
ROM[18372] <= 32'b00000000000000010010010000000011;
ROM[18373] <= 32'b00000000011101000000001110110011;
ROM[18374] <= 32'b00000000011100010010000000100011;
ROM[18375] <= 32'b00000000010000010000000100010011;
ROM[18376] <= 32'b11111111110000010000000100010011;
ROM[18377] <= 32'b00000000000000010010001110000011;
ROM[18378] <= 32'b00000000011100011010000000100011;
ROM[18379] <= 32'b00000000010000100010001110000011;
ROM[18380] <= 32'b00000000011100010010000000100011;
ROM[18381] <= 32'b00000000010000010000000100010011;
ROM[18382] <= 32'b00000000000000100010001110000011;
ROM[18383] <= 32'b00000000011100010010000000100011;
ROM[18384] <= 32'b00000000010000010000000100010011;
ROM[18385] <= 32'b11111111110000010000000100010011;
ROM[18386] <= 32'b00000000000000010010001110000011;
ROM[18387] <= 32'b11111111110000010000000100010011;
ROM[18388] <= 32'b00000000000000010010010000000011;
ROM[18389] <= 32'b00000000100000111010001110110011;
ROM[18390] <= 32'b00000000011100010010000000100011;
ROM[18391] <= 32'b00000000010000010000000100010011;
ROM[18392] <= 32'b11111111110000010000000100010011;
ROM[18393] <= 32'b00000000000000010010001110000011;
ROM[18394] <= 32'b01000000011100000000001110110011;
ROM[18395] <= 32'b00000000000100111000001110010011;
ROM[18396] <= 32'b00000000011100010010000000100011;
ROM[18397] <= 32'b00000000010000010000000100010011;
ROM[18398] <= 32'b11111111110000010000000100010011;
ROM[18399] <= 32'b00000000000000010010001110000011;
ROM[18400] <= 32'b00000000011100011010010000100011;
ROM[18401] <= 32'b11101110100111111111000011101111;
ROM[18402] <= 32'b00000000010000011010001110000011;
ROM[18403] <= 32'b00000000011100010010000000100011;
ROM[18404] <= 32'b00000000010000010000000100010011;
ROM[18405] <= 32'b11111111110000010000000100010011;
ROM[18406] <= 32'b00000000000000010010001110000011;
ROM[18407] <= 32'b00000000000000111000101001100011;
ROM[18408] <= 32'b00000000000000010010001110110111;
ROM[18409] <= 32'b11111011010000111000001110010011;
ROM[18410] <= 32'b00000000111000111000001110110011;
ROM[18411] <= 32'b00000000000000111000000011100111;
ROM[18412] <= 32'b00000011000000000000000011101111;
ROM[18413] <= 32'b00000000000000011010001110000011;
ROM[18414] <= 32'b00000000011100010010000000100011;
ROM[18415] <= 32'b00000000010000010000000100010011;
ROM[18416] <= 32'b11111111110000010000000100010011;
ROM[18417] <= 32'b00000000000000010010001110000011;
ROM[18418] <= 32'b01000000011100000000001110110011;
ROM[18419] <= 32'b00000000011100010010000000100011;
ROM[18420] <= 32'b00000000010000010000000100010011;
ROM[18421] <= 32'b11111111110000010000000100010011;
ROM[18422] <= 32'b00000000000000010010001110000011;
ROM[18423] <= 32'b00000000011100011010000000100011;
ROM[18424] <= 32'b00000000000000011010001110000011;
ROM[18425] <= 32'b00000000011100010010000000100011;
ROM[18426] <= 32'b00000000010000010000000100010011;
ROM[18427] <= 32'b00000001010000000000001110010011;
ROM[18428] <= 32'b01000000011100011000001110110011;
ROM[18429] <= 32'b00000000000000111010000010000011;
ROM[18430] <= 32'b11111111110000010000000100010011;
ROM[18431] <= 32'b00000000000000010010001110000011;
ROM[18432] <= 32'b00000000011100100010000000100011;
ROM[18433] <= 32'b00000000010000100000000100010011;
ROM[18434] <= 32'b00000001010000000000001110010011;
ROM[18435] <= 32'b01000000011100011000001110110011;
ROM[18436] <= 32'b00000000010000111010000110000011;
ROM[18437] <= 32'b00000000100000111010001000000011;
ROM[18438] <= 32'b00000000110000111010001010000011;
ROM[18439] <= 32'b00000001000000111010001100000011;
ROM[18440] <= 32'b00000000000000001000000011100111;
ROM[18441] <= 32'b00000000000000010010000000100011;
ROM[18442] <= 32'b00000000010000010000000100010011;
ROM[18443] <= 32'b00000000000000010010000000100011;
ROM[18444] <= 32'b00000000010000010000000100010011;
ROM[18445] <= 32'b00000000000000010010000000100011;
ROM[18446] <= 32'b00000000010000010000000100010011;
ROM[18447] <= 32'b00000000000000010010000000100011;
ROM[18448] <= 32'b00000000010000010000000100010011;
ROM[18449] <= 32'b00000000000000100010001110000011;
ROM[18450] <= 32'b00000000011100010010000000100011;
ROM[18451] <= 32'b00000000010000010000000100010011;
ROM[18452] <= 32'b00000000000000000000001110010011;
ROM[18453] <= 32'b00000000011100010010000000100011;
ROM[18454] <= 32'b00000000010000010000000100010011;
ROM[18455] <= 32'b11111111110000010000000100010011;
ROM[18456] <= 32'b00000000000000010010001110000011;
ROM[18457] <= 32'b11111111110000010000000100010011;
ROM[18458] <= 32'b00000000000000010010010000000011;
ROM[18459] <= 32'b00000000011101000010001110110011;
ROM[18460] <= 32'b00000000011100010010000000100011;
ROM[18461] <= 32'b00000000010000010000000100010011;
ROM[18462] <= 32'b11111111110000010000000100010011;
ROM[18463] <= 32'b00000000000000010010001110000011;
ROM[18464] <= 32'b00000000000000111000101001100011;
ROM[18465] <= 32'b00000000000000010010001110110111;
ROM[18466] <= 32'b00001001100000111000001110010011;
ROM[18467] <= 32'b00000000111000111000001110110011;
ROM[18468] <= 32'b00000000000000111000000011100111;
ROM[18469] <= 32'b00110000010100000000000011101111;
ROM[18470] <= 32'b00000001110000000000001110010011;
ROM[18471] <= 32'b00000000011100010010000000100011;
ROM[18472] <= 32'b00000000010000010000000100010011;
ROM[18473] <= 32'b00000000000000010010001110110111;
ROM[18474] <= 32'b00001111000000111000001110010011;
ROM[18475] <= 32'b00000000111000111000001110110011;
ROM[18476] <= 32'b00000000011100010010000000100011;
ROM[18477] <= 32'b00000000010000010000000100010011;
ROM[18478] <= 32'b00000000001100010010000000100011;
ROM[18479] <= 32'b00000000010000010000000100010011;
ROM[18480] <= 32'b00000000010000010010000000100011;
ROM[18481] <= 32'b00000000010000010000000100010011;
ROM[18482] <= 32'b00000000010100010010000000100011;
ROM[18483] <= 32'b00000000010000010000000100010011;
ROM[18484] <= 32'b00000000011000010010000000100011;
ROM[18485] <= 32'b00000000010000010000000100010011;
ROM[18486] <= 32'b00000001010000000000001110010011;
ROM[18487] <= 32'b00000000010000111000001110010011;
ROM[18488] <= 32'b01000000011100010000001110110011;
ROM[18489] <= 32'b00000000011100000000001000110011;
ROM[18490] <= 32'b00000000001000000000000110110011;
ROM[18491] <= 32'b01100101000000010111000011101111;
ROM[18492] <= 32'b00000111001100000000001110010011;
ROM[18493] <= 32'b00000000011100010010000000100011;
ROM[18494] <= 32'b00000000010000010000000100010011;
ROM[18495] <= 32'b00000000000000010010001110110111;
ROM[18496] <= 32'b00010100100000111000001110010011;
ROM[18497] <= 32'b00000000111000111000001110110011;
ROM[18498] <= 32'b00000000011100010010000000100011;
ROM[18499] <= 32'b00000000010000010000000100010011;
ROM[18500] <= 32'b00000000001100010010000000100011;
ROM[18501] <= 32'b00000000010000010000000100010011;
ROM[18502] <= 32'b00000000010000010010000000100011;
ROM[18503] <= 32'b00000000010000010000000100010011;
ROM[18504] <= 32'b00000000010100010010000000100011;
ROM[18505] <= 32'b00000000010000010000000100010011;
ROM[18506] <= 32'b00000000011000010010000000100011;
ROM[18507] <= 32'b00000000010000010000000100010011;
ROM[18508] <= 32'b00000001010000000000001110010011;
ROM[18509] <= 32'b00000000100000111000001110010011;
ROM[18510] <= 32'b01000000011100010000001110110011;
ROM[18511] <= 32'b00000000011100000000001000110011;
ROM[18512] <= 32'b00000000001000000000000110110011;
ROM[18513] <= 32'b00100110100100010111000011101111;
ROM[18514] <= 32'b00000111000100000000001110010011;
ROM[18515] <= 32'b00000000011100010010000000100011;
ROM[18516] <= 32'b00000000010000010000000100010011;
ROM[18517] <= 32'b00000000000000010010001110110111;
ROM[18518] <= 32'b00011010000000111000001110010011;
ROM[18519] <= 32'b00000000111000111000001110110011;
ROM[18520] <= 32'b00000000011100010010000000100011;
ROM[18521] <= 32'b00000000010000010000000100010011;
ROM[18522] <= 32'b00000000001100010010000000100011;
ROM[18523] <= 32'b00000000010000010000000100010011;
ROM[18524] <= 32'b00000000010000010010000000100011;
ROM[18525] <= 32'b00000000010000010000000100010011;
ROM[18526] <= 32'b00000000010100010010000000100011;
ROM[18527] <= 32'b00000000010000010000000100010011;
ROM[18528] <= 32'b00000000011000010010000000100011;
ROM[18529] <= 32'b00000000010000010000000100010011;
ROM[18530] <= 32'b00000001010000000000001110010011;
ROM[18531] <= 32'b00000000100000111000001110010011;
ROM[18532] <= 32'b01000000011100010000001110110011;
ROM[18533] <= 32'b00000000011100000000001000110011;
ROM[18534] <= 32'b00000000001000000000000110110011;
ROM[18535] <= 32'b00100001000100010111000011101111;
ROM[18536] <= 32'b00000111001000000000001110010011;
ROM[18537] <= 32'b00000000011100010010000000100011;
ROM[18538] <= 32'b00000000010000010000000100010011;
ROM[18539] <= 32'b00000000000000010010001110110111;
ROM[18540] <= 32'b00011111100000111000001110010011;
ROM[18541] <= 32'b00000000111000111000001110110011;
ROM[18542] <= 32'b00000000011100010010000000100011;
ROM[18543] <= 32'b00000000010000010000000100010011;
ROM[18544] <= 32'b00000000001100010010000000100011;
ROM[18545] <= 32'b00000000010000010000000100010011;
ROM[18546] <= 32'b00000000010000010010000000100011;
ROM[18547] <= 32'b00000000010000010000000100010011;
ROM[18548] <= 32'b00000000010100010010000000100011;
ROM[18549] <= 32'b00000000010000010000000100010011;
ROM[18550] <= 32'b00000000011000010010000000100011;
ROM[18551] <= 32'b00000000010000010000000100010011;
ROM[18552] <= 32'b00000001010000000000001110010011;
ROM[18553] <= 32'b00000000100000111000001110010011;
ROM[18554] <= 32'b01000000011100010000001110110011;
ROM[18555] <= 32'b00000000011100000000001000110011;
ROM[18556] <= 32'b00000000001000000000000110110011;
ROM[18557] <= 32'b00011011100100010111000011101111;
ROM[18558] <= 32'b00000111010000000000001110010011;
ROM[18559] <= 32'b00000000011100010010000000100011;
ROM[18560] <= 32'b00000000010000010000000100010011;
ROM[18561] <= 32'b00000000000000010010001110110111;
ROM[18562] <= 32'b00100101000000111000001110010011;
ROM[18563] <= 32'b00000000111000111000001110110011;
ROM[18564] <= 32'b00000000011100010010000000100011;
ROM[18565] <= 32'b00000000010000010000000100010011;
ROM[18566] <= 32'b00000000001100010010000000100011;
ROM[18567] <= 32'b00000000010000010000000100010011;
ROM[18568] <= 32'b00000000010000010010000000100011;
ROM[18569] <= 32'b00000000010000010000000100010011;
ROM[18570] <= 32'b00000000010100010010000000100011;
ROM[18571] <= 32'b00000000010000010000000100010011;
ROM[18572] <= 32'b00000000011000010010000000100011;
ROM[18573] <= 32'b00000000010000010000000100010011;
ROM[18574] <= 32'b00000001010000000000001110010011;
ROM[18575] <= 32'b00000000100000111000001110010011;
ROM[18576] <= 32'b01000000011100010000001110110011;
ROM[18577] <= 32'b00000000011100000000001000110011;
ROM[18578] <= 32'b00000000001000000000000110110011;
ROM[18579] <= 32'b00010110000100010111000011101111;
ROM[18580] <= 32'b00000011101000000000001110010011;
ROM[18581] <= 32'b00000000011100010010000000100011;
ROM[18582] <= 32'b00000000010000010000000100010011;
ROM[18583] <= 32'b00000000000000010010001110110111;
ROM[18584] <= 32'b00101010100000111000001110010011;
ROM[18585] <= 32'b00000000111000111000001110110011;
ROM[18586] <= 32'b00000000011100010010000000100011;
ROM[18587] <= 32'b00000000010000010000000100010011;
ROM[18588] <= 32'b00000000001100010010000000100011;
ROM[18589] <= 32'b00000000010000010000000100010011;
ROM[18590] <= 32'b00000000010000010010000000100011;
ROM[18591] <= 32'b00000000010000010000000100010011;
ROM[18592] <= 32'b00000000010100010010000000100011;
ROM[18593] <= 32'b00000000010000010000000100010011;
ROM[18594] <= 32'b00000000011000010010000000100011;
ROM[18595] <= 32'b00000000010000010000000100010011;
ROM[18596] <= 32'b00000001010000000000001110010011;
ROM[18597] <= 32'b00000000100000111000001110010011;
ROM[18598] <= 32'b01000000011100010000001110110011;
ROM[18599] <= 32'b00000000011100000000001000110011;
ROM[18600] <= 32'b00000000001000000000000110110011;
ROM[18601] <= 32'b00010000100100010111000011101111;
ROM[18602] <= 32'b00000010000000000000001110010011;
ROM[18603] <= 32'b00000000011100010010000000100011;
ROM[18604] <= 32'b00000000010000010000000100010011;
ROM[18605] <= 32'b00000000000000010010001110110111;
ROM[18606] <= 32'b00110000000000111000001110010011;
ROM[18607] <= 32'b00000000111000111000001110110011;
ROM[18608] <= 32'b00000000011100010010000000100011;
ROM[18609] <= 32'b00000000010000010000000100010011;
ROM[18610] <= 32'b00000000001100010010000000100011;
ROM[18611] <= 32'b00000000010000010000000100010011;
ROM[18612] <= 32'b00000000010000010010000000100011;
ROM[18613] <= 32'b00000000010000010000000100010011;
ROM[18614] <= 32'b00000000010100010010000000100011;
ROM[18615] <= 32'b00000000010000010000000100010011;
ROM[18616] <= 32'b00000000011000010010000000100011;
ROM[18617] <= 32'b00000000010000010000000100010011;
ROM[18618] <= 32'b00000001010000000000001110010011;
ROM[18619] <= 32'b00000000100000111000001110010011;
ROM[18620] <= 32'b01000000011100010000001110110011;
ROM[18621] <= 32'b00000000011100000000001000110011;
ROM[18622] <= 32'b00000000001000000000000110110011;
ROM[18623] <= 32'b00001011000100010111000011101111;
ROM[18624] <= 32'b00000110000100000000001110010011;
ROM[18625] <= 32'b00000000011100010010000000100011;
ROM[18626] <= 32'b00000000010000010000000100010011;
ROM[18627] <= 32'b00000000000000010010001110110111;
ROM[18628] <= 32'b00110101100000111000001110010011;
ROM[18629] <= 32'b00000000111000111000001110110011;
ROM[18630] <= 32'b00000000011100010010000000100011;
ROM[18631] <= 32'b00000000010000010000000100010011;
ROM[18632] <= 32'b00000000001100010010000000100011;
ROM[18633] <= 32'b00000000010000010000000100010011;
ROM[18634] <= 32'b00000000010000010010000000100011;
ROM[18635] <= 32'b00000000010000010000000100010011;
ROM[18636] <= 32'b00000000010100010010000000100011;
ROM[18637] <= 32'b00000000010000010000000100010011;
ROM[18638] <= 32'b00000000011000010010000000100011;
ROM[18639] <= 32'b00000000010000010000000100010011;
ROM[18640] <= 32'b00000001010000000000001110010011;
ROM[18641] <= 32'b00000000100000111000001110010011;
ROM[18642] <= 32'b01000000011100010000001110110011;
ROM[18643] <= 32'b00000000011100000000001000110011;
ROM[18644] <= 32'b00000000001000000000000110110011;
ROM[18645] <= 32'b00000101100100010111000011101111;
ROM[18646] <= 32'b00000111001000000000001110010011;
ROM[18647] <= 32'b00000000011100010010000000100011;
ROM[18648] <= 32'b00000000010000010000000100010011;
ROM[18649] <= 32'b00000000000000010010001110110111;
ROM[18650] <= 32'b00111011000000111000001110010011;
ROM[18651] <= 32'b00000000111000111000001110110011;
ROM[18652] <= 32'b00000000011100010010000000100011;
ROM[18653] <= 32'b00000000010000010000000100010011;
ROM[18654] <= 32'b00000000001100010010000000100011;
ROM[18655] <= 32'b00000000010000010000000100010011;
ROM[18656] <= 32'b00000000010000010010000000100011;
ROM[18657] <= 32'b00000000010000010000000100010011;
ROM[18658] <= 32'b00000000010100010010000000100011;
ROM[18659] <= 32'b00000000010000010000000100010011;
ROM[18660] <= 32'b00000000011000010010000000100011;
ROM[18661] <= 32'b00000000010000010000000100010011;
ROM[18662] <= 32'b00000001010000000000001110010011;
ROM[18663] <= 32'b00000000100000111000001110010011;
ROM[18664] <= 32'b01000000011100010000001110110011;
ROM[18665] <= 32'b00000000011100000000001000110011;
ROM[18666] <= 32'b00000000001000000000000110110011;
ROM[18667] <= 32'b00000000000100010111000011101111;
ROM[18668] <= 32'b00000110011100000000001110010011;
ROM[18669] <= 32'b00000000011100010010000000100011;
ROM[18670] <= 32'b00000000010000010000000100010011;
ROM[18671] <= 32'b00000000000000010010001110110111;
ROM[18672] <= 32'b01000000100000111000001110010011;
ROM[18673] <= 32'b00000000111000111000001110110011;
ROM[18674] <= 32'b00000000011100010010000000100011;
ROM[18675] <= 32'b00000000010000010000000100010011;
ROM[18676] <= 32'b00000000001100010010000000100011;
ROM[18677] <= 32'b00000000010000010000000100010011;
ROM[18678] <= 32'b00000000010000010010000000100011;
ROM[18679] <= 32'b00000000010000010000000100010011;
ROM[18680] <= 32'b00000000010100010010000000100011;
ROM[18681] <= 32'b00000000010000010000000100010011;
ROM[18682] <= 32'b00000000011000010010000000100011;
ROM[18683] <= 32'b00000000010000010000000100010011;
ROM[18684] <= 32'b00000001010000000000001110010011;
ROM[18685] <= 32'b00000000100000111000001110010011;
ROM[18686] <= 32'b01000000011100010000001110110011;
ROM[18687] <= 32'b00000000011100000000001000110011;
ROM[18688] <= 32'b00000000001000000000000110110011;
ROM[18689] <= 32'b01111010100000010111000011101111;
ROM[18690] <= 32'b00000111010100000000001110010011;
ROM[18691] <= 32'b00000000011100010010000000100011;
ROM[18692] <= 32'b00000000010000010000000100010011;
ROM[18693] <= 32'b00000000000000010010001110110111;
ROM[18694] <= 32'b01000110000000111000001110010011;
ROM[18695] <= 32'b00000000111000111000001110110011;
ROM[18696] <= 32'b00000000011100010010000000100011;
ROM[18697] <= 32'b00000000010000010000000100010011;
ROM[18698] <= 32'b00000000001100010010000000100011;
ROM[18699] <= 32'b00000000010000010000000100010011;
ROM[18700] <= 32'b00000000010000010010000000100011;
ROM[18701] <= 32'b00000000010000010000000100010011;
ROM[18702] <= 32'b00000000010100010010000000100011;
ROM[18703] <= 32'b00000000010000010000000100010011;
ROM[18704] <= 32'b00000000011000010010000000100011;
ROM[18705] <= 32'b00000000010000010000000100010011;
ROM[18706] <= 32'b00000001010000000000001110010011;
ROM[18707] <= 32'b00000000100000111000001110010011;
ROM[18708] <= 32'b01000000011100010000001110110011;
ROM[18709] <= 32'b00000000011100000000001000110011;
ROM[18710] <= 32'b00000000001000000000000110110011;
ROM[18711] <= 32'b01110101000000010111000011101111;
ROM[18712] <= 32'b00000110110100000000001110010011;
ROM[18713] <= 32'b00000000011100010010000000100011;
ROM[18714] <= 32'b00000000010000010000000100010011;
ROM[18715] <= 32'b00000000000000010010001110110111;
ROM[18716] <= 32'b01001011100000111000001110010011;
ROM[18717] <= 32'b00000000111000111000001110110011;
ROM[18718] <= 32'b00000000011100010010000000100011;
ROM[18719] <= 32'b00000000010000010000000100010011;
ROM[18720] <= 32'b00000000001100010010000000100011;
ROM[18721] <= 32'b00000000010000010000000100010011;
ROM[18722] <= 32'b00000000010000010010000000100011;
ROM[18723] <= 32'b00000000010000010000000100010011;
ROM[18724] <= 32'b00000000010100010010000000100011;
ROM[18725] <= 32'b00000000010000010000000100010011;
ROM[18726] <= 32'b00000000011000010010000000100011;
ROM[18727] <= 32'b00000000010000010000000100010011;
ROM[18728] <= 32'b00000001010000000000001110010011;
ROM[18729] <= 32'b00000000100000111000001110010011;
ROM[18730] <= 32'b01000000011100010000001110110011;
ROM[18731] <= 32'b00000000011100000000001000110011;
ROM[18732] <= 32'b00000000001000000000000110110011;
ROM[18733] <= 32'b01101111100000010111000011101111;
ROM[18734] <= 32'b00000110010100000000001110010011;
ROM[18735] <= 32'b00000000011100010010000000100011;
ROM[18736] <= 32'b00000000010000010000000100010011;
ROM[18737] <= 32'b00000000000000010010001110110111;
ROM[18738] <= 32'b01010001000000111000001110010011;
ROM[18739] <= 32'b00000000111000111000001110110011;
ROM[18740] <= 32'b00000000011100010010000000100011;
ROM[18741] <= 32'b00000000010000010000000100010011;
ROM[18742] <= 32'b00000000001100010010000000100011;
ROM[18743] <= 32'b00000000010000010000000100010011;
ROM[18744] <= 32'b00000000010000010010000000100011;
ROM[18745] <= 32'b00000000010000010000000100010011;
ROM[18746] <= 32'b00000000010100010010000000100011;
ROM[18747] <= 32'b00000000010000010000000100010011;
ROM[18748] <= 32'b00000000011000010010000000100011;
ROM[18749] <= 32'b00000000010000010000000100010011;
ROM[18750] <= 32'b00000001010000000000001110010011;
ROM[18751] <= 32'b00000000100000111000001110010011;
ROM[18752] <= 32'b01000000011100010000001110110011;
ROM[18753] <= 32'b00000000011100000000001000110011;
ROM[18754] <= 32'b00000000001000000000000110110011;
ROM[18755] <= 32'b01101010000000010111000011101111;
ROM[18756] <= 32'b00000110111000000000001110010011;
ROM[18757] <= 32'b00000000011100010010000000100011;
ROM[18758] <= 32'b00000000010000010000000100010011;
ROM[18759] <= 32'b00000000000000010010001110110111;
ROM[18760] <= 32'b01010110100000111000001110010011;
ROM[18761] <= 32'b00000000111000111000001110110011;
ROM[18762] <= 32'b00000000011100010010000000100011;
ROM[18763] <= 32'b00000000010000010000000100010011;
ROM[18764] <= 32'b00000000001100010010000000100011;
ROM[18765] <= 32'b00000000010000010000000100010011;
ROM[18766] <= 32'b00000000010000010010000000100011;
ROM[18767] <= 32'b00000000010000010000000100010011;
ROM[18768] <= 32'b00000000010100010010000000100011;
ROM[18769] <= 32'b00000000010000010000000100010011;
ROM[18770] <= 32'b00000000011000010010000000100011;
ROM[18771] <= 32'b00000000010000010000000100010011;
ROM[18772] <= 32'b00000001010000000000001110010011;
ROM[18773] <= 32'b00000000100000111000001110010011;
ROM[18774] <= 32'b01000000011100010000001110110011;
ROM[18775] <= 32'b00000000011100000000001000110011;
ROM[18776] <= 32'b00000000001000000000000110110011;
ROM[18777] <= 32'b01100100100000010111000011101111;
ROM[18778] <= 32'b00000111010000000000001110010011;
ROM[18779] <= 32'b00000000011100010010000000100011;
ROM[18780] <= 32'b00000000010000010000000100010011;
ROM[18781] <= 32'b00000000000000010010001110110111;
ROM[18782] <= 32'b01011100000000111000001110010011;
ROM[18783] <= 32'b00000000111000111000001110110011;
ROM[18784] <= 32'b00000000011100010010000000100011;
ROM[18785] <= 32'b00000000010000010000000100010011;
ROM[18786] <= 32'b00000000001100010010000000100011;
ROM[18787] <= 32'b00000000010000010000000100010011;
ROM[18788] <= 32'b00000000010000010010000000100011;
ROM[18789] <= 32'b00000000010000010000000100010011;
ROM[18790] <= 32'b00000000010100010010000000100011;
ROM[18791] <= 32'b00000000010000010000000100010011;
ROM[18792] <= 32'b00000000011000010010000000100011;
ROM[18793] <= 32'b00000000010000010000000100010011;
ROM[18794] <= 32'b00000001010000000000001110010011;
ROM[18795] <= 32'b00000000100000111000001110010011;
ROM[18796] <= 32'b01000000011100010000001110110011;
ROM[18797] <= 32'b00000000011100000000001000110011;
ROM[18798] <= 32'b00000000001000000000000110110011;
ROM[18799] <= 32'b01011111000000010111000011101111;
ROM[18800] <= 32'b00000010000000000000001110010011;
ROM[18801] <= 32'b00000000011100010010000000100011;
ROM[18802] <= 32'b00000000010000010000000100010011;
ROM[18803] <= 32'b00000000000000010010001110110111;
ROM[18804] <= 32'b01100001100000111000001110010011;
ROM[18805] <= 32'b00000000111000111000001110110011;
ROM[18806] <= 32'b00000000011100010010000000100011;
ROM[18807] <= 32'b00000000010000010000000100010011;
ROM[18808] <= 32'b00000000001100010010000000100011;
ROM[18809] <= 32'b00000000010000010000000100010011;
ROM[18810] <= 32'b00000000010000010010000000100011;
ROM[18811] <= 32'b00000000010000010000000100010011;
ROM[18812] <= 32'b00000000010100010010000000100011;
ROM[18813] <= 32'b00000000010000010000000100010011;
ROM[18814] <= 32'b00000000011000010010000000100011;
ROM[18815] <= 32'b00000000010000010000000100010011;
ROM[18816] <= 32'b00000001010000000000001110010011;
ROM[18817] <= 32'b00000000100000111000001110010011;
ROM[18818] <= 32'b01000000011100010000001110110011;
ROM[18819] <= 32'b00000000011100000000001000110011;
ROM[18820] <= 32'b00000000001000000000000110110011;
ROM[18821] <= 32'b01011001100000010111000011101111;
ROM[18822] <= 32'b00000110100100000000001110010011;
ROM[18823] <= 32'b00000000011100010010000000100011;
ROM[18824] <= 32'b00000000010000010000000100010011;
ROM[18825] <= 32'b00000000000000010010001110110111;
ROM[18826] <= 32'b01100111000000111000001110010011;
ROM[18827] <= 32'b00000000111000111000001110110011;
ROM[18828] <= 32'b00000000011100010010000000100011;
ROM[18829] <= 32'b00000000010000010000000100010011;
ROM[18830] <= 32'b00000000001100010010000000100011;
ROM[18831] <= 32'b00000000010000010000000100010011;
ROM[18832] <= 32'b00000000010000010010000000100011;
ROM[18833] <= 32'b00000000010000010000000100010011;
ROM[18834] <= 32'b00000000010100010010000000100011;
ROM[18835] <= 32'b00000000010000010000000100010011;
ROM[18836] <= 32'b00000000011000010010000000100011;
ROM[18837] <= 32'b00000000010000010000000100010011;
ROM[18838] <= 32'b00000001010000000000001110010011;
ROM[18839] <= 32'b00000000100000111000001110010011;
ROM[18840] <= 32'b01000000011100010000001110110011;
ROM[18841] <= 32'b00000000011100000000001000110011;
ROM[18842] <= 32'b00000000001000000000000110110011;
ROM[18843] <= 32'b01010100000000010111000011101111;
ROM[18844] <= 32'b00000111001100000000001110010011;
ROM[18845] <= 32'b00000000011100010010000000100011;
ROM[18846] <= 32'b00000000010000010000000100010011;
ROM[18847] <= 32'b00000000000000010010001110110111;
ROM[18848] <= 32'b01101100100000111000001110010011;
ROM[18849] <= 32'b00000000111000111000001110110011;
ROM[18850] <= 32'b00000000011100010010000000100011;
ROM[18851] <= 32'b00000000010000010000000100010011;
ROM[18852] <= 32'b00000000001100010010000000100011;
ROM[18853] <= 32'b00000000010000010000000100010011;
ROM[18854] <= 32'b00000000010000010010000000100011;
ROM[18855] <= 32'b00000000010000010000000100010011;
ROM[18856] <= 32'b00000000010100010010000000100011;
ROM[18857] <= 32'b00000000010000010000000100010011;
ROM[18858] <= 32'b00000000011000010010000000100011;
ROM[18859] <= 32'b00000000010000010000000100010011;
ROM[18860] <= 32'b00000001010000000000001110010011;
ROM[18861] <= 32'b00000000100000111000001110010011;
ROM[18862] <= 32'b01000000011100010000001110110011;
ROM[18863] <= 32'b00000000011100000000001000110011;
ROM[18864] <= 32'b00000000001000000000000110110011;
ROM[18865] <= 32'b01001110100000010111000011101111;
ROM[18866] <= 32'b00000010000000000000001110010011;
ROM[18867] <= 32'b00000000011100010010000000100011;
ROM[18868] <= 32'b00000000010000010000000100010011;
ROM[18869] <= 32'b00000000000000010010001110110111;
ROM[18870] <= 32'b01110010000000111000001110010011;
ROM[18871] <= 32'b00000000111000111000001110110011;
ROM[18872] <= 32'b00000000011100010010000000100011;
ROM[18873] <= 32'b00000000010000010000000100010011;
ROM[18874] <= 32'b00000000001100010010000000100011;
ROM[18875] <= 32'b00000000010000010000000100010011;
ROM[18876] <= 32'b00000000010000010010000000100011;
ROM[18877] <= 32'b00000000010000010000000100010011;
ROM[18878] <= 32'b00000000010100010010000000100011;
ROM[18879] <= 32'b00000000010000010000000100010011;
ROM[18880] <= 32'b00000000011000010010000000100011;
ROM[18881] <= 32'b00000000010000010000000100010011;
ROM[18882] <= 32'b00000001010000000000001110010011;
ROM[18883] <= 32'b00000000100000111000001110010011;
ROM[18884] <= 32'b01000000011100010000001110110011;
ROM[18885] <= 32'b00000000011100000000001000110011;
ROM[18886] <= 32'b00000000001000000000000110110011;
ROM[18887] <= 32'b01001001000000010111000011101111;
ROM[18888] <= 32'b00000110111000000000001110010011;
ROM[18889] <= 32'b00000000011100010010000000100011;
ROM[18890] <= 32'b00000000010000010000000100010011;
ROM[18891] <= 32'b00000000000000010010001110110111;
ROM[18892] <= 32'b01110111100000111000001110010011;
ROM[18893] <= 32'b00000000111000111000001110110011;
ROM[18894] <= 32'b00000000011100010010000000100011;
ROM[18895] <= 32'b00000000010000010000000100010011;
ROM[18896] <= 32'b00000000001100010010000000100011;
ROM[18897] <= 32'b00000000010000010000000100010011;
ROM[18898] <= 32'b00000000010000010010000000100011;
ROM[18899] <= 32'b00000000010000010000000100010011;
ROM[18900] <= 32'b00000000010100010010000000100011;
ROM[18901] <= 32'b00000000010000010000000100010011;
ROM[18902] <= 32'b00000000011000010010000000100011;
ROM[18903] <= 32'b00000000010000010000000100010011;
ROM[18904] <= 32'b00000001010000000000001110010011;
ROM[18905] <= 32'b00000000100000111000001110010011;
ROM[18906] <= 32'b01000000011100010000001110110011;
ROM[18907] <= 32'b00000000011100000000001000110011;
ROM[18908] <= 32'b00000000001000000000000110110011;
ROM[18909] <= 32'b01000011100000010111000011101111;
ROM[18910] <= 32'b00000110010100000000001110010011;
ROM[18911] <= 32'b00000000011100010010000000100011;
ROM[18912] <= 32'b00000000010000010000000100010011;
ROM[18913] <= 32'b00000000000000010010001110110111;
ROM[18914] <= 32'b01111101000000111000001110010011;
ROM[18915] <= 32'b00000000111000111000001110110011;
ROM[18916] <= 32'b00000000011100010010000000100011;
ROM[18917] <= 32'b00000000010000010000000100010011;
ROM[18918] <= 32'b00000000001100010010000000100011;
ROM[18919] <= 32'b00000000010000010000000100010011;
ROM[18920] <= 32'b00000000010000010010000000100011;
ROM[18921] <= 32'b00000000010000010000000100010011;
ROM[18922] <= 32'b00000000010100010010000000100011;
ROM[18923] <= 32'b00000000010000010000000100010011;
ROM[18924] <= 32'b00000000011000010010000000100011;
ROM[18925] <= 32'b00000000010000010000000100010011;
ROM[18926] <= 32'b00000001010000000000001110010011;
ROM[18927] <= 32'b00000000100000111000001110010011;
ROM[18928] <= 32'b01000000011100010000001110110011;
ROM[18929] <= 32'b00000000011100000000001000110011;
ROM[18930] <= 32'b00000000001000000000000110110011;
ROM[18931] <= 32'b00111110000000010111000011101111;
ROM[18932] <= 32'b00000110011100000000001110010011;
ROM[18933] <= 32'b00000000011100010010000000100011;
ROM[18934] <= 32'b00000000010000010000000100010011;
ROM[18935] <= 32'b00000000000000010011001110110111;
ROM[18936] <= 32'b10000010100000111000001110010011;
ROM[18937] <= 32'b00000000111000111000001110110011;
ROM[18938] <= 32'b00000000011100010010000000100011;
ROM[18939] <= 32'b00000000010000010000000100010011;
ROM[18940] <= 32'b00000000001100010010000000100011;
ROM[18941] <= 32'b00000000010000010000000100010011;
ROM[18942] <= 32'b00000000010000010010000000100011;
ROM[18943] <= 32'b00000000010000010000000100010011;
ROM[18944] <= 32'b00000000010100010010000000100011;
ROM[18945] <= 32'b00000000010000010000000100010011;
ROM[18946] <= 32'b00000000011000010010000000100011;
ROM[18947] <= 32'b00000000010000010000000100010011;
ROM[18948] <= 32'b00000001010000000000001110010011;
ROM[18949] <= 32'b00000000100000111000001110010011;
ROM[18950] <= 32'b01000000011100010000001110110011;
ROM[18951] <= 32'b00000000011100000000001000110011;
ROM[18952] <= 32'b00000000001000000000000110110011;
ROM[18953] <= 32'b00111000100000010111000011101111;
ROM[18954] <= 32'b00000110000100000000001110010011;
ROM[18955] <= 32'b00000000011100010010000000100011;
ROM[18956] <= 32'b00000000010000010000000100010011;
ROM[18957] <= 32'b00000000000000010011001110110111;
ROM[18958] <= 32'b10001000000000111000001110010011;
ROM[18959] <= 32'b00000000111000111000001110110011;
ROM[18960] <= 32'b00000000011100010010000000100011;
ROM[18961] <= 32'b00000000010000010000000100010011;
ROM[18962] <= 32'b00000000001100010010000000100011;
ROM[18963] <= 32'b00000000010000010000000100010011;
ROM[18964] <= 32'b00000000010000010010000000100011;
ROM[18965] <= 32'b00000000010000010000000100010011;
ROM[18966] <= 32'b00000000010100010010000000100011;
ROM[18967] <= 32'b00000000010000010000000100010011;
ROM[18968] <= 32'b00000000011000010010000000100011;
ROM[18969] <= 32'b00000000010000010000000100010011;
ROM[18970] <= 32'b00000001010000000000001110010011;
ROM[18971] <= 32'b00000000100000111000001110010011;
ROM[18972] <= 32'b01000000011100010000001110110011;
ROM[18973] <= 32'b00000000011100000000001000110011;
ROM[18974] <= 32'b00000000001000000000000110110011;
ROM[18975] <= 32'b00110011000000010111000011101111;
ROM[18976] <= 32'b00000111010000000000001110010011;
ROM[18977] <= 32'b00000000011100010010000000100011;
ROM[18978] <= 32'b00000000010000010000000100010011;
ROM[18979] <= 32'b00000000000000010011001110110111;
ROM[18980] <= 32'b10001101100000111000001110010011;
ROM[18981] <= 32'b00000000111000111000001110110011;
ROM[18982] <= 32'b00000000011100010010000000100011;
ROM[18983] <= 32'b00000000010000010000000100010011;
ROM[18984] <= 32'b00000000001100010010000000100011;
ROM[18985] <= 32'b00000000010000010000000100010011;
ROM[18986] <= 32'b00000000010000010010000000100011;
ROM[18987] <= 32'b00000000010000010000000100010011;
ROM[18988] <= 32'b00000000010100010010000000100011;
ROM[18989] <= 32'b00000000010000010000000100010011;
ROM[18990] <= 32'b00000000011000010010000000100011;
ROM[18991] <= 32'b00000000010000010000000100010011;
ROM[18992] <= 32'b00000001010000000000001110010011;
ROM[18993] <= 32'b00000000100000111000001110010011;
ROM[18994] <= 32'b01000000011100010000001110110011;
ROM[18995] <= 32'b00000000011100000000001000110011;
ROM[18996] <= 32'b00000000001000000000000110110011;
ROM[18997] <= 32'b00101101100000010111000011101111;
ROM[18998] <= 32'b00000110100100000000001110010011;
ROM[18999] <= 32'b00000000011100010010000000100011;
ROM[19000] <= 32'b00000000010000010000000100010011;
ROM[19001] <= 32'b00000000000000010011001110110111;
ROM[19002] <= 32'b10010011000000111000001110010011;
ROM[19003] <= 32'b00000000111000111000001110110011;
ROM[19004] <= 32'b00000000011100010010000000100011;
ROM[19005] <= 32'b00000000010000010000000100010011;
ROM[19006] <= 32'b00000000001100010010000000100011;
ROM[19007] <= 32'b00000000010000010000000100010011;
ROM[19008] <= 32'b00000000010000010010000000100011;
ROM[19009] <= 32'b00000000010000010000000100010011;
ROM[19010] <= 32'b00000000010100010010000000100011;
ROM[19011] <= 32'b00000000010000010000000100010011;
ROM[19012] <= 32'b00000000011000010010000000100011;
ROM[19013] <= 32'b00000000010000010000000100010011;
ROM[19014] <= 32'b00000001010000000000001110010011;
ROM[19015] <= 32'b00000000100000111000001110010011;
ROM[19016] <= 32'b01000000011100010000001110110011;
ROM[19017] <= 32'b00000000011100000000001000110011;
ROM[19018] <= 32'b00000000001000000000000110110011;
ROM[19019] <= 32'b00101000000000010111000011101111;
ROM[19020] <= 32'b00000111011000000000001110010011;
ROM[19021] <= 32'b00000000011100010010000000100011;
ROM[19022] <= 32'b00000000010000010000000100010011;
ROM[19023] <= 32'b00000000000000010011001110110111;
ROM[19024] <= 32'b10011000100000111000001110010011;
ROM[19025] <= 32'b00000000111000111000001110110011;
ROM[19026] <= 32'b00000000011100010010000000100011;
ROM[19027] <= 32'b00000000010000010000000100010011;
ROM[19028] <= 32'b00000000001100010010000000100011;
ROM[19029] <= 32'b00000000010000010000000100010011;
ROM[19030] <= 32'b00000000010000010010000000100011;
ROM[19031] <= 32'b00000000010000010000000100010011;
ROM[19032] <= 32'b00000000010100010010000000100011;
ROM[19033] <= 32'b00000000010000010000000100010011;
ROM[19034] <= 32'b00000000011000010010000000100011;
ROM[19035] <= 32'b00000000010000010000000100010011;
ROM[19036] <= 32'b00000001010000000000001110010011;
ROM[19037] <= 32'b00000000100000111000001110010011;
ROM[19038] <= 32'b01000000011100010000001110110011;
ROM[19039] <= 32'b00000000011100000000001000110011;
ROM[19040] <= 32'b00000000001000000000000110110011;
ROM[19041] <= 32'b00100010100000010111000011101111;
ROM[19042] <= 32'b00000110010100000000001110010011;
ROM[19043] <= 32'b00000000011100010010000000100011;
ROM[19044] <= 32'b00000000010000010000000100010011;
ROM[19045] <= 32'b00000000000000010011001110110111;
ROM[19046] <= 32'b10011110000000111000001110010011;
ROM[19047] <= 32'b00000000111000111000001110110011;
ROM[19048] <= 32'b00000000011100010010000000100011;
ROM[19049] <= 32'b00000000010000010000000100010011;
ROM[19050] <= 32'b00000000001100010010000000100011;
ROM[19051] <= 32'b00000000010000010000000100010011;
ROM[19052] <= 32'b00000000010000010010000000100011;
ROM[19053] <= 32'b00000000010000010000000100010011;
ROM[19054] <= 32'b00000000010100010010000000100011;
ROM[19055] <= 32'b00000000010000010000000100010011;
ROM[19056] <= 32'b00000000011000010010000000100011;
ROM[19057] <= 32'b00000000010000010000000100010011;
ROM[19058] <= 32'b00000001010000000000001110010011;
ROM[19059] <= 32'b00000000100000111000001110010011;
ROM[19060] <= 32'b01000000011100010000001110110011;
ROM[19061] <= 32'b00000000011100000000001000110011;
ROM[19062] <= 32'b00000000001000000000000110110011;
ROM[19063] <= 32'b00011101000000010111000011101111;
ROM[19064] <= 32'b00000101110000000000001110010011;
ROM[19065] <= 32'b00000000011100010010000000100011;
ROM[19066] <= 32'b00000000010000010000000100010011;
ROM[19067] <= 32'b00000000000000010011001110110111;
ROM[19068] <= 32'b10100011100000111000001110010011;
ROM[19069] <= 32'b00000000111000111000001110110011;
ROM[19070] <= 32'b00000000011100010010000000100011;
ROM[19071] <= 32'b00000000010000010000000100010011;
ROM[19072] <= 32'b00000000001100010010000000100011;
ROM[19073] <= 32'b00000000010000010000000100010011;
ROM[19074] <= 32'b00000000010000010010000000100011;
ROM[19075] <= 32'b00000000010000010000000100010011;
ROM[19076] <= 32'b00000000010100010010000000100011;
ROM[19077] <= 32'b00000000010000010000000100010011;
ROM[19078] <= 32'b00000000011000010010000000100011;
ROM[19079] <= 32'b00000000010000010000000100010011;
ROM[19080] <= 32'b00000001010000000000001110010011;
ROM[19081] <= 32'b00000000100000111000001110010011;
ROM[19082] <= 32'b01000000011100010000001110110011;
ROM[19083] <= 32'b00000000011100000000001000110011;
ROM[19084] <= 32'b00000000001000000000000110110011;
ROM[19085] <= 32'b00010111100000010111000011101111;
ROM[19086] <= 32'b00000110111000000000001110010011;
ROM[19087] <= 32'b00000000011100010010000000100011;
ROM[19088] <= 32'b00000000010000010000000100010011;
ROM[19089] <= 32'b00000000000000010011001110110111;
ROM[19090] <= 32'b10101001000000111000001110010011;
ROM[19091] <= 32'b00000000111000111000001110110011;
ROM[19092] <= 32'b00000000011100010010000000100011;
ROM[19093] <= 32'b00000000010000010000000100010011;
ROM[19094] <= 32'b00000000001100010010000000100011;
ROM[19095] <= 32'b00000000010000010000000100010011;
ROM[19096] <= 32'b00000000010000010010000000100011;
ROM[19097] <= 32'b00000000010000010000000100010011;
ROM[19098] <= 32'b00000000010100010010000000100011;
ROM[19099] <= 32'b00000000010000010000000100010011;
ROM[19100] <= 32'b00000000011000010010000000100011;
ROM[19101] <= 32'b00000000010000010000000100010011;
ROM[19102] <= 32'b00000001010000000000001110010011;
ROM[19103] <= 32'b00000000100000111000001110010011;
ROM[19104] <= 32'b01000000011100010000001110110011;
ROM[19105] <= 32'b00000000011100000000001000110011;
ROM[19106] <= 32'b00000000001000000000000110110011;
ROM[19107] <= 32'b00010010000000010111000011101111;
ROM[19108] <= 32'b00000000000000010011001110110111;
ROM[19109] <= 32'b10101101110000111000001110010011;
ROM[19110] <= 32'b00000000111000111000001110110011;
ROM[19111] <= 32'b00000000011100010010000000100011;
ROM[19112] <= 32'b00000000010000010000000100010011;
ROM[19113] <= 32'b00000000001100010010000000100011;
ROM[19114] <= 32'b00000000010000010000000100010011;
ROM[19115] <= 32'b00000000010000010010000000100011;
ROM[19116] <= 32'b00000000010000010000000100010011;
ROM[19117] <= 32'b00000000010100010010000000100011;
ROM[19118] <= 32'b00000000010000010000000100010011;
ROM[19119] <= 32'b00000000011000010010000000100011;
ROM[19120] <= 32'b00000000010000010000000100010011;
ROM[19121] <= 32'b00000001010000000000001110010011;
ROM[19122] <= 32'b00000000010000111000001110010011;
ROM[19123] <= 32'b01000000011100010000001110110011;
ROM[19124] <= 32'b00000000011100000000001000110011;
ROM[19125] <= 32'b00000000001000000000000110110011;
ROM[19126] <= 32'b00000000000000011001000011101111;
ROM[19127] <= 32'b11111111110000010000000100010011;
ROM[19128] <= 32'b00000000000000010010001110000011;
ROM[19129] <= 32'b00000000011101100010000000100011;
ROM[19130] <= 32'b00000000000000010011001110110111;
ROM[19131] <= 32'b10110011010000111000001110010011;
ROM[19132] <= 32'b00000000111000111000001110110011;
ROM[19133] <= 32'b00000000011100010010000000100011;
ROM[19134] <= 32'b00000000010000010000000100010011;
ROM[19135] <= 32'b00000000001100010010000000100011;
ROM[19136] <= 32'b00000000010000010000000100010011;
ROM[19137] <= 32'b00000000010000010010000000100011;
ROM[19138] <= 32'b00000000010000010000000100010011;
ROM[19139] <= 32'b00000000010100010010000000100011;
ROM[19140] <= 32'b00000000010000010000000100010011;
ROM[19141] <= 32'b00000000011000010010000000100011;
ROM[19142] <= 32'b00000000010000010000000100010011;
ROM[19143] <= 32'b00000001010000000000001110010011;
ROM[19144] <= 32'b00000000000000111000001110010011;
ROM[19145] <= 32'b01000000011100010000001110110011;
ROM[19146] <= 32'b00000000011100000000001000110011;
ROM[19147] <= 32'b00000000001000000000000110110011;
ROM[19148] <= 32'b01001111100000011000000011101111;
ROM[19149] <= 32'b11111111110000010000000100010011;
ROM[19150] <= 32'b00000000000000010010001110000011;
ROM[19151] <= 32'b00000000011101100010000000100011;
ROM[19152] <= 32'b00000000000100000000001110010011;
ROM[19153] <= 32'b00000000011100010010000000100011;
ROM[19154] <= 32'b00000000010000010000000100010011;
ROM[19155] <= 32'b11111111110000010000000100010011;
ROM[19156] <= 32'b00000000000000010010001110000011;
ROM[19157] <= 32'b01000000011100000000001110110011;
ROM[19158] <= 32'b00000000011100010010000000100011;
ROM[19159] <= 32'b00000000010000010000000100010011;
ROM[19160] <= 32'b00000001010000000000001110010011;
ROM[19161] <= 32'b01000000011100011000001110110011;
ROM[19162] <= 32'b00000000000000111010000010000011;
ROM[19163] <= 32'b11111111110000010000000100010011;
ROM[19164] <= 32'b00000000000000010010001110000011;
ROM[19165] <= 32'b00000000011100100010000000100011;
ROM[19166] <= 32'b00000000010000100000000100010011;
ROM[19167] <= 32'b00000001010000000000001110010011;
ROM[19168] <= 32'b01000000011100011000001110110011;
ROM[19169] <= 32'b00000000010000111010000110000011;
ROM[19170] <= 32'b00000000100000111010001000000011;
ROM[19171] <= 32'b00000000110000111010001010000011;
ROM[19172] <= 32'b00000001000000111010001100000011;
ROM[19173] <= 32'b00000000000000001000000011100111;
ROM[19174] <= 32'b00000000000000000000001110010011;
ROM[19175] <= 32'b00000000011100010010000000100011;
ROM[19176] <= 32'b00000000010000010000000100010011;
ROM[19177] <= 32'b11111111110000010000000100010011;
ROM[19178] <= 32'b00000000000000010010001110000011;
ROM[19179] <= 32'b00000000011100011010000000100011;
ROM[19180] <= 32'b00000111110000000000001110010011;
ROM[19181] <= 32'b00000000011100010010000000100011;
ROM[19182] <= 32'b00000000010000010000000100010011;
ROM[19183] <= 32'b11111111110000010000000100010011;
ROM[19184] <= 32'b00000000000000010010001110000011;
ROM[19185] <= 32'b00000000011100011010001000100011;
ROM[19186] <= 32'b00000000010000011010001110000011;
ROM[19187] <= 32'b00000000011100010010000000100011;
ROM[19188] <= 32'b00000000010000010000000100010011;
ROM[19189] <= 32'b00000000000000000000001110010011;
ROM[19190] <= 32'b00000000011100010010000000100011;
ROM[19191] <= 32'b00000000010000010000000100010011;
ROM[19192] <= 32'b11111111110000010000000100010011;
ROM[19193] <= 32'b00000000000000010010001110000011;
ROM[19194] <= 32'b11111111110000010000000100010011;
ROM[19195] <= 32'b00000000000000010010010000000011;
ROM[19196] <= 32'b00000000011101000010001110110011;
ROM[19197] <= 32'b00000000011100010010000000100011;
ROM[19198] <= 32'b00000000010000010000000100010011;
ROM[19199] <= 32'b11111111110000010000000100010011;
ROM[19200] <= 32'b00000000000000010010001110000011;
ROM[19201] <= 32'b01000000011100000000001110110011;
ROM[19202] <= 32'b00000000000100111000001110010011;
ROM[19203] <= 32'b00000000011100010010000000100011;
ROM[19204] <= 32'b00000000010000010000000100010011;
ROM[19205] <= 32'b11111111110000010000000100010011;
ROM[19206] <= 32'b00000000000000010010001110000011;
ROM[19207] <= 32'b01000000011100000000001110110011;
ROM[19208] <= 32'b00000000000100111000001110010011;
ROM[19209] <= 32'b00000000011100010010000000100011;
ROM[19210] <= 32'b00000000010000010000000100010011;
ROM[19211] <= 32'b11111111110000010000000100010011;
ROM[19212] <= 32'b00000000000000010010001110000011;
ROM[19213] <= 32'b00000000000000111000101001100011;
ROM[19214] <= 32'b00000000000000010011001110110111;
ROM[19215] <= 32'b11100101010000111000001110010011;
ROM[19216] <= 32'b00000000111000111000001110110011;
ROM[19217] <= 32'b00000000000000111000000011100111;
ROM[19218] <= 32'b00000000000000011010001110000011;
ROM[19219] <= 32'b00000000011100010010000000100011;
ROM[19220] <= 32'b00000000010000010000000100010011;
ROM[19221] <= 32'b00000100010001101010001110000011;
ROM[19222] <= 32'b00000000011100010010000000100011;
ROM[19223] <= 32'b00000000010000010000000100010011;
ROM[19224] <= 32'b00000000010000011010001110000011;
ROM[19225] <= 32'b00000000011100010010000000100011;
ROM[19226] <= 32'b00000000010000010000000100010011;
ROM[19227] <= 32'b11111111110000010000000100010011;
ROM[19228] <= 32'b00000000000000010010001110000011;
ROM[19229] <= 32'b11111111110000010000000100010011;
ROM[19230] <= 32'b00000000000000010010010000000011;
ROM[19231] <= 32'b00000000011101000000001110110011;
ROM[19232] <= 32'b00000000011100010010000000100011;
ROM[19233] <= 32'b00000000010000010000000100010011;
ROM[19234] <= 32'b11111111110000010000000100010011;
ROM[19235] <= 32'b00000000000000010010001110000011;
ROM[19236] <= 32'b00000000000000111000001100010011;
ROM[19237] <= 32'b00000000110100110000010000110011;
ROM[19238] <= 32'b00000000000001000010001110000011;
ROM[19239] <= 32'b00000000011100010010000000100011;
ROM[19240] <= 32'b00000000010000010000000100010011;
ROM[19241] <= 32'b11111111110000010000000100010011;
ROM[19242] <= 32'b00000000000000010010001110000011;
ROM[19243] <= 32'b11111111110000010000000100010011;
ROM[19244] <= 32'b00000000000000010010010000000011;
ROM[19245] <= 32'b00000000011101000000001110110011;
ROM[19246] <= 32'b00000000011100010010000000100011;
ROM[19247] <= 32'b00000000010000010000000100010011;
ROM[19248] <= 32'b11111111110000010000000100010011;
ROM[19249] <= 32'b00000000000000010010001110000011;
ROM[19250] <= 32'b00000000011100011010010000100011;
ROM[19251] <= 32'b00000000100000011010001110000011;
ROM[19252] <= 32'b00000000011100010010000000100011;
ROM[19253] <= 32'b00000000010000010000000100010011;
ROM[19254] <= 32'b00000000100000011010001110000011;
ROM[19255] <= 32'b00000000011100010010000000100011;
ROM[19256] <= 32'b00000000010000010000000100010011;
ROM[19257] <= 32'b00000000000000010011001110110111;
ROM[19258] <= 32'b11010011000000111000001110010011;
ROM[19259] <= 32'b00000000111000111000001110110011;
ROM[19260] <= 32'b00000000011100010010000000100011;
ROM[19261] <= 32'b00000000010000010000000100010011;
ROM[19262] <= 32'b00000000001100010010000000100011;
ROM[19263] <= 32'b00000000010000010000000100010011;
ROM[19264] <= 32'b00000000010000010010000000100011;
ROM[19265] <= 32'b00000000010000010000000100010011;
ROM[19266] <= 32'b00000000010100010010000000100011;
ROM[19267] <= 32'b00000000010000010000000100010011;
ROM[19268] <= 32'b00000000011000010010000000100011;
ROM[19269] <= 32'b00000000010000010000000100010011;
ROM[19270] <= 32'b00000001010000000000001110010011;
ROM[19271] <= 32'b00000000100000111000001110010011;
ROM[19272] <= 32'b01000000011100010000001110110011;
ROM[19273] <= 32'b00000000011100000000001000110011;
ROM[19274] <= 32'b00000000001000000000000110110011;
ROM[19275] <= 32'b10110000000111111110000011101111;
ROM[19276] <= 32'b11111111110000010000000100010011;
ROM[19277] <= 32'b00000000000000010010001110000011;
ROM[19278] <= 32'b00000000011100011010011000100011;
ROM[19279] <= 32'b00000000110000011010001110000011;
ROM[19280] <= 32'b00000000011100010010000000100011;
ROM[19281] <= 32'b00000000010000010000000100010011;
ROM[19282] <= 32'b00000000000000100010001110000011;
ROM[19283] <= 32'b00000000011100010010000000100011;
ROM[19284] <= 32'b00000000010000010000000100010011;
ROM[19285] <= 32'b11111111110000010000000100010011;
ROM[19286] <= 32'b00000000000000010010001110000011;
ROM[19287] <= 32'b11111111110000010000000100010011;
ROM[19288] <= 32'b00000000000000010010010000000011;
ROM[19289] <= 32'b00000000100000111010001110110011;
ROM[19290] <= 32'b00000000011100010010000000100011;
ROM[19291] <= 32'b00000000010000010000000100010011;
ROM[19292] <= 32'b11111111110000010000000100010011;
ROM[19293] <= 32'b00000000000000010010001110000011;
ROM[19294] <= 32'b01000000011100000000001110110011;
ROM[19295] <= 32'b00000000000100111000001110010011;
ROM[19296] <= 32'b00000000011100010010000000100011;
ROM[19297] <= 32'b00000000010000010000000100010011;
ROM[19298] <= 32'b00000000110000011010001110000011;
ROM[19299] <= 32'b00000000011100010010000000100011;
ROM[19300] <= 32'b00000000010000010000000100010011;
ROM[19301] <= 32'b00000000000000000000001110010011;
ROM[19302] <= 32'b00000000011100010010000000100011;
ROM[19303] <= 32'b00000000010000010000000100010011;
ROM[19304] <= 32'b11111111110000010000000100010011;
ROM[19305] <= 32'b00000000000000010010001110000011;
ROM[19306] <= 32'b11111111110000010000000100010011;
ROM[19307] <= 32'b00000000000000010010010000000011;
ROM[19308] <= 32'b00000000100000111010001110110011;
ROM[19309] <= 32'b00000000011100010010000000100011;
ROM[19310] <= 32'b00000000010000010000000100010011;
ROM[19311] <= 32'b11111111110000010000000100010011;
ROM[19312] <= 32'b00000000000000010010001110000011;
ROM[19313] <= 32'b11111111110000010000000100010011;
ROM[19314] <= 32'b00000000000000010010010000000011;
ROM[19315] <= 32'b00000000011101000111001110110011;
ROM[19316] <= 32'b00000000011100010010000000100011;
ROM[19317] <= 32'b00000000010000010000000100010011;
ROM[19318] <= 32'b11111111110000010000000100010011;
ROM[19319] <= 32'b00000000000000010010001110000011;
ROM[19320] <= 32'b00000000000000111000101001100011;
ROM[19321] <= 32'b00000000000000010011001110110111;
ROM[19322] <= 32'b11011111100000111000001110010011;
ROM[19323] <= 32'b00000000111000111000001110110011;
ROM[19324] <= 32'b00000000000000111000000011100111;
ROM[19325] <= 32'b00000001110000000000000011101111;
ROM[19326] <= 32'b00000000100000011010001110000011;
ROM[19327] <= 32'b00000000011100010010000000100011;
ROM[19328] <= 32'b00000000010000010000000100010011;
ROM[19329] <= 32'b11111111110000010000000100010011;
ROM[19330] <= 32'b00000000000000010010001110000011;
ROM[19331] <= 32'b00000000011100011010000000100011;
ROM[19332] <= 32'b00000000010000011010001110000011;
ROM[19333] <= 32'b00000000011100010010000000100011;
ROM[19334] <= 32'b00000000010000010000000100010011;
ROM[19335] <= 32'b00000000010000000000001110010011;
ROM[19336] <= 32'b00000000011100010010000000100011;
ROM[19337] <= 32'b00000000010000010000000100010011;
ROM[19338] <= 32'b11111111110000010000000100010011;
ROM[19339] <= 32'b00000000000000010010001110000011;
ROM[19340] <= 32'b11111111110000010000000100010011;
ROM[19341] <= 32'b00000000000000010010010000000011;
ROM[19342] <= 32'b01000000011101000000001110110011;
ROM[19343] <= 32'b00000000011100010010000000100011;
ROM[19344] <= 32'b00000000010000010000000100010011;
ROM[19345] <= 32'b11111111110000010000000100010011;
ROM[19346] <= 32'b00000000000000010010001110000011;
ROM[19347] <= 32'b00000000011100011010001000100011;
ROM[19348] <= 32'b11010111100111111111000011101111;
ROM[19349] <= 32'b00000000000000011010001110000011;
ROM[19350] <= 32'b00000000011100010010000000100011;
ROM[19351] <= 32'b00000000010000010000000100010011;
ROM[19352] <= 32'b00000001010000000000001110010011;
ROM[19353] <= 32'b01000000011100011000001110110011;
ROM[19354] <= 32'b00000000000000111010000010000011;
ROM[19355] <= 32'b11111111110000010000000100010011;
ROM[19356] <= 32'b00000000000000010010001110000011;
ROM[19357] <= 32'b00000000011100100010000000100011;
ROM[19358] <= 32'b00000000010000100000000100010011;
ROM[19359] <= 32'b00000001010000000000001110010011;
ROM[19360] <= 32'b01000000011100011000001110110011;
ROM[19361] <= 32'b00000000010000111010000110000011;
ROM[19362] <= 32'b00000000100000111010001000000011;
ROM[19363] <= 32'b00000000110000111010001010000011;
ROM[19364] <= 32'b00000001000000111010001100000011;
ROM[19365] <= 32'b00000000000000001000000011100111;
ROM[19366] <= 32'b00000000000000100010001110000011;
ROM[19367] <= 32'b00000000011100010010000000100011;
ROM[19368] <= 32'b00000000010000010000000100010011;
ROM[19369] <= 32'b00000000010000100010001110000011;
ROM[19370] <= 32'b00000000011100010010000000100011;
ROM[19371] <= 32'b00000000010000010000000100010011;
ROM[19372] <= 32'b11111111110000010000000100010011;
ROM[19373] <= 32'b00000000000000010010001110000011;
ROM[19374] <= 32'b11111111110000010000000100010011;
ROM[19375] <= 32'b00000000000000010010010000000011;
ROM[19376] <= 32'b00000000100000111010001110110011;
ROM[19377] <= 32'b00000000011100010010000000100011;
ROM[19378] <= 32'b00000000010000010000000100010011;
ROM[19379] <= 32'b11111111110000010000000100010011;
ROM[19380] <= 32'b00000000000000010010001110000011;
ROM[19381] <= 32'b00000000000000111000101001100011;
ROM[19382] <= 32'b00000000000000010011001110110111;
ROM[19383] <= 32'b11101110110000111000001110010011;
ROM[19384] <= 32'b00000000111000111000001110110011;
ROM[19385] <= 32'b00000000000000111000000011100111;
ROM[19386] <= 32'b00000100100000000000000011101111;
ROM[19387] <= 32'b00000000000000100010001110000011;
ROM[19388] <= 32'b00000000011100010010000000100011;
ROM[19389] <= 32'b00000000010000010000000100010011;
ROM[19390] <= 32'b00000001010000000000001110010011;
ROM[19391] <= 32'b01000000011100011000001110110011;
ROM[19392] <= 32'b00000000000000111010000010000011;
ROM[19393] <= 32'b11111111110000010000000100010011;
ROM[19394] <= 32'b00000000000000010010001110000011;
ROM[19395] <= 32'b00000000011100100010000000100011;
ROM[19396] <= 32'b00000000010000100000000100010011;
ROM[19397] <= 32'b00000001010000000000001110010011;
ROM[19398] <= 32'b01000000011100011000001110110011;
ROM[19399] <= 32'b00000000010000111010000110000011;
ROM[19400] <= 32'b00000000100000111010001000000011;
ROM[19401] <= 32'b00000000110000111010001010000011;
ROM[19402] <= 32'b00000001000000111010001100000011;
ROM[19403] <= 32'b00000000000000001000000011100111;
ROM[19404] <= 32'b00000000010000100010001110000011;
ROM[19405] <= 32'b00000000011100010010000000100011;
ROM[19406] <= 32'b00000000010000010000000100010011;
ROM[19407] <= 32'b00000001010000000000001110010011;
ROM[19408] <= 32'b01000000011100011000001110110011;
ROM[19409] <= 32'b00000000000000111010000010000011;
ROM[19410] <= 32'b11111111110000010000000100010011;
ROM[19411] <= 32'b00000000000000010010001110000011;
ROM[19412] <= 32'b00000000011100100010000000100011;
ROM[19413] <= 32'b00000000010000100000000100010011;
ROM[19414] <= 32'b00000001010000000000001110010011;
ROM[19415] <= 32'b01000000011100011000001110110011;
ROM[19416] <= 32'b00000000010000111010000110000011;
ROM[19417] <= 32'b00000000100000111010001000000011;
ROM[19418] <= 32'b00000000110000111010001010000011;
ROM[19419] <= 32'b00000001000000111010001100000011;
ROM[19420] <= 32'b00000000000000001000000011100111;
ROM[19421] <= 32'b00000000000000100010001110000011;
ROM[19422] <= 32'b00000000011100010010000000100011;
ROM[19423] <= 32'b00000000010000010000000100010011;
ROM[19424] <= 32'b00000000010000100010001110000011;
ROM[19425] <= 32'b00000000011100010010000000100011;
ROM[19426] <= 32'b00000000010000010000000100010011;
ROM[19427] <= 32'b11111111110000010000000100010011;
ROM[19428] <= 32'b00000000000000010010001110000011;
ROM[19429] <= 32'b11111111110000010000000100010011;
ROM[19430] <= 32'b00000000000000010010010000000011;
ROM[19431] <= 32'b00000000011101000010001110110011;
ROM[19432] <= 32'b00000000011100010010000000100011;
ROM[19433] <= 32'b00000000010000010000000100010011;
ROM[19434] <= 32'b11111111110000010000000100010011;
ROM[19435] <= 32'b00000000000000010010001110000011;
ROM[19436] <= 32'b00000000000000111000101001100011;
ROM[19437] <= 32'b00000000000000010011001110110111;
ROM[19438] <= 32'b11111100100000111000001110010011;
ROM[19439] <= 32'b00000000111000111000001110110011;
ROM[19440] <= 32'b00000000000000111000000011100111;
ROM[19441] <= 32'b00000100100000000000000011101111;
ROM[19442] <= 32'b00000000000000100010001110000011;
ROM[19443] <= 32'b00000000011100010010000000100011;
ROM[19444] <= 32'b00000000010000010000000100010011;
ROM[19445] <= 32'b00000001010000000000001110010011;
ROM[19446] <= 32'b01000000011100011000001110110011;
ROM[19447] <= 32'b00000000000000111010000010000011;
ROM[19448] <= 32'b11111111110000010000000100010011;
ROM[19449] <= 32'b00000000000000010010001110000011;
ROM[19450] <= 32'b00000000011100100010000000100011;
ROM[19451] <= 32'b00000000010000100000000100010011;
ROM[19452] <= 32'b00000001010000000000001110010011;
ROM[19453] <= 32'b01000000011100011000001110110011;
ROM[19454] <= 32'b00000000010000111010000110000011;
ROM[19455] <= 32'b00000000100000111010001000000011;
ROM[19456] <= 32'b00000000110000111010001010000011;
ROM[19457] <= 32'b00000001000000111010001100000011;
ROM[19458] <= 32'b00000000000000001000000011100111;
ROM[19459] <= 32'b00000000010000100010001110000011;
ROM[19460] <= 32'b00000000011100010010000000100011;
ROM[19461] <= 32'b00000000010000010000000100010011;
ROM[19462] <= 32'b00000001010000000000001110010011;
ROM[19463] <= 32'b01000000011100011000001110110011;
ROM[19464] <= 32'b00000000000000111010000010000011;
ROM[19465] <= 32'b11111111110000010000000100010011;
ROM[19466] <= 32'b00000000000000010010001110000011;
ROM[19467] <= 32'b00000000011100100010000000100011;
ROM[19468] <= 32'b00000000010000100000000100010011;
ROM[19469] <= 32'b00000001010000000000001110010011;
ROM[19470] <= 32'b01000000011100011000001110110011;
ROM[19471] <= 32'b00000000010000111010000110000011;
ROM[19472] <= 32'b00000000100000111010001000000011;
ROM[19473] <= 32'b00000000110000111010001010000011;
ROM[19474] <= 32'b00000001000000111010001100000011;
ROM[19475] <= 32'b00000000000000001000000011100111;
ROM[19476] <= 32'b00000000000000100010001110000011;
ROM[19477] <= 32'b00000000011100010010000000100011;
ROM[19478] <= 32'b00000000010000010000000100010011;
ROM[19479] <= 32'b00000000000000100010001110000011;
ROM[19480] <= 32'b00000000011100010010000000100011;
ROM[19481] <= 32'b00000000010000010000000100010011;
ROM[19482] <= 32'b00000000010000100010001110000011;
ROM[19483] <= 32'b00000000011100010010000000100011;
ROM[19484] <= 32'b00000000010000010000000100010011;
ROM[19485] <= 32'b00000000000000010011001110110111;
ROM[19486] <= 32'b00001100000000111000001110010011;
ROM[19487] <= 32'b00000000111000111000001110110011;
ROM[19488] <= 32'b00000000011100010010000000100011;
ROM[19489] <= 32'b00000000010000010000000100010011;
ROM[19490] <= 32'b00000000001100010010000000100011;
ROM[19491] <= 32'b00000000010000010000000100010011;
ROM[19492] <= 32'b00000000010000010010000000100011;
ROM[19493] <= 32'b00000000010000010000000100010011;
ROM[19494] <= 32'b00000000010100010010000000100011;
ROM[19495] <= 32'b00000000010000010000000100010011;
ROM[19496] <= 32'b00000000011000010010000000100011;
ROM[19497] <= 32'b00000000010000010000000100010011;
ROM[19498] <= 32'b00000001010000000000001110010011;
ROM[19499] <= 32'b00000000100000111000001110010011;
ROM[19500] <= 32'b01000000011100010000001110110011;
ROM[19501] <= 32'b00000000011100000000001000110011;
ROM[19502] <= 32'b00000000001000000000000110110011;
ROM[19503] <= 32'b10101110110111111110000011101111;
ROM[19504] <= 32'b00000000010000100010001110000011;
ROM[19505] <= 32'b00000000011100010010000000100011;
ROM[19506] <= 32'b00000000010000010000000100010011;
ROM[19507] <= 32'b00000000000000010011001110110111;
ROM[19508] <= 32'b00010001100000111000001110010011;
ROM[19509] <= 32'b00000000111000111000001110110011;
ROM[19510] <= 32'b00000000011100010010000000100011;
ROM[19511] <= 32'b00000000010000010000000100010011;
ROM[19512] <= 32'b00000000001100010010000000100011;
ROM[19513] <= 32'b00000000010000010000000100010011;
ROM[19514] <= 32'b00000000010000010010000000100011;
ROM[19515] <= 32'b00000000010000010000000100010011;
ROM[19516] <= 32'b00000000010100010010000000100011;
ROM[19517] <= 32'b00000000010000010000000100010011;
ROM[19518] <= 32'b00000000011000010010000000100011;
ROM[19519] <= 32'b00000000010000010000000100010011;
ROM[19520] <= 32'b00000001010000000000001110010011;
ROM[19521] <= 32'b00000000100000111000001110010011;
ROM[19522] <= 32'b01000000011100010000001110110011;
ROM[19523] <= 32'b00000000011100000000001000110011;
ROM[19524] <= 32'b00000000001000000000000110110011;
ROM[19525] <= 32'b11110001100011111110000011101111;
ROM[19526] <= 32'b11111111110000010000000100010011;
ROM[19527] <= 32'b00000000000000010010001110000011;
ROM[19528] <= 32'b11111111110000010000000100010011;
ROM[19529] <= 32'b00000000000000010010010000000011;
ROM[19530] <= 32'b01000000011101000000001110110011;
ROM[19531] <= 32'b00000000011100010010000000100011;
ROM[19532] <= 32'b00000000010000010000000100010011;
ROM[19533] <= 32'b00000001010000000000001110010011;
ROM[19534] <= 32'b01000000011100011000001110110011;
ROM[19535] <= 32'b00000000000000111010000010000011;
ROM[19536] <= 32'b11111111110000010000000100010011;
ROM[19537] <= 32'b00000000000000010010001110000011;
ROM[19538] <= 32'b00000000011100100010000000100011;
ROM[19539] <= 32'b00000000010000100000000100010011;
ROM[19540] <= 32'b00000001010000000000001110010011;
ROM[19541] <= 32'b01000000011100011000001110110011;
ROM[19542] <= 32'b00000000010000111010000110000011;
ROM[19543] <= 32'b00000000100000111010001000000011;
ROM[19544] <= 32'b00000000110000111010001010000011;
ROM[19545] <= 32'b00000001000000111010001100000011;
ROM[19546] <= 32'b00000000000000001000000011100111;
ROM[19547] <= 32'b00000000000000100010001110000011;
ROM[19548] <= 32'b00000000011100010010000000100011;
ROM[19549] <= 32'b00000000010000010000000100010011;
ROM[19550] <= 32'b00000000010000000000001110010011;
ROM[19551] <= 32'b00000000011100010010000000100011;
ROM[19552] <= 32'b00000000010000010000000100010011;
ROM[19553] <= 32'b00000000000000010011001110110111;
ROM[19554] <= 32'b00011101000000111000001110010011;
ROM[19555] <= 32'b00000000111000111000001110110011;
ROM[19556] <= 32'b00000000011100010010000000100011;
ROM[19557] <= 32'b00000000010000010000000100010011;
ROM[19558] <= 32'b00000000001100010010000000100011;
ROM[19559] <= 32'b00000000010000010000000100010011;
ROM[19560] <= 32'b00000000010000010010000000100011;
ROM[19561] <= 32'b00000000010000010000000100010011;
ROM[19562] <= 32'b00000000010100010010000000100011;
ROM[19563] <= 32'b00000000010000010000000100010011;
ROM[19564] <= 32'b00000000011000010010000000100011;
ROM[19565] <= 32'b00000000010000010000000100010011;
ROM[19566] <= 32'b00000001010000000000001110010011;
ROM[19567] <= 32'b00000000100000111000001110010011;
ROM[19568] <= 32'b01000000011100010000001110110011;
ROM[19569] <= 32'b00000000011100000000001000110011;
ROM[19570] <= 32'b00000000001000000000000110110011;
ROM[19571] <= 32'b11100110000011111110000011101111;
ROM[19572] <= 32'b11111111110000010000000100010011;
ROM[19573] <= 32'b00000000000000010010001110000011;
ROM[19574] <= 32'b00000000011100100010000000100011;
ROM[19575] <= 32'b00000100010001101010001110000011;
ROM[19576] <= 32'b00000000011100010010000000100011;
ROM[19577] <= 32'b00000000010000010000000100010011;
ROM[19578] <= 32'b00000000000000100010001110000011;
ROM[19579] <= 32'b00000000011100010010000000100011;
ROM[19580] <= 32'b00000000010000010000000100010011;
ROM[19581] <= 32'b11111111110000010000000100010011;
ROM[19582] <= 32'b00000000000000010010001110000011;
ROM[19583] <= 32'b11111111110000010000000100010011;
ROM[19584] <= 32'b00000000000000010010010000000011;
ROM[19585] <= 32'b00000000011101000000001110110011;
ROM[19586] <= 32'b00000000011100010010000000100011;
ROM[19587] <= 32'b00000000010000010000000100010011;
ROM[19588] <= 32'b11111111110000010000000100010011;
ROM[19589] <= 32'b00000000000000010010001110000011;
ROM[19590] <= 32'b00000000000000111000001100010011;
ROM[19591] <= 32'b00000000110100110000010000110011;
ROM[19592] <= 32'b00000000000001000010001110000011;
ROM[19593] <= 32'b00000000011100010010000000100011;
ROM[19594] <= 32'b00000000010000010000000100010011;
ROM[19595] <= 32'b00000001010000000000001110010011;
ROM[19596] <= 32'b01000000011100011000001110110011;
ROM[19597] <= 32'b00000000000000111010000010000011;
ROM[19598] <= 32'b11111111110000010000000100010011;
ROM[19599] <= 32'b00000000000000010010001110000011;
ROM[19600] <= 32'b00000000011100100010000000100011;
ROM[19601] <= 32'b00000000010000100000000100010011;
ROM[19602] <= 32'b00000001010000000000001110010011;
ROM[19603] <= 32'b01000000011100011000001110110011;
ROM[19604] <= 32'b00000000010000111010000110000011;
ROM[19605] <= 32'b00000000100000111010001000000011;
ROM[19606] <= 32'b00000000110000111010001010000011;
ROM[19607] <= 32'b00000001000000111010001100000011;
ROM[19608] <= 32'b00000000000000001000000011100111;
ROM[19609] <= 32'b00000000000000000010001110110111;
ROM[19610] <= 32'b00000000000000111000001110010011;
ROM[19611] <= 32'b00000000011100010010000000100011;
ROM[19612] <= 32'b00000000010000010000000100010011;
ROM[19613] <= 32'b11111111110000010000000100010011;
ROM[19614] <= 32'b00000000000000010010001110000011;
ROM[19615] <= 32'b00000100011101101010010000100011;
ROM[19616] <= 32'b00000000000000000100001110110111;
ROM[19617] <= 32'b00000000000000111000001110010011;
ROM[19618] <= 32'b00000000011100010010000000100011;
ROM[19619] <= 32'b00000000010000010000000100010011;
ROM[19620] <= 32'b11111111110000010000000100010011;
ROM[19621] <= 32'b00000000000000010010001110000011;
ROM[19622] <= 32'b00000100011101101010011000100011;
ROM[19623] <= 32'b00000100110001101010001110000011;
ROM[19624] <= 32'b00000000011100010010000000100011;
ROM[19625] <= 32'b00000000010000010000000100010011;
ROM[19626] <= 32'b00000100110001101010001110000011;
ROM[19627] <= 32'b00000000011100010010000000100011;
ROM[19628] <= 32'b00000000010000010000000100010011;
ROM[19629] <= 32'b11111111110000010000000100010011;
ROM[19630] <= 32'b00000000000000010010001110000011;
ROM[19631] <= 32'b11111111110000010000000100010011;
ROM[19632] <= 32'b00000000000000010010010000000011;
ROM[19633] <= 32'b00000000011101000000001110110011;
ROM[19634] <= 32'b00000000011100010010000000100011;
ROM[19635] <= 32'b00000000010000010000000100010011;
ROM[19636] <= 32'b00000100110001101010001110000011;
ROM[19637] <= 32'b00000000011100010010000000100011;
ROM[19638] <= 32'b00000000010000010000000100010011;
ROM[19639] <= 32'b11111111110000010000000100010011;
ROM[19640] <= 32'b00000000000000010010001110000011;
ROM[19641] <= 32'b11111111110000010000000100010011;
ROM[19642] <= 32'b00000000000000010010010000000011;
ROM[19643] <= 32'b00000000011101000000001110110011;
ROM[19644] <= 32'b00000000011100010010000000100011;
ROM[19645] <= 32'b00000000010000010000000100010011;
ROM[19646] <= 32'b00000100110001101010001110000011;
ROM[19647] <= 32'b00000000011100010010000000100011;
ROM[19648] <= 32'b00000000010000010000000100010011;
ROM[19649] <= 32'b11111111110000010000000100010011;
ROM[19650] <= 32'b00000000000000010010001110000011;
ROM[19651] <= 32'b11111111110000010000000100010011;
ROM[19652] <= 32'b00000000000000010010010000000011;
ROM[19653] <= 32'b00000000011101000000001110110011;
ROM[19654] <= 32'b00000000011100010010000000100011;
ROM[19655] <= 32'b00000000010000010000000100010011;
ROM[19656] <= 32'b11111111110000010000000100010011;
ROM[19657] <= 32'b00000000000000010010001110000011;
ROM[19658] <= 32'b00000100011101101010011000100011;
ROM[19659] <= 32'b00000000000000000001001110110111;
ROM[19660] <= 32'b10000000000000111000001110010011;
ROM[19661] <= 32'b00000000011100010010000000100011;
ROM[19662] <= 32'b00000000010000010000000100010011;
ROM[19663] <= 32'b11111111110000010000000100010011;
ROM[19664] <= 32'b00000000000000010010001110000011;
ROM[19665] <= 32'b00000100011101101010100000100011;
ROM[19666] <= 32'b00000000000000000100001110110111;
ROM[19667] <= 32'b00000000000000111000001110010011;
ROM[19668] <= 32'b00000000011100010010000000100011;
ROM[19669] <= 32'b00000000010000010000000100010011;
ROM[19670] <= 32'b11111111110000010000000100010011;
ROM[19671] <= 32'b00000000000000010010001110000011;
ROM[19672] <= 32'b00000100011101101010101000100011;
ROM[19673] <= 32'b00000000000000000000001110010011;
ROM[19674] <= 32'b00000000011100010010000000100011;
ROM[19675] <= 32'b00000000010000010000000100010011;
ROM[19676] <= 32'b11111111110000010000000100010011;
ROM[19677] <= 32'b00000000000000010010001110000011;
ROM[19678] <= 32'b00000100011101101010110000100011;
ROM[19679] <= 32'b00000100100001101010001110000011;
ROM[19680] <= 32'b00000000011100010010000000100011;
ROM[19681] <= 32'b00000000010000010000000100010011;
ROM[19682] <= 32'b11111111110000010000000100010011;
ROM[19683] <= 32'b00000000000000010010001110000011;
ROM[19684] <= 32'b00000100011101101010111000100011;
ROM[19685] <= 32'b00000000000000000000001110010011;
ROM[19686] <= 32'b00000000011100010010000000100011;
ROM[19687] <= 32'b00000000010000010000000100010011;
ROM[19688] <= 32'b11111111110000010000000100010011;
ROM[19689] <= 32'b00000000000000010010001110000011;
ROM[19690] <= 32'b00000110011101101010000000100011;
ROM[19691] <= 32'b00000000010000000000001110010011;
ROM[19692] <= 32'b00000000011100010010000000100011;
ROM[19693] <= 32'b00000000010000010000000100010011;
ROM[19694] <= 32'b11111111110000010000000100010011;
ROM[19695] <= 32'b00000000000000010010001110000011;
ROM[19696] <= 32'b00000110011101101010001000100011;
ROM[19697] <= 32'b00000101010001101010001110000011;
ROM[19698] <= 32'b00000000011100010010000000100011;
ROM[19699] <= 32'b00000000010000010000000100010011;
ROM[19700] <= 32'b00000101000001101010001110000011;
ROM[19701] <= 32'b00000000011100010010000000100011;
ROM[19702] <= 32'b00000000010000010000000100010011;
ROM[19703] <= 32'b11111111110000010000000100010011;
ROM[19704] <= 32'b00000000000000010010001110000011;
ROM[19705] <= 32'b11111111110000010000000100010011;
ROM[19706] <= 32'b00000000000000010010010000000011;
ROM[19707] <= 32'b01000000011101000000001110110011;
ROM[19708] <= 32'b00000000011100010010000000100011;
ROM[19709] <= 32'b00000000010000010000000100010011;
ROM[19710] <= 32'b00000101110001101010001110000011;
ROM[19711] <= 32'b00000000011100010010000000100011;
ROM[19712] <= 32'b00000000010000010000000100010011;
ROM[19713] <= 32'b00000110000001101010001110000011;
ROM[19714] <= 32'b00000000011100010010000000100011;
ROM[19715] <= 32'b00000000010000010000000100010011;
ROM[19716] <= 32'b11111111110000010000000100010011;
ROM[19717] <= 32'b00000000000000010010001110000011;
ROM[19718] <= 32'b11111111110000010000000100010011;
ROM[19719] <= 32'b00000000000000010010010000000011;
ROM[19720] <= 32'b00000000011101000000001110110011;
ROM[19721] <= 32'b00000000011100010010000000100011;
ROM[19722] <= 32'b00000000010000010000000100010011;
ROM[19723] <= 32'b11111111110000010000000100010011;
ROM[19724] <= 32'b00000000000000010010001110000011;
ROM[19725] <= 32'b00000000000000111000001100010011;
ROM[19726] <= 32'b11111111110000010000000100010011;
ROM[19727] <= 32'b00000000000000010010001110000011;
ROM[19728] <= 32'b00000000110100110000010000110011;
ROM[19729] <= 32'b00000000011101000010000000100011;
ROM[19730] <= 32'b00000000000000000000001110010011;
ROM[19731] <= 32'b00000000011100010010000000100011;
ROM[19732] <= 32'b00000000010000010000000100010011;
ROM[19733] <= 32'b00000101110001101010001110000011;
ROM[19734] <= 32'b00000000011100010010000000100011;
ROM[19735] <= 32'b00000000010000010000000100010011;
ROM[19736] <= 32'b00000110010001101010001110000011;
ROM[19737] <= 32'b00000000011100010010000000100011;
ROM[19738] <= 32'b00000000010000010000000100010011;
ROM[19739] <= 32'b11111111110000010000000100010011;
ROM[19740] <= 32'b00000000000000010010001110000011;
ROM[19741] <= 32'b11111111110000010000000100010011;
ROM[19742] <= 32'b00000000000000010010010000000011;
ROM[19743] <= 32'b00000000011101000000001110110011;
ROM[19744] <= 32'b00000000011100010010000000100011;
ROM[19745] <= 32'b00000000010000010000000100010011;
ROM[19746] <= 32'b11111111110000010000000100010011;
ROM[19747] <= 32'b00000000000000010010001110000011;
ROM[19748] <= 32'b00000000000000111000001100010011;
ROM[19749] <= 32'b11111111110000010000000100010011;
ROM[19750] <= 32'b00000000000000010010001110000011;
ROM[19751] <= 32'b00000000110100110000010000110011;
ROM[19752] <= 32'b00000000011101000010000000100011;
ROM[19753] <= 32'b00000000010000000000001110010011;
ROM[19754] <= 32'b00000000011100010010000000100011;
ROM[19755] <= 32'b00000000010000010000000100010011;
ROM[19756] <= 32'b11111111110000010000000100010011;
ROM[19757] <= 32'b00000000000000010010001110000011;
ROM[19758] <= 32'b01000000011100000000001110110011;
ROM[19759] <= 32'b00000000011100010010000000100011;
ROM[19760] <= 32'b00000000010000010000000100010011;
ROM[19761] <= 32'b11111111110000010000000100010011;
ROM[19762] <= 32'b00000000000000010010001110000011;
ROM[19763] <= 32'b00000110011101101010010000100011;
ROM[19764] <= 32'b00000000000000000000001110010011;
ROM[19765] <= 32'b00000000011100010010000000100011;
ROM[19766] <= 32'b00000000010000010000000100010011;
ROM[19767] <= 32'b00000001010000000000001110010011;
ROM[19768] <= 32'b01000000011100011000001110110011;
ROM[19769] <= 32'b00000000000000111010000010000011;
ROM[19770] <= 32'b11111111110000010000000100010011;
ROM[19771] <= 32'b00000000000000010010001110000011;
ROM[19772] <= 32'b00000000011100100010000000100011;
ROM[19773] <= 32'b00000000010000100000000100010011;
ROM[19774] <= 32'b00000001010000000000001110010011;
ROM[19775] <= 32'b01000000011100011000001110110011;
ROM[19776] <= 32'b00000000010000111010000110000011;
ROM[19777] <= 32'b00000000100000111010001000000011;
ROM[19778] <= 32'b00000000110000111010001010000011;
ROM[19779] <= 32'b00000001000000111010001100000011;
ROM[19780] <= 32'b00000000000000001000000011100111;
ROM[19781] <= 32'b00000000000000100010001110000011;
ROM[19782] <= 32'b00000000011100010010000000100011;
ROM[19783] <= 32'b00000000010000010000000100010011;
ROM[19784] <= 32'b00000000000000100010001110000011;
ROM[19785] <= 32'b00000000011100010010000000100011;
ROM[19786] <= 32'b00000000010000010000000100010011;
ROM[19787] <= 32'b11111111110000010000000100010011;
ROM[19788] <= 32'b00000000000000010010001110000011;
ROM[19789] <= 32'b11111111110000010000000100010011;
ROM[19790] <= 32'b00000000000000010010010000000011;
ROM[19791] <= 32'b00000000011101000000001110110011;
ROM[19792] <= 32'b00000000011100010010000000100011;
ROM[19793] <= 32'b00000000010000010000000100010011;
ROM[19794] <= 32'b11111111110000010000000100010011;
ROM[19795] <= 32'b00000000000000010010001110000011;
ROM[19796] <= 32'b00000000011100100010000000100011;
ROM[19797] <= 32'b00000000000000100010001110000011;
ROM[19798] <= 32'b00000000011100010010000000100011;
ROM[19799] <= 32'b00000000010000010000000100010011;
ROM[19800] <= 32'b00000000000000100010001110000011;
ROM[19801] <= 32'b00000000011100010010000000100011;
ROM[19802] <= 32'b00000000010000010000000100010011;
ROM[19803] <= 32'b11111111110000010000000100010011;
ROM[19804] <= 32'b00000000000000010010001110000011;
ROM[19805] <= 32'b11111111110000010000000100010011;
ROM[19806] <= 32'b00000000000000010010010000000011;
ROM[19807] <= 32'b00000000011101000000001110110011;
ROM[19808] <= 32'b00000000011100010010000000100011;
ROM[19809] <= 32'b00000000010000010000000100010011;
ROM[19810] <= 32'b11111111110000010000000100010011;
ROM[19811] <= 32'b00000000000000010010001110000011;
ROM[19812] <= 32'b00000000011100100010000000100011;
ROM[19813] <= 32'b00000101100001101010001110000011;
ROM[19814] <= 32'b00000000011100010010000000100011;
ROM[19815] <= 32'b00000000010000010000000100010011;
ROM[19816] <= 32'b00000000000000100010001110000011;
ROM[19817] <= 32'b00000000011100010010000000100011;
ROM[19818] <= 32'b00000000010000010000000100010011;
ROM[19819] <= 32'b11111111110000010000000100010011;
ROM[19820] <= 32'b00000000000000010010001110000011;
ROM[19821] <= 32'b11111111110000010000000100010011;
ROM[19822] <= 32'b00000000000000010010010000000011;
ROM[19823] <= 32'b00000000011101000000001110110011;
ROM[19824] <= 32'b00000000011100010010000000100011;
ROM[19825] <= 32'b00000000010000010000000100010011;
ROM[19826] <= 32'b11111111110000010000000100010011;
ROM[19827] <= 32'b00000000000000010010001110000011;
ROM[19828] <= 32'b00000000000000111000001100010011;
ROM[19829] <= 32'b00000000110100110000010000110011;
ROM[19830] <= 32'b00000000000001000010001110000011;
ROM[19831] <= 32'b00000000011100010010000000100011;
ROM[19832] <= 32'b00000000010000010000000100010011;
ROM[19833] <= 32'b00000001010000000000001110010011;
ROM[19834] <= 32'b01000000011100011000001110110011;
ROM[19835] <= 32'b00000000000000111010000010000011;
ROM[19836] <= 32'b11111111110000010000000100010011;
ROM[19837] <= 32'b00000000000000010010001110000011;
ROM[19838] <= 32'b00000000011100100010000000100011;
ROM[19839] <= 32'b00000000010000100000000100010011;
ROM[19840] <= 32'b00000001010000000000001110010011;
ROM[19841] <= 32'b01000000011100011000001110110011;
ROM[19842] <= 32'b00000000010000111010000110000011;
ROM[19843] <= 32'b00000000100000111010001000000011;
ROM[19844] <= 32'b00000000110000111010001010000011;
ROM[19845] <= 32'b00000001000000111010001100000011;
ROM[19846] <= 32'b00000000000000001000000011100111;
ROM[19847] <= 32'b00000000000000100010001110000011;
ROM[19848] <= 32'b00000000011100010010000000100011;
ROM[19849] <= 32'b00000000010000010000000100010011;
ROM[19850] <= 32'b00000000000000100010001110000011;
ROM[19851] <= 32'b00000000011100010010000000100011;
ROM[19852] <= 32'b00000000010000010000000100010011;
ROM[19853] <= 32'b11111111110000010000000100010011;
ROM[19854] <= 32'b00000000000000010010001110000011;
ROM[19855] <= 32'b11111111110000010000000100010011;
ROM[19856] <= 32'b00000000000000010010010000000011;
ROM[19857] <= 32'b00000000011101000000001110110011;
ROM[19858] <= 32'b00000000011100010010000000100011;
ROM[19859] <= 32'b00000000010000010000000100010011;
ROM[19860] <= 32'b11111111110000010000000100010011;
ROM[19861] <= 32'b00000000000000010010001110000011;
ROM[19862] <= 32'b00000000011100100010000000100011;
ROM[19863] <= 32'b00000000000000100010001110000011;
ROM[19864] <= 32'b00000000011100010010000000100011;
ROM[19865] <= 32'b00000000010000010000000100010011;
ROM[19866] <= 32'b00000000000000100010001110000011;
ROM[19867] <= 32'b00000000011100010010000000100011;
ROM[19868] <= 32'b00000000010000010000000100010011;
ROM[19869] <= 32'b11111111110000010000000100010011;
ROM[19870] <= 32'b00000000000000010010001110000011;
ROM[19871] <= 32'b11111111110000010000000100010011;
ROM[19872] <= 32'b00000000000000010010010000000011;
ROM[19873] <= 32'b00000000011101000000001110110011;
ROM[19874] <= 32'b00000000011100010010000000100011;
ROM[19875] <= 32'b00000000010000010000000100010011;
ROM[19876] <= 32'b11111111110000010000000100010011;
ROM[19877] <= 32'b00000000000000010010001110000011;
ROM[19878] <= 32'b00000000011100100010000000100011;
ROM[19879] <= 32'b00000000010000100010001110000011;
ROM[19880] <= 32'b00000000011100010010000000100011;
ROM[19881] <= 32'b00000000010000010000000100010011;
ROM[19882] <= 32'b00000101100001101010001110000011;
ROM[19883] <= 32'b00000000011100010010000000100011;
ROM[19884] <= 32'b00000000010000010000000100010011;
ROM[19885] <= 32'b00000000000000100010001110000011;
ROM[19886] <= 32'b00000000011100010010000000100011;
ROM[19887] <= 32'b00000000010000010000000100010011;
ROM[19888] <= 32'b11111111110000010000000100010011;
ROM[19889] <= 32'b00000000000000010010001110000011;
ROM[19890] <= 32'b11111111110000010000000100010011;
ROM[19891] <= 32'b00000000000000010010010000000011;
ROM[19892] <= 32'b00000000011101000000001110110011;
ROM[19893] <= 32'b00000000011100010010000000100011;
ROM[19894] <= 32'b00000000010000010000000100010011;
ROM[19895] <= 32'b11111111110000010000000100010011;
ROM[19896] <= 32'b00000000000000010010001110000011;
ROM[19897] <= 32'b00000000000000111000001100010011;
ROM[19898] <= 32'b11111111110000010000000100010011;
ROM[19899] <= 32'b00000000000000010010001110000011;
ROM[19900] <= 32'b00000000110100110000010000110011;
ROM[19901] <= 32'b00000000011101000010000000100011;
ROM[19902] <= 32'b00000000000000000000001110010011;
ROM[19903] <= 32'b00000000011100010010000000100011;
ROM[19904] <= 32'b00000000010000010000000100010011;
ROM[19905] <= 32'b00000001010000000000001110010011;
ROM[19906] <= 32'b01000000011100011000001110110011;
ROM[19907] <= 32'b00000000000000111010000010000011;
ROM[19908] <= 32'b11111111110000010000000100010011;
ROM[19909] <= 32'b00000000000000010010001110000011;
ROM[19910] <= 32'b00000000011100100010000000100011;
ROM[19911] <= 32'b00000000010000100000000100010011;
ROM[19912] <= 32'b00000001010000000000001110010011;
ROM[19913] <= 32'b01000000011100011000001110110011;
ROM[19914] <= 32'b00000000010000111010000110000011;
ROM[19915] <= 32'b00000000100000111010001000000011;
ROM[19916] <= 32'b00000000110000111010001010000011;
ROM[19917] <= 32'b00000001000000111010001100000011;
ROM[19918] <= 32'b00000000000000001000000011100111;
ROM[19919] <= 32'b00000000000000010010000000100011;
ROM[19920] <= 32'b00000000010000010000000100010011;
ROM[19921] <= 32'b00000000000000010010000000100011;
ROM[19922] <= 32'b00000000010000010000000100010011;
ROM[19923] <= 32'b00000000000000010010000000100011;
ROM[19924] <= 32'b00000000010000010000000100010011;
ROM[19925] <= 32'b00000000000000010010000000100011;
ROM[19926] <= 32'b00000000010000010000000100010011;
ROM[19927] <= 32'b00000000000000000000001110010011;
ROM[19928] <= 32'b00000000011100010010000000100011;
ROM[19929] <= 32'b00000000010000010000000100010011;
ROM[19930] <= 32'b11111111110000010000000100010011;
ROM[19931] <= 32'b00000000000000010010001110000011;
ROM[19932] <= 32'b00000000011100011010001000100011;
ROM[19933] <= 32'b00000101010001101010001110000011;
ROM[19934] <= 32'b00000000011100010010000000100011;
ROM[19935] <= 32'b00000000010000010000000100010011;
ROM[19936] <= 32'b00000101000001101010001110000011;
ROM[19937] <= 32'b00000000011100010010000000100011;
ROM[19938] <= 32'b00000000010000010000000100010011;
ROM[19939] <= 32'b11111111110000010000000100010011;
ROM[19940] <= 32'b00000000000000010010001110000011;
ROM[19941] <= 32'b11111111110000010000000100010011;
ROM[19942] <= 32'b00000000000000010010010000000011;
ROM[19943] <= 32'b01000000011101000000001110110011;
ROM[19944] <= 32'b00000000011100010010000000100011;
ROM[19945] <= 32'b00000000010000010000000100010011;
ROM[19946] <= 32'b11111111110000010000000100010011;
ROM[19947] <= 32'b00000000000000010010001110000011;
ROM[19948] <= 32'b00000000011100011010010000100011;
ROM[19949] <= 32'b00000101110001101010001110000011;
ROM[19950] <= 32'b00000000011100010010000000100011;
ROM[19951] <= 32'b00000000010000010000000100010011;
ROM[19952] <= 32'b11111111110000010000000100010011;
ROM[19953] <= 32'b00000000000000010010001110000011;
ROM[19954] <= 32'b00000000011100011010000000100011;
ROM[19955] <= 32'b00000000000000011010001110000011;
ROM[19956] <= 32'b00000000011100010010000000100011;
ROM[19957] <= 32'b00000000010000010000000100010011;
ROM[19958] <= 32'b00000110010001101010001110000011;
ROM[19959] <= 32'b00000000011100010010000000100011;
ROM[19960] <= 32'b00000000010000010000000100010011;
ROM[19961] <= 32'b11111111110000010000000100010011;
ROM[19962] <= 32'b00000000000000010010001110000011;
ROM[19963] <= 32'b11111111110000010000000100010011;
ROM[19964] <= 32'b00000000000000010010010000000011;
ROM[19965] <= 32'b00000000011101000000001110110011;
ROM[19966] <= 32'b00000000011100010010000000100011;
ROM[19967] <= 32'b00000000010000010000000100010011;
ROM[19968] <= 32'b11111111110000010000000100010011;
ROM[19969] <= 32'b00000000000000010010001110000011;
ROM[19970] <= 32'b00000000000000111000001100010011;
ROM[19971] <= 32'b00000000110100110000010000110011;
ROM[19972] <= 32'b00000000000001000010001110000011;
ROM[19973] <= 32'b00000000011100010010000000100011;
ROM[19974] <= 32'b00000000010000010000000100010011;
ROM[19975] <= 32'b00000000000000000000001110010011;
ROM[19976] <= 32'b00000000011100010010000000100011;
ROM[19977] <= 32'b00000000010000010000000100010011;
ROM[19978] <= 32'b11111111110000010000000100010011;
ROM[19979] <= 32'b00000000000000010010001110000011;
ROM[19980] <= 32'b11111111110000010000000100010011;
ROM[19981] <= 32'b00000000000000010010010000000011;
ROM[19982] <= 32'b00000000011101000010010010110011;
ROM[19983] <= 32'b00000000100000111010010100110011;
ROM[19984] <= 32'b00000000101001001000001110110011;
ROM[19985] <= 32'b00000000000100111000001110010011;
ROM[19986] <= 32'b00000000000100111111001110010011;
ROM[19987] <= 32'b00000000011100010010000000100011;
ROM[19988] <= 32'b00000000010000010000000100010011;
ROM[19989] <= 32'b11111111110000010000000100010011;
ROM[19990] <= 32'b00000000000000010010001110000011;
ROM[19991] <= 32'b00000000000000111000101001100011;
ROM[19992] <= 32'b00000000000000010100001110110111;
ROM[19993] <= 32'b10000111010000111000001110010011;
ROM[19994] <= 32'b00000000111000111000001110110011;
ROM[19995] <= 32'b00000000000000111000000011100111;
ROM[19996] <= 32'b00000100100000000000000011101111;
ROM[19997] <= 32'b00000000000000011010001110000011;
ROM[19998] <= 32'b00000000011100010010000000100011;
ROM[19999] <= 32'b00000000010000010000000100010011;
ROM[20000] <= 32'b00000001010000000000001110010011;
ROM[20001] <= 32'b01000000011100011000001110110011;
ROM[20002] <= 32'b00000000000000111010000010000011;
ROM[20003] <= 32'b11111111110000010000000100010011;
ROM[20004] <= 32'b00000000000000010010001110000011;
ROM[20005] <= 32'b00000000011100100010000000100011;
ROM[20006] <= 32'b00000000010000100000000100010011;
ROM[20007] <= 32'b00000001010000000000001110010011;
ROM[20008] <= 32'b01000000011100011000001110110011;
ROM[20009] <= 32'b00000000010000111010000110000011;
ROM[20010] <= 32'b00000000100000111010001000000011;
ROM[20011] <= 32'b00000000110000111010001010000011;
ROM[20012] <= 32'b00000001000000111010001100000011;
ROM[20013] <= 32'b00000000000000001000000011100111;
ROM[20014] <= 32'b00000000000000011010001110000011;
ROM[20015] <= 32'b00000000011100010010000000100011;
ROM[20016] <= 32'b00000000010000010000000100010011;
ROM[20017] <= 32'b00000000000000000000001110010011;
ROM[20018] <= 32'b00000000011100010010000000100011;
ROM[20019] <= 32'b00000000010000010000000100010011;
ROM[20020] <= 32'b11111111110000010000000100010011;
ROM[20021] <= 32'b00000000000000010010001110000011;
ROM[20022] <= 32'b11111111110000010000000100010011;
ROM[20023] <= 32'b00000000000000010010010000000011;
ROM[20024] <= 32'b00000000011101000010010010110011;
ROM[20025] <= 32'b00000000100000111010010100110011;
ROM[20026] <= 32'b00000000101001001000001110110011;
ROM[20027] <= 32'b00000000000100111000001110010011;
ROM[20028] <= 32'b00000000000100111111001110010011;
ROM[20029] <= 32'b00000000011100010010000000100011;
ROM[20030] <= 32'b00000000010000010000000100010011;
ROM[20031] <= 32'b11111111110000010000000100010011;
ROM[20032] <= 32'b00000000000000010010001110000011;
ROM[20033] <= 32'b01000000011100000000001110110011;
ROM[20034] <= 32'b00000000000100111000001110010011;
ROM[20035] <= 32'b00000000011100010010000000100011;
ROM[20036] <= 32'b00000000010000010000000100010011;
ROM[20037] <= 32'b11111111110000010000000100010011;
ROM[20038] <= 32'b00000000000000010010001110000011;
ROM[20039] <= 32'b01000000011100000000001110110011;
ROM[20040] <= 32'b00000000000100111000001110010011;
ROM[20041] <= 32'b00000000011100010010000000100011;
ROM[20042] <= 32'b00000000010000010000000100010011;
ROM[20043] <= 32'b11111111110000010000000100010011;
ROM[20044] <= 32'b00000000000000010010001110000011;
ROM[20045] <= 32'b00000000000000111000101001100011;
ROM[20046] <= 32'b00000000000000010100001110110111;
ROM[20047] <= 32'b10110001100000111000001110010011;
ROM[20048] <= 32'b00000000111000111000001110110011;
ROM[20049] <= 32'b00000000000000111000000011100111;
ROM[20050] <= 32'b00000000000000011010001110000011;
ROM[20051] <= 32'b00000000011100010010000000100011;
ROM[20052] <= 32'b00000000010000010000000100010011;
ROM[20053] <= 32'b00000110000001101010001110000011;
ROM[20054] <= 32'b00000000011100010010000000100011;
ROM[20055] <= 32'b00000000010000010000000100010011;
ROM[20056] <= 32'b11111111110000010000000100010011;
ROM[20057] <= 32'b00000000000000010010001110000011;
ROM[20058] <= 32'b11111111110000010000000100010011;
ROM[20059] <= 32'b00000000000000010010010000000011;
ROM[20060] <= 32'b00000000011101000000001110110011;
ROM[20061] <= 32'b00000000011100010010000000100011;
ROM[20062] <= 32'b00000000010000010000000100010011;
ROM[20063] <= 32'b11111111110000010000000100010011;
ROM[20064] <= 32'b00000000000000010010001110000011;
ROM[20065] <= 32'b00000000000000111000001100010011;
ROM[20066] <= 32'b00000000110100110000010000110011;
ROM[20067] <= 32'b00000000000001000010001110000011;
ROM[20068] <= 32'b00000000011100010010000000100011;
ROM[20069] <= 32'b00000000010000010000000100010011;
ROM[20070] <= 32'b00000000000100000000001110010011;
ROM[20071] <= 32'b00000000011100010010000000100011;
ROM[20072] <= 32'b00000000010000010000000100010011;
ROM[20073] <= 32'b11111111110000010000000100010011;
ROM[20074] <= 32'b00000000000000010010001110000011;
ROM[20075] <= 32'b11111111110000010000000100010011;
ROM[20076] <= 32'b00000000000000010010010000000011;
ROM[20077] <= 32'b01000000011101000000001110110011;
ROM[20078] <= 32'b00000000011100010010000000100011;
ROM[20079] <= 32'b00000000010000010000000100010011;
ROM[20080] <= 32'b11111111110000010000000100010011;
ROM[20081] <= 32'b00000000000000010010001110000011;
ROM[20082] <= 32'b00000000011100011010011000100011;
ROM[20083] <= 32'b00000000110000011010001110000011;
ROM[20084] <= 32'b00000000011100010010000000100011;
ROM[20085] <= 32'b00000000010000010000000100010011;
ROM[20086] <= 32'b00000000000000100010001110000011;
ROM[20087] <= 32'b00000000011100010010000000100011;
ROM[20088] <= 32'b00000000010000010000000100010011;
ROM[20089] <= 32'b11111111110000010000000100010011;
ROM[20090] <= 32'b00000000000000010010001110000011;
ROM[20091] <= 32'b11111111110000010000000100010011;
ROM[20092] <= 32'b00000000000000010010010000000011;
ROM[20093] <= 32'b00000000011101000010001110110011;
ROM[20094] <= 32'b00000000011100010010000000100011;
ROM[20095] <= 32'b00000000010000010000000100010011;
ROM[20096] <= 32'b11111111110000010000000100010011;
ROM[20097] <= 32'b00000000000000010010001110000011;
ROM[20098] <= 32'b01000000011100000000001110110011;
ROM[20099] <= 32'b00000000000100111000001110010011;
ROM[20100] <= 32'b00000000011100010010000000100011;
ROM[20101] <= 32'b00000000010000010000000100010011;
ROM[20102] <= 32'b00000000110000011010001110000011;
ROM[20103] <= 32'b00000000011100010010000000100011;
ROM[20104] <= 32'b00000000010000010000000100010011;
ROM[20105] <= 32'b00000000100000011010001110000011;
ROM[20106] <= 32'b00000000011100010010000000100011;
ROM[20107] <= 32'b00000000010000010000000100010011;
ROM[20108] <= 32'b11111111110000010000000100010011;
ROM[20109] <= 32'b00000000000000010010001110000011;
ROM[20110] <= 32'b11111111110000010000000100010011;
ROM[20111] <= 32'b00000000000000010010010000000011;
ROM[20112] <= 32'b00000000011101000010001110110011;
ROM[20113] <= 32'b00000000011100010010000000100011;
ROM[20114] <= 32'b00000000010000010000000100010011;
ROM[20115] <= 32'b11111111110000010000000100010011;
ROM[20116] <= 32'b00000000000000010010001110000011;
ROM[20117] <= 32'b11111111110000010000000100010011;
ROM[20118] <= 32'b00000000000000010010010000000011;
ROM[20119] <= 32'b00000000011101000111001110110011;
ROM[20120] <= 32'b00000000011100010010000000100011;
ROM[20121] <= 32'b00000000010000010000000100010011;
ROM[20122] <= 32'b11111111110000010000000100010011;
ROM[20123] <= 32'b00000000000000010010001110000011;
ROM[20124] <= 32'b00000000000000111000101001100011;
ROM[20125] <= 32'b00000000000000010100001110110111;
ROM[20126] <= 32'b10101000100000111000001110010011;
ROM[20127] <= 32'b00000000111000111000001110110011;
ROM[20128] <= 32'b00000000000000111000000011100111;
ROM[20129] <= 32'b00000011010000000000000011101111;
ROM[20130] <= 32'b00000000000000011010001110000011;
ROM[20131] <= 32'b00000000011100010010000000100011;
ROM[20132] <= 32'b00000000010000010000000100010011;
ROM[20133] <= 32'b11111111110000010000000100010011;
ROM[20134] <= 32'b00000000000000010010001110000011;
ROM[20135] <= 32'b00000000011100011010001000100011;
ROM[20136] <= 32'b00000000110000011010001110000011;
ROM[20137] <= 32'b00000000011100010010000000100011;
ROM[20138] <= 32'b00000000010000010000000100010011;
ROM[20139] <= 32'b11111111110000010000000100010011;
ROM[20140] <= 32'b00000000000000010010001110000011;
ROM[20141] <= 32'b00000000011100011010010000100011;
ROM[20142] <= 32'b00000000000000011010001110000011;
ROM[20143] <= 32'b00000000011100010010000000100011;
ROM[20144] <= 32'b00000000010000010000000100010011;
ROM[20145] <= 32'b00000110010001101010001110000011;
ROM[20146] <= 32'b00000000011100010010000000100011;
ROM[20147] <= 32'b00000000010000010000000100010011;
ROM[20148] <= 32'b11111111110000010000000100010011;
ROM[20149] <= 32'b00000000000000010010001110000011;
ROM[20150] <= 32'b11111111110000010000000100010011;
ROM[20151] <= 32'b00000000000000010010010000000011;
ROM[20152] <= 32'b00000000011101000000001110110011;
ROM[20153] <= 32'b00000000011100010010000000100011;
ROM[20154] <= 32'b00000000010000010000000100010011;
ROM[20155] <= 32'b11111111110000010000000100010011;
ROM[20156] <= 32'b00000000000000010010001110000011;
ROM[20157] <= 32'b00000000000000111000001100010011;
ROM[20158] <= 32'b00000000110100110000010000110011;
ROM[20159] <= 32'b00000000000001000010001110000011;
ROM[20160] <= 32'b00000000011100010010000000100011;
ROM[20161] <= 32'b00000000010000010000000100010011;
ROM[20162] <= 32'b11111111110000010000000100010011;
ROM[20163] <= 32'b00000000000000010010001110000011;
ROM[20164] <= 32'b00000000011100011010000000100011;
ROM[20165] <= 32'b11011010010111111111000011101111;
ROM[20166] <= 32'b00000000010000011010001110000011;
ROM[20167] <= 32'b00000000011100010010000000100011;
ROM[20168] <= 32'b00000000010000010000000100010011;
ROM[20169] <= 32'b00000001010000000000001110010011;
ROM[20170] <= 32'b01000000011100011000001110110011;
ROM[20171] <= 32'b00000000000000111010000010000011;
ROM[20172] <= 32'b11111111110000010000000100010011;
ROM[20173] <= 32'b00000000000000010010001110000011;
ROM[20174] <= 32'b00000000011100100010000000100011;
ROM[20175] <= 32'b00000000010000100000000100010011;
ROM[20176] <= 32'b00000001010000000000001110010011;
ROM[20177] <= 32'b01000000011100011000001110110011;
ROM[20178] <= 32'b00000000010000111010000110000011;
ROM[20179] <= 32'b00000000100000111010001000000011;
ROM[20180] <= 32'b00000000110000111010001010000011;
ROM[20181] <= 32'b00000001000000111010001100000011;
ROM[20182] <= 32'b00000000000000001000000011100111;
ROM[20183] <= 32'b00000000000000010010000000100011;
ROM[20184] <= 32'b00000000010000010000000100010011;
ROM[20185] <= 32'b00000000000000010010000000100011;
ROM[20186] <= 32'b00000000010000010000000100010011;
ROM[20187] <= 32'b00000000000000010010000000100011;
ROM[20188] <= 32'b00000000010000010000000100010011;
ROM[20189] <= 32'b00000000000000100010001110000011;
ROM[20190] <= 32'b00000000011100010010000000100011;
ROM[20191] <= 32'b00000000010000010000000100010011;
ROM[20192] <= 32'b00000110100001101010001110000011;
ROM[20193] <= 32'b00000000011100010010000000100011;
ROM[20194] <= 32'b00000000010000010000000100010011;
ROM[20195] <= 32'b11111111110000010000000100010011;
ROM[20196] <= 32'b00000000000000010010001110000011;
ROM[20197] <= 32'b11111111110000010000000100010011;
ROM[20198] <= 32'b00000000000000010010010000000011;
ROM[20199] <= 32'b00000000011101000000001110110011;
ROM[20200] <= 32'b00000000011100010010000000100011;
ROM[20201] <= 32'b00000000010000010000000100010011;
ROM[20202] <= 32'b11111111110000010000000100010011;
ROM[20203] <= 32'b00000000000000010010001110000011;
ROM[20204] <= 32'b00000000000000111000001100010011;
ROM[20205] <= 32'b00000000110100110000010000110011;
ROM[20206] <= 32'b00000000000001000010001110000011;
ROM[20207] <= 32'b00000000011100010010000000100011;
ROM[20208] <= 32'b00000000010000010000000100010011;
ROM[20209] <= 32'b11111111110000010000000100010011;
ROM[20210] <= 32'b00000000000000010010001110000011;
ROM[20211] <= 32'b00000000011100011010010000100011;
ROM[20212] <= 32'b00000000000000100010001110000011;
ROM[20213] <= 32'b00000000011100010010000000100011;
ROM[20214] <= 32'b00000000010000010000000100010011;
ROM[20215] <= 32'b00000000000100000000001110010011;
ROM[20216] <= 32'b00000000011100010010000000100011;
ROM[20217] <= 32'b00000000010000010000000100010011;
ROM[20218] <= 32'b11111111110000010000000100010011;
ROM[20219] <= 32'b00000000000000010010001110000011;
ROM[20220] <= 32'b11111111110000010000000100010011;
ROM[20221] <= 32'b00000000000000010010010000000011;
ROM[20222] <= 32'b00000000011101000000001110110011;
ROM[20223] <= 32'b00000000011100010010000000100011;
ROM[20224] <= 32'b00000000010000010000000100010011;
ROM[20225] <= 32'b11111111110000010000000100010011;
ROM[20226] <= 32'b00000000000000010010001110000011;
ROM[20227] <= 32'b00000000011100100010000000100011;
ROM[20228] <= 32'b00000000000000100010001110000011;
ROM[20229] <= 32'b00000000011100010010000000100011;
ROM[20230] <= 32'b00000000010000010000000100010011;
ROM[20231] <= 32'b00000000000000010100001110110111;
ROM[20232] <= 32'b11000110100000111000001110010011;
ROM[20233] <= 32'b00000000111000111000001110110011;
ROM[20234] <= 32'b00000000011100010010000000100011;
ROM[20235] <= 32'b00000000010000010000000100010011;
ROM[20236] <= 32'b00000000001100010010000000100011;
ROM[20237] <= 32'b00000000010000010000000100010011;
ROM[20238] <= 32'b00000000010000010010000000100011;
ROM[20239] <= 32'b00000000010000010000000100010011;
ROM[20240] <= 32'b00000000010100010010000000100011;
ROM[20241] <= 32'b00000000010000010000000100010011;
ROM[20242] <= 32'b00000000011000010010000000100011;
ROM[20243] <= 32'b00000000010000010000000100010011;
ROM[20244] <= 32'b00000001010000000000001110010011;
ROM[20245] <= 32'b00000000010000111000001110010011;
ROM[20246] <= 32'b01000000011100010000001110110011;
ROM[20247] <= 32'b00000000011100000000001000110011;
ROM[20248] <= 32'b00000000001000000000000110110011;
ROM[20249] <= 32'b01111010110000000000000011101111;
ROM[20250] <= 32'b11111111110000010000000100010011;
ROM[20251] <= 32'b00000000000000010010001110000011;
ROM[20252] <= 32'b00000000011100011010000000100011;
ROM[20253] <= 32'b00000000000000011010001110000011;
ROM[20254] <= 32'b00000000011100010010000000100011;
ROM[20255] <= 32'b00000000010000010000000100010011;
ROM[20256] <= 32'b00000000000000000000001110010011;
ROM[20257] <= 32'b00000000011100010010000000100011;
ROM[20258] <= 32'b00000000010000010000000100010011;
ROM[20259] <= 32'b11111111110000010000000100010011;
ROM[20260] <= 32'b00000000000000010010001110000011;
ROM[20261] <= 32'b11111111110000010000000100010011;
ROM[20262] <= 32'b00000000000000010010010000000011;
ROM[20263] <= 32'b00000000011101000010010010110011;
ROM[20264] <= 32'b00000000100000111010010100110011;
ROM[20265] <= 32'b00000000101001001000001110110011;
ROM[20266] <= 32'b00000000000100111000001110010011;
ROM[20267] <= 32'b00000000000100111111001110010011;
ROM[20268] <= 32'b00000000011100010010000000100011;
ROM[20269] <= 32'b00000000010000010000000100010011;
ROM[20270] <= 32'b11111111110000010000000100010011;
ROM[20271] <= 32'b00000000000000010010001110000011;
ROM[20272] <= 32'b00000000000000111000101001100011;
ROM[20273] <= 32'b00000000000000010100001110110111;
ROM[20274] <= 32'b11111110000000111000001110010011;
ROM[20275] <= 32'b00000000111000111000001110110011;
ROM[20276] <= 32'b00000000000000111000000011100111;
ROM[20277] <= 32'b00000000000000011010001110000011;
ROM[20278] <= 32'b00000000011100010010000000100011;
ROM[20279] <= 32'b00000000010000010000000100010011;
ROM[20280] <= 32'b00000000000000011010001110000011;
ROM[20281] <= 32'b00000000011100010010000000100011;
ROM[20282] <= 32'b00000000010000010000000100010011;
ROM[20283] <= 32'b00000110000001101010001110000011;
ROM[20284] <= 32'b00000000011100010010000000100011;
ROM[20285] <= 32'b00000000010000010000000100010011;
ROM[20286] <= 32'b11111111110000010000000100010011;
ROM[20287] <= 32'b00000000000000010010001110000011;
ROM[20288] <= 32'b11111111110000010000000100010011;
ROM[20289] <= 32'b00000000000000010010010000000011;
ROM[20290] <= 32'b00000000011101000000001110110011;
ROM[20291] <= 32'b00000000011100010010000000100011;
ROM[20292] <= 32'b00000000010000010000000100010011;
ROM[20293] <= 32'b11111111110000010000000100010011;
ROM[20294] <= 32'b00000000000000010010001110000011;
ROM[20295] <= 32'b00000000000000111000001100010011;
ROM[20296] <= 32'b00000000110100110000010000110011;
ROM[20297] <= 32'b00000000000001000010001110000011;
ROM[20298] <= 32'b00000000011100010010000000100011;
ROM[20299] <= 32'b00000000010000010000000100010011;
ROM[20300] <= 32'b11111111110000010000000100010011;
ROM[20301] <= 32'b00000000000000010010001110000011;
ROM[20302] <= 32'b11111111110000010000000100010011;
ROM[20303] <= 32'b00000000000000010010010000000011;
ROM[20304] <= 32'b01000000011101000000001110110011;
ROM[20305] <= 32'b00000000011100010010000000100011;
ROM[20306] <= 32'b00000000010000010000000100010011;
ROM[20307] <= 32'b00000000000000100010001110000011;
ROM[20308] <= 32'b00000000011100010010000000100011;
ROM[20309] <= 32'b00000000010000010000000100010011;
ROM[20310] <= 32'b11111111110000010000000100010011;
ROM[20311] <= 32'b00000000000000010010001110000011;
ROM[20312] <= 32'b11111111110000010000000100010011;
ROM[20313] <= 32'b00000000000000010010010000000011;
ROM[20314] <= 32'b00000000011101000010010010110011;
ROM[20315] <= 32'b00000000100000111010010100110011;
ROM[20316] <= 32'b00000000101001001000001110110011;
ROM[20317] <= 32'b00000000000100111000001110010011;
ROM[20318] <= 32'b00000000000100111111001110010011;
ROM[20319] <= 32'b00000000011100010010000000100011;
ROM[20320] <= 32'b00000000010000010000000100010011;
ROM[20321] <= 32'b11111111110000010000000100010011;
ROM[20322] <= 32'b00000000000000010010001110000011;
ROM[20323] <= 32'b00000000000000111000101001100011;
ROM[20324] <= 32'b00000000000000010100001110110111;
ROM[20325] <= 32'b11101111110000111000001110010011;
ROM[20326] <= 32'b00000000111000111000001110110011;
ROM[20327] <= 32'b00000000000000111000000011100111;
ROM[20328] <= 32'b00000000100000011010001110000011;
ROM[20329] <= 32'b00000000011100010010000000100011;
ROM[20330] <= 32'b00000000010000010000000100010011;
ROM[20331] <= 32'b00000000000000100010001110000011;
ROM[20332] <= 32'b00000000011100010010000000100011;
ROM[20333] <= 32'b00000000010000010000000100010011;
ROM[20334] <= 32'b00000110000001101010001110000011;
ROM[20335] <= 32'b00000000011100010010000000100011;
ROM[20336] <= 32'b00000000010000010000000100010011;
ROM[20337] <= 32'b11111111110000010000000100010011;
ROM[20338] <= 32'b00000000000000010010001110000011;
ROM[20339] <= 32'b11111111110000010000000100010011;
ROM[20340] <= 32'b00000000000000010010010000000011;
ROM[20341] <= 32'b00000000011101000000001110110011;
ROM[20342] <= 32'b00000000011100010010000000100011;
ROM[20343] <= 32'b00000000010000010000000100010011;
ROM[20344] <= 32'b11111111110000010000000100010011;
ROM[20345] <= 32'b00000000000000010010001110000011;
ROM[20346] <= 32'b00000000000000111000001100010011;
ROM[20347] <= 32'b11111111110000010000000100010011;
ROM[20348] <= 32'b00000000000000010010001110000011;
ROM[20349] <= 32'b00000000110100110000010000110011;
ROM[20350] <= 32'b00000000011101000010000000100011;
ROM[20351] <= 32'b00000000000000011010001110000011;
ROM[20352] <= 32'b00000000011100010010000000100011;
ROM[20353] <= 32'b00000000010000010000000100010011;
ROM[20354] <= 32'b00000110010001101010001110000011;
ROM[20355] <= 32'b00000000011100010010000000100011;
ROM[20356] <= 32'b00000000010000010000000100010011;
ROM[20357] <= 32'b11111111110000010000000100010011;
ROM[20358] <= 32'b00000000000000010010001110000011;
ROM[20359] <= 32'b11111111110000010000000100010011;
ROM[20360] <= 32'b00000000000000010010010000000011;
ROM[20361] <= 32'b00000000011101000000001110110011;
ROM[20362] <= 32'b00000000011100010010000000100011;
ROM[20363] <= 32'b00000000010000010000000100010011;
ROM[20364] <= 32'b11111111110000010000000100010011;
ROM[20365] <= 32'b00000000000000010010001110000011;
ROM[20366] <= 32'b00000000000000111000001100010011;
ROM[20367] <= 32'b00000000110100110000010000110011;
ROM[20368] <= 32'b00000000000001000010001110000011;
ROM[20369] <= 32'b00000000011100010010000000100011;
ROM[20370] <= 32'b00000000010000010000000100010011;
ROM[20371] <= 32'b00000000000000100010001110000011;
ROM[20372] <= 32'b00000000011100010010000000100011;
ROM[20373] <= 32'b00000000010000010000000100010011;
ROM[20374] <= 32'b00000110010001101010001110000011;
ROM[20375] <= 32'b00000000011100010010000000100011;
ROM[20376] <= 32'b00000000010000010000000100010011;
ROM[20377] <= 32'b11111111110000010000000100010011;
ROM[20378] <= 32'b00000000000000010010001110000011;
ROM[20379] <= 32'b11111111110000010000000100010011;
ROM[20380] <= 32'b00000000000000010010010000000011;
ROM[20381] <= 32'b00000000011101000000001110110011;
ROM[20382] <= 32'b00000000011100010010000000100011;
ROM[20383] <= 32'b00000000010000010000000100010011;
ROM[20384] <= 32'b11111111110000010000000100010011;
ROM[20385] <= 32'b00000000000000010010001110000011;
ROM[20386] <= 32'b00000000000000111000001100010011;
ROM[20387] <= 32'b11111111110000010000000100010011;
ROM[20388] <= 32'b00000000000000010010001110000011;
ROM[20389] <= 32'b00000000110100110000010000110011;
ROM[20390] <= 32'b00000000011101000010000000100011;
ROM[20391] <= 32'b00000000000000100010001110000011;
ROM[20392] <= 32'b00000000011100010010000000100011;
ROM[20393] <= 32'b00000000010000010000000100010011;
ROM[20394] <= 32'b00000000000000011010001110000011;
ROM[20395] <= 32'b00000000011100010010000000100011;
ROM[20396] <= 32'b00000000010000010000000100010011;
ROM[20397] <= 32'b00000110010001101010001110000011;
ROM[20398] <= 32'b00000000011100010010000000100011;
ROM[20399] <= 32'b00000000010000010000000100010011;
ROM[20400] <= 32'b11111111110000010000000100010011;
ROM[20401] <= 32'b00000000000000010010001110000011;
ROM[20402] <= 32'b11111111110000010000000100010011;
ROM[20403] <= 32'b00000000000000010010010000000011;
ROM[20404] <= 32'b00000000011101000000001110110011;
ROM[20405] <= 32'b00000000011100010010000000100011;
ROM[20406] <= 32'b00000000010000010000000100010011;
ROM[20407] <= 32'b11111111110000010000000100010011;
ROM[20408] <= 32'b00000000000000010010001110000011;
ROM[20409] <= 32'b00000000000000111000001100010011;
ROM[20410] <= 32'b11111111110000010000000100010011;
ROM[20411] <= 32'b00000000000000010010001110000011;
ROM[20412] <= 32'b00000000110100110000010000110011;
ROM[20413] <= 32'b00000000011101000010000000100011;
ROM[20414] <= 32'b00001110010000000000000011101111;
ROM[20415] <= 32'b00000000000000011010001110000011;
ROM[20416] <= 32'b00000000011100010010000000100011;
ROM[20417] <= 32'b00000000010000010000000100010011;
ROM[20418] <= 32'b00000110000001101010001110000011;
ROM[20419] <= 32'b00000000011100010010000000100011;
ROM[20420] <= 32'b00000000010000010000000100010011;
ROM[20421] <= 32'b11111111110000010000000100010011;
ROM[20422] <= 32'b00000000000000010010001110000011;
ROM[20423] <= 32'b11111111110000010000000100010011;
ROM[20424] <= 32'b00000000000000010010010000000011;
ROM[20425] <= 32'b00000000011101000000001110110011;
ROM[20426] <= 32'b00000000011100010010000000100011;
ROM[20427] <= 32'b00000000010000010000000100010011;
ROM[20428] <= 32'b11111111110000010000000100010011;
ROM[20429] <= 32'b00000000000000010010001110000011;
ROM[20430] <= 32'b00000000000000111000001100010011;
ROM[20431] <= 32'b00000000110100110000010000110011;
ROM[20432] <= 32'b00000000000001000010001110000011;
ROM[20433] <= 32'b00000000011100010010000000100011;
ROM[20434] <= 32'b00000000010000010000000100010011;
ROM[20435] <= 32'b00000000100000011010001110000011;
ROM[20436] <= 32'b00000000011100010010000000100011;
ROM[20437] <= 32'b00000000010000010000000100010011;
ROM[20438] <= 32'b11111111110000010000000100010011;
ROM[20439] <= 32'b00000000000000010010001110000011;
ROM[20440] <= 32'b11111111110000010000000100010011;
ROM[20441] <= 32'b00000000000000010010010000000011;
ROM[20442] <= 32'b00000000011101000000001110110011;
ROM[20443] <= 32'b00000000011100010010000000100011;
ROM[20444] <= 32'b00000000010000010000000100010011;
ROM[20445] <= 32'b00000000000000011010001110000011;
ROM[20446] <= 32'b00000000011100010010000000100011;
ROM[20447] <= 32'b00000000010000010000000100010011;
ROM[20448] <= 32'b00000110000001101010001110000011;
ROM[20449] <= 32'b00000000011100010010000000100011;
ROM[20450] <= 32'b00000000010000010000000100010011;
ROM[20451] <= 32'b11111111110000010000000100010011;
ROM[20452] <= 32'b00000000000000010010001110000011;
ROM[20453] <= 32'b11111111110000010000000100010011;
ROM[20454] <= 32'b00000000000000010010010000000011;
ROM[20455] <= 32'b00000000011101000000001110110011;
ROM[20456] <= 32'b00000000011100010010000000100011;
ROM[20457] <= 32'b00000000010000010000000100010011;
ROM[20458] <= 32'b11111111110000010000000100010011;
ROM[20459] <= 32'b00000000000000010010001110000011;
ROM[20460] <= 32'b00000000000000111000001100010011;
ROM[20461] <= 32'b11111111110000010000000100010011;
ROM[20462] <= 32'b00000000000000010010001110000011;
ROM[20463] <= 32'b00000000110100110000010000110011;
ROM[20464] <= 32'b00000000011101000010000000100011;
ROM[20465] <= 32'b00000000000000011010001110000011;
ROM[20466] <= 32'b00000000011100010010000000100011;
ROM[20467] <= 32'b00000000010000010000000100010011;
ROM[20468] <= 32'b11111111110000010000000100010011;
ROM[20469] <= 32'b00000000000000010010001110000011;
ROM[20470] <= 32'b00000000011100100010000000100011;
ROM[20471] <= 32'b00001101010000000000000011101111;
ROM[20472] <= 32'b00000000100000011010001110000011;
ROM[20473] <= 32'b00000000011100010010000000100011;
ROM[20474] <= 32'b00000000010000010000000100010011;
ROM[20475] <= 32'b00000000000000100010001110000011;
ROM[20476] <= 32'b00000000011100010010000000100011;
ROM[20477] <= 32'b00000000010000010000000100010011;
ROM[20478] <= 32'b00000110000001101010001110000011;
ROM[20479] <= 32'b00000000011100010010000000100011;
ROM[20480] <= 32'b00000000010000010000000100010011;
ROM[20481] <= 32'b11111111110000010000000100010011;
ROM[20482] <= 32'b00000000000000010010001110000011;
ROM[20483] <= 32'b11111111110000010000000100010011;
ROM[20484] <= 32'b00000000000000010010010000000011;
ROM[20485] <= 32'b00000000011101000000001110110011;
ROM[20486] <= 32'b00000000011100010010000000100011;
ROM[20487] <= 32'b00000000010000010000000100010011;
ROM[20488] <= 32'b11111111110000010000000100010011;
ROM[20489] <= 32'b00000000000000010010001110000011;
ROM[20490] <= 32'b00000000000000111000001100010011;
ROM[20491] <= 32'b11111111110000010000000100010011;
ROM[20492] <= 32'b00000000000000010010001110000011;
ROM[20493] <= 32'b00000000110100110000010000110011;
ROM[20494] <= 32'b00000000011101000010000000100011;
ROM[20495] <= 32'b00000101110001101010001110000011;
ROM[20496] <= 32'b00000000011100010010000000100011;
ROM[20497] <= 32'b00000000010000010000000100010011;
ROM[20498] <= 32'b00000000000000100010001110000011;
ROM[20499] <= 32'b00000000011100010010000000100011;
ROM[20500] <= 32'b00000000010000010000000100010011;
ROM[20501] <= 32'b00000110010001101010001110000011;
ROM[20502] <= 32'b00000000011100010010000000100011;
ROM[20503] <= 32'b00000000010000010000000100010011;
ROM[20504] <= 32'b11111111110000010000000100010011;
ROM[20505] <= 32'b00000000000000010010001110000011;
ROM[20506] <= 32'b11111111110000010000000100010011;
ROM[20507] <= 32'b00000000000000010010010000000011;
ROM[20508] <= 32'b00000000011101000000001110110011;
ROM[20509] <= 32'b00000000011100010010000000100011;
ROM[20510] <= 32'b00000000010000010000000100010011;
ROM[20511] <= 32'b11111111110000010000000100010011;
ROM[20512] <= 32'b00000000000000010010001110000011;
ROM[20513] <= 32'b00000000000000111000001100010011;
ROM[20514] <= 32'b11111111110000010000000100010011;
ROM[20515] <= 32'b00000000000000010010001110000011;
ROM[20516] <= 32'b00000000110100110000010000110011;
ROM[20517] <= 32'b00000000011101000010000000100011;
ROM[20518] <= 32'b00000000000000100010001110000011;
ROM[20519] <= 32'b00000000011100010010000000100011;
ROM[20520] <= 32'b00000000010000010000000100010011;
ROM[20521] <= 32'b11111111110000010000000100010011;
ROM[20522] <= 32'b00000000000000010010001110000011;
ROM[20523] <= 32'b00000100011101101010111000100011;
ROM[20524] <= 32'b00000000000000100010001110000011;
ROM[20525] <= 32'b00000000011100010010000000100011;
ROM[20526] <= 32'b00000000010000010000000100010011;
ROM[20527] <= 32'b00000000000000100010001110000011;
ROM[20528] <= 32'b00000000011100010010000000100011;
ROM[20529] <= 32'b00000000010000010000000100010011;
ROM[20530] <= 32'b00000110000001101010001110000011;
ROM[20531] <= 32'b00000000011100010010000000100011;
ROM[20532] <= 32'b00000000010000010000000100010011;
ROM[20533] <= 32'b11111111110000010000000100010011;
ROM[20534] <= 32'b00000000000000010010001110000011;
ROM[20535] <= 32'b11111111110000010000000100010011;
ROM[20536] <= 32'b00000000000000010010010000000011;
ROM[20537] <= 32'b00000000011101000000001110110011;
ROM[20538] <= 32'b00000000011100010010000000100011;
ROM[20539] <= 32'b00000000010000010000000100010011;
ROM[20540] <= 32'b11111111110000010000000100010011;
ROM[20541] <= 32'b00000000000000010010001110000011;
ROM[20542] <= 32'b00000000000000111000001100010011;
ROM[20543] <= 32'b00000000110100110000010000110011;
ROM[20544] <= 32'b00000000000001000010001110000011;
ROM[20545] <= 32'b00000000011100010010000000100011;
ROM[20546] <= 32'b00000000010000010000000100010011;
ROM[20547] <= 32'b11111111110000010000000100010011;
ROM[20548] <= 32'b00000000000000010010001110000011;
ROM[20549] <= 32'b11111111110000010000000100010011;
ROM[20550] <= 32'b00000000000000010010010000000011;
ROM[20551] <= 32'b01000000011101000000001110110011;
ROM[20552] <= 32'b00000000011100010010000000100011;
ROM[20553] <= 32'b00000000010000010000000100010011;
ROM[20554] <= 32'b00000000000000100010001110000011;
ROM[20555] <= 32'b00000000011100010010000000100011;
ROM[20556] <= 32'b00000000010000010000000100010011;
ROM[20557] <= 32'b00000110010001101010001110000011;
ROM[20558] <= 32'b00000000011100010010000000100011;
ROM[20559] <= 32'b00000000010000010000000100010011;
ROM[20560] <= 32'b11111111110000010000000100010011;
ROM[20561] <= 32'b00000000000000010010001110000011;
ROM[20562] <= 32'b11111111110000010000000100010011;
ROM[20563] <= 32'b00000000000000010010010000000011;
ROM[20564] <= 32'b00000000011101000000001110110011;
ROM[20565] <= 32'b00000000011100010010000000100011;
ROM[20566] <= 32'b00000000010000010000000100010011;
ROM[20567] <= 32'b11111111110000010000000100010011;
ROM[20568] <= 32'b00000000000000010010001110000011;
ROM[20569] <= 32'b00000000000000111000001100010011;
ROM[20570] <= 32'b00000000110100110000010000110011;
ROM[20571] <= 32'b00000000000001000010001110000011;
ROM[20572] <= 32'b00000000011100010010000000100011;
ROM[20573] <= 32'b00000000010000010000000100010011;
ROM[20574] <= 32'b11111111110000010000000100010011;
ROM[20575] <= 32'b00000000000000010010001110000011;
ROM[20576] <= 32'b11111111110000010000000100010011;
ROM[20577] <= 32'b00000000000000010010010000000011;
ROM[20578] <= 32'b00000000011101000010010010110011;
ROM[20579] <= 32'b00000000100000111010010100110011;
ROM[20580] <= 32'b00000000101001001000001110110011;
ROM[20581] <= 32'b00000000000100111000001110010011;
ROM[20582] <= 32'b00000000000100111111001110010011;
ROM[20583] <= 32'b00000000011100010010000000100011;
ROM[20584] <= 32'b00000000010000010000000100010011;
ROM[20585] <= 32'b11111111110000010000000100010011;
ROM[20586] <= 32'b00000000000000010010001110000011;
ROM[20587] <= 32'b00000000000000111000101001100011;
ROM[20588] <= 32'b00000000000000010100001110110111;
ROM[20589] <= 32'b00011100010000111000001110010011;
ROM[20590] <= 32'b00000000111000111000001110110011;
ROM[20591] <= 32'b00000000000000111000000011100111;
ROM[20592] <= 32'b00100000110000000000000011101111;
ROM[20593] <= 32'b00000000000000100010001110000011;
ROM[20594] <= 32'b00000000011100010010000000100011;
ROM[20595] <= 32'b00000000010000010000000100010011;
ROM[20596] <= 32'b00000110010001101010001110000011;
ROM[20597] <= 32'b00000000011100010010000000100011;
ROM[20598] <= 32'b00000000010000010000000100010011;
ROM[20599] <= 32'b11111111110000010000000100010011;
ROM[20600] <= 32'b00000000000000010010001110000011;
ROM[20601] <= 32'b11111111110000010000000100010011;
ROM[20602] <= 32'b00000000000000010010010000000011;
ROM[20603] <= 32'b00000000011101000000001110110011;
ROM[20604] <= 32'b00000000011100010010000000100011;
ROM[20605] <= 32'b00000000010000010000000100010011;
ROM[20606] <= 32'b11111111110000010000000100010011;
ROM[20607] <= 32'b00000000000000010010001110000011;
ROM[20608] <= 32'b00000000000000111000001100010011;
ROM[20609] <= 32'b00000000110100110000010000110011;
ROM[20610] <= 32'b00000000000001000010001110000011;
ROM[20611] <= 32'b00000000011100010010000000100011;
ROM[20612] <= 32'b00000000010000010000000100010011;
ROM[20613] <= 32'b11111111110000010000000100010011;
ROM[20614] <= 32'b00000000000000010010001110000011;
ROM[20615] <= 32'b00000000011100011010001000100011;
ROM[20616] <= 32'b00000000000000100010001110000011;
ROM[20617] <= 32'b00000000011100010010000000100011;
ROM[20618] <= 32'b00000000010000010000000100010011;
ROM[20619] <= 32'b00000110000001101010001110000011;
ROM[20620] <= 32'b00000000011100010010000000100011;
ROM[20621] <= 32'b00000000010000010000000100010011;
ROM[20622] <= 32'b11111111110000010000000100010011;
ROM[20623] <= 32'b00000000000000010010001110000011;
ROM[20624] <= 32'b11111111110000010000000100010011;
ROM[20625] <= 32'b00000000000000010010010000000011;
ROM[20626] <= 32'b00000000011101000000001110110011;
ROM[20627] <= 32'b00000000011100010010000000100011;
ROM[20628] <= 32'b00000000010000010000000100010011;
ROM[20629] <= 32'b11111111110000010000000100010011;
ROM[20630] <= 32'b00000000000000010010001110000011;
ROM[20631] <= 32'b00000000000000111000001100010011;
ROM[20632] <= 32'b00000000110100110000010000110011;
ROM[20633] <= 32'b00000000000001000010001110000011;
ROM[20634] <= 32'b00000000011100010010000000100011;
ROM[20635] <= 32'b00000000010000010000000100010011;
ROM[20636] <= 32'b00000000010000011010001110000011;
ROM[20637] <= 32'b00000000011100010010000000100011;
ROM[20638] <= 32'b00000000010000010000000100010011;
ROM[20639] <= 32'b00000110000001101010001110000011;
ROM[20640] <= 32'b00000000011100010010000000100011;
ROM[20641] <= 32'b00000000010000010000000100010011;
ROM[20642] <= 32'b11111111110000010000000100010011;
ROM[20643] <= 32'b00000000000000010010001110000011;
ROM[20644] <= 32'b11111111110000010000000100010011;
ROM[20645] <= 32'b00000000000000010010010000000011;
ROM[20646] <= 32'b00000000011101000000001110110011;
ROM[20647] <= 32'b00000000011100010010000000100011;
ROM[20648] <= 32'b00000000010000010000000100010011;
ROM[20649] <= 32'b11111111110000010000000100010011;
ROM[20650] <= 32'b00000000000000010010001110000011;
ROM[20651] <= 32'b00000000000000111000001100010011;
ROM[20652] <= 32'b00000000110100110000010000110011;
ROM[20653] <= 32'b00000000000001000010001110000011;
ROM[20654] <= 32'b00000000011100010010000000100011;
ROM[20655] <= 32'b00000000010000010000000100010011;
ROM[20656] <= 32'b11111111110000010000000100010011;
ROM[20657] <= 32'b00000000000000010010001110000011;
ROM[20658] <= 32'b11111111110000010000000100010011;
ROM[20659] <= 32'b00000000000000010010010000000011;
ROM[20660] <= 32'b00000000011101000000001110110011;
ROM[20661] <= 32'b00000000011100010010000000100011;
ROM[20662] <= 32'b00000000010000010000000100010011;
ROM[20663] <= 32'b00000000000000100010001110000011;
ROM[20664] <= 32'b00000000011100010010000000100011;
ROM[20665] <= 32'b00000000010000010000000100010011;
ROM[20666] <= 32'b00000110000001101010001110000011;
ROM[20667] <= 32'b00000000011100010010000000100011;
ROM[20668] <= 32'b00000000010000010000000100010011;
ROM[20669] <= 32'b11111111110000010000000100010011;
ROM[20670] <= 32'b00000000000000010010001110000011;
ROM[20671] <= 32'b11111111110000010000000100010011;
ROM[20672] <= 32'b00000000000000010010010000000011;
ROM[20673] <= 32'b00000000011101000000001110110011;
ROM[20674] <= 32'b00000000011100010010000000100011;
ROM[20675] <= 32'b00000000010000010000000100010011;
ROM[20676] <= 32'b11111111110000010000000100010011;
ROM[20677] <= 32'b00000000000000010010001110000011;
ROM[20678] <= 32'b00000000000000111000001100010011;
ROM[20679] <= 32'b11111111110000010000000100010011;
ROM[20680] <= 32'b00000000000000010010001110000011;
ROM[20681] <= 32'b00000000110100110000010000110011;
ROM[20682] <= 32'b00000000011101000010000000100011;
ROM[20683] <= 32'b00000000010000011010001110000011;
ROM[20684] <= 32'b00000000011100010010000000100011;
ROM[20685] <= 32'b00000000010000010000000100010011;
ROM[20686] <= 32'b00000110010001101010001110000011;
ROM[20687] <= 32'b00000000011100010010000000100011;
ROM[20688] <= 32'b00000000010000010000000100010011;
ROM[20689] <= 32'b11111111110000010000000100010011;
ROM[20690] <= 32'b00000000000000010010001110000011;
ROM[20691] <= 32'b11111111110000010000000100010011;
ROM[20692] <= 32'b00000000000000010010010000000011;
ROM[20693] <= 32'b00000000011101000000001110110011;
ROM[20694] <= 32'b00000000011100010010000000100011;
ROM[20695] <= 32'b00000000010000010000000100010011;
ROM[20696] <= 32'b11111111110000010000000100010011;
ROM[20697] <= 32'b00000000000000010010001110000011;
ROM[20698] <= 32'b00000000000000111000001100010011;
ROM[20699] <= 32'b00000000110100110000010000110011;
ROM[20700] <= 32'b00000000000001000010001110000011;
ROM[20701] <= 32'b00000000011100010010000000100011;
ROM[20702] <= 32'b00000000010000010000000100010011;
ROM[20703] <= 32'b00000000000000100010001110000011;
ROM[20704] <= 32'b00000000011100010010000000100011;
ROM[20705] <= 32'b00000000010000010000000100010011;
ROM[20706] <= 32'b00000110010001101010001110000011;
ROM[20707] <= 32'b00000000011100010010000000100011;
ROM[20708] <= 32'b00000000010000010000000100010011;
ROM[20709] <= 32'b11111111110000010000000100010011;
ROM[20710] <= 32'b00000000000000010010001110000011;
ROM[20711] <= 32'b11111111110000010000000100010011;
ROM[20712] <= 32'b00000000000000010010010000000011;
ROM[20713] <= 32'b00000000011101000000001110110011;
ROM[20714] <= 32'b00000000011100010010000000100011;
ROM[20715] <= 32'b00000000010000010000000100010011;
ROM[20716] <= 32'b11111111110000010000000100010011;
ROM[20717] <= 32'b00000000000000010010001110000011;
ROM[20718] <= 32'b00000000000000111000001100010011;
ROM[20719] <= 32'b11111111110000010000000100010011;
ROM[20720] <= 32'b00000000000000010010001110000011;
ROM[20721] <= 32'b00000000110100110000010000110011;
ROM[20722] <= 32'b00000000011101000010000000100011;
ROM[20723] <= 32'b00000000000000000000001110010011;
ROM[20724] <= 32'b00000000011100010010000000100011;
ROM[20725] <= 32'b00000000010000010000000100010011;
ROM[20726] <= 32'b00000001010000000000001110010011;
ROM[20727] <= 32'b01000000011100011000001110110011;
ROM[20728] <= 32'b00000000000000111010000010000011;
ROM[20729] <= 32'b11111111110000010000000100010011;
ROM[20730] <= 32'b00000000000000010010001110000011;
ROM[20731] <= 32'b00000000011100100010000000100011;
ROM[20732] <= 32'b00000000010000100000000100010011;
ROM[20733] <= 32'b00000001010000000000001110010011;
ROM[20734] <= 32'b01000000011100011000001110110011;
ROM[20735] <= 32'b00000000010000111010000110000011;
ROM[20736] <= 32'b00000000100000111010001000000011;
ROM[20737] <= 32'b00000000110000111010001010000011;
ROM[20738] <= 32'b00000001000000111010001100000011;
ROM[20739] <= 32'b00000000000000001000000011100111;
ROM[20740] <= 32'b00000000000000010010000000100011;
ROM[20741] <= 32'b00000000010000010000000100010011;
ROM[20742] <= 32'b00000101110001101010001110000011;
ROM[20743] <= 32'b00000000011100010010000000100011;
ROM[20744] <= 32'b00000000010000010000000100010011;
ROM[20745] <= 32'b00000000000000100010001110000011;
ROM[20746] <= 32'b00000000011100010010000000100011;
ROM[20747] <= 32'b00000000010000010000000100010011;
ROM[20748] <= 32'b11111111110000010000000100010011;
ROM[20749] <= 32'b00000000000000010010001110000011;
ROM[20750] <= 32'b11111111110000010000000100010011;
ROM[20751] <= 32'b00000000000000010010010000000011;
ROM[20752] <= 32'b00000000011101000010001110110011;
ROM[20753] <= 32'b00000000011100010010000000100011;
ROM[20754] <= 32'b00000000010000010000000100010011;
ROM[20755] <= 32'b11111111110000010000000100010011;
ROM[20756] <= 32'b00000000000000010010001110000011;
ROM[20757] <= 32'b00000000000000111000101001100011;
ROM[20758] <= 32'b00000000000000010100001110110111;
ROM[20759] <= 32'b01000110110000111000001110010011;
ROM[20760] <= 32'b00000000111000111000001110110011;
ROM[20761] <= 32'b00000000000000111000000011100111;
ROM[20762] <= 32'b00000100100000000000000011101111;
ROM[20763] <= 32'b00000000000000000000001110010011;
ROM[20764] <= 32'b00000000011100010010000000100011;
ROM[20765] <= 32'b00000000010000010000000100010011;
ROM[20766] <= 32'b00000001010000000000001110010011;
ROM[20767] <= 32'b01000000011100011000001110110011;
ROM[20768] <= 32'b00000000000000111010000010000011;
ROM[20769] <= 32'b11111111110000010000000100010011;
ROM[20770] <= 32'b00000000000000010010001110000011;
ROM[20771] <= 32'b00000000011100100010000000100011;
ROM[20772] <= 32'b00000000010000100000000100010011;
ROM[20773] <= 32'b00000001010000000000001110010011;
ROM[20774] <= 32'b01000000011100011000001110110011;
ROM[20775] <= 32'b00000000010000111010000110000011;
ROM[20776] <= 32'b00000000100000111010001000000011;
ROM[20777] <= 32'b00000000110000111010001010000011;
ROM[20778] <= 32'b00000001000000111010001100000011;
ROM[20779] <= 32'b00000000000000001000000011100111;
ROM[20780] <= 32'b00000101110001101010001110000011;
ROM[20781] <= 32'b00000000011100010010000000100011;
ROM[20782] <= 32'b00000000010000010000000100010011;
ROM[20783] <= 32'b11111111110000010000000100010011;
ROM[20784] <= 32'b00000000000000010010001110000011;
ROM[20785] <= 32'b00000000011100011010000000100011;
ROM[20786] <= 32'b00000000000000011010001110000011;
ROM[20787] <= 32'b00000000011100010010000000100011;
ROM[20788] <= 32'b00000000010000010000000100010011;
ROM[20789] <= 32'b00000110010001101010001110000011;
ROM[20790] <= 32'b00000000011100010010000000100011;
ROM[20791] <= 32'b00000000010000010000000100010011;
ROM[20792] <= 32'b11111111110000010000000100010011;
ROM[20793] <= 32'b00000000000000010010001110000011;
ROM[20794] <= 32'b11111111110000010000000100010011;
ROM[20795] <= 32'b00000000000000010010010000000011;
ROM[20796] <= 32'b00000000011101000000001110110011;
ROM[20797] <= 32'b00000000011100010010000000100011;
ROM[20798] <= 32'b00000000010000010000000100010011;
ROM[20799] <= 32'b11111111110000010000000100010011;
ROM[20800] <= 32'b00000000000000010010001110000011;
ROM[20801] <= 32'b00000000000000111000001100010011;
ROM[20802] <= 32'b00000000110100110000010000110011;
ROM[20803] <= 32'b00000000000001000010001110000011;
ROM[20804] <= 32'b00000000011100010010000000100011;
ROM[20805] <= 32'b00000000010000010000000100010011;
ROM[20806] <= 32'b00000000000000000000001110010011;
ROM[20807] <= 32'b00000000011100010010000000100011;
ROM[20808] <= 32'b00000000010000010000000100010011;
ROM[20809] <= 32'b11111111110000010000000100010011;
ROM[20810] <= 32'b00000000000000010010001110000011;
ROM[20811] <= 32'b11111111110000010000000100010011;
ROM[20812] <= 32'b00000000000000010010010000000011;
ROM[20813] <= 32'b00000000011101000010010010110011;
ROM[20814] <= 32'b00000000100000111010010100110011;
ROM[20815] <= 32'b00000000101001001000001110110011;
ROM[20816] <= 32'b00000000000100111000001110010011;
ROM[20817] <= 32'b00000000000100111111001110010011;
ROM[20818] <= 32'b00000000011100010010000000100011;
ROM[20819] <= 32'b00000000010000010000000100010011;
ROM[20820] <= 32'b11111111110000010000000100010011;
ROM[20821] <= 32'b00000000000000010010001110000011;
ROM[20822] <= 32'b01000000011100000000001110110011;
ROM[20823] <= 32'b00000000000100111000001110010011;
ROM[20824] <= 32'b00000000011100010010000000100011;
ROM[20825] <= 32'b00000000010000010000000100010011;
ROM[20826] <= 32'b00000000000000011010001110000011;
ROM[20827] <= 32'b00000000011100010010000000100011;
ROM[20828] <= 32'b00000000010000010000000100010011;
ROM[20829] <= 32'b00000110010001101010001110000011;
ROM[20830] <= 32'b00000000011100010010000000100011;
ROM[20831] <= 32'b00000000010000010000000100010011;
ROM[20832] <= 32'b11111111110000010000000100010011;
ROM[20833] <= 32'b00000000000000010010001110000011;
ROM[20834] <= 32'b11111111110000010000000100010011;
ROM[20835] <= 32'b00000000000000010010010000000011;
ROM[20836] <= 32'b00000000011101000000001110110011;
ROM[20837] <= 32'b00000000011100010010000000100011;
ROM[20838] <= 32'b00000000010000010000000100010011;
ROM[20839] <= 32'b11111111110000010000000100010011;
ROM[20840] <= 32'b00000000000000010010001110000011;
ROM[20841] <= 32'b00000000000000111000001100010011;
ROM[20842] <= 32'b00000000110100110000010000110011;
ROM[20843] <= 32'b00000000000001000010001110000011;
ROM[20844] <= 32'b00000000011100010010000000100011;
ROM[20845] <= 32'b00000000010000010000000100010011;
ROM[20846] <= 32'b00000000000000100010001110000011;
ROM[20847] <= 32'b00000000011100010010000000100011;
ROM[20848] <= 32'b00000000010000010000000100010011;
ROM[20849] <= 32'b11111111110000010000000100010011;
ROM[20850] <= 32'b00000000000000010010001110000011;
ROM[20851] <= 32'b11111111110000010000000100010011;
ROM[20852] <= 32'b00000000000000010010010000000011;
ROM[20853] <= 32'b00000000100000111010001110110011;
ROM[20854] <= 32'b00000000011100010010000000100011;
ROM[20855] <= 32'b00000000010000010000000100010011;
ROM[20856] <= 32'b11111111110000010000000100010011;
ROM[20857] <= 32'b00000000000000010010001110000011;
ROM[20858] <= 32'b11111111110000010000000100010011;
ROM[20859] <= 32'b00000000000000010010010000000011;
ROM[20860] <= 32'b00000000011101000111001110110011;
ROM[20861] <= 32'b00000000011100010010000000100011;
ROM[20862] <= 32'b00000000010000010000000100010011;
ROM[20863] <= 32'b11111111110000010000000100010011;
ROM[20864] <= 32'b00000000000000010010001110000011;
ROM[20865] <= 32'b01000000011100000000001110110011;
ROM[20866] <= 32'b00000000000100111000001110010011;
ROM[20867] <= 32'b00000000011100010010000000100011;
ROM[20868] <= 32'b00000000010000010000000100010011;
ROM[20869] <= 32'b11111111110000010000000100010011;
ROM[20870] <= 32'b00000000000000010010001110000011;
ROM[20871] <= 32'b00000000000000111000101001100011;
ROM[20872] <= 32'b00000000000000010100001110110111;
ROM[20873] <= 32'b01101001000000111000001110010011;
ROM[20874] <= 32'b00000000111000111000001110110011;
ROM[20875] <= 32'b00000000000000111000000011100111;
ROM[20876] <= 32'b00000000000000011010001110000011;
ROM[20877] <= 32'b00000000011100010010000000100011;
ROM[20878] <= 32'b00000000010000010000000100010011;
ROM[20879] <= 32'b00000110010001101010001110000011;
ROM[20880] <= 32'b00000000011100010010000000100011;
ROM[20881] <= 32'b00000000010000010000000100010011;
ROM[20882] <= 32'b11111111110000010000000100010011;
ROM[20883] <= 32'b00000000000000010010001110000011;
ROM[20884] <= 32'b11111111110000010000000100010011;
ROM[20885] <= 32'b00000000000000010010010000000011;
ROM[20886] <= 32'b00000000011101000000001110110011;
ROM[20887] <= 32'b00000000011100010010000000100011;
ROM[20888] <= 32'b00000000010000010000000100010011;
ROM[20889] <= 32'b11111111110000010000000100010011;
ROM[20890] <= 32'b00000000000000010010001110000011;
ROM[20891] <= 32'b00000000000000111000001100010011;
ROM[20892] <= 32'b00000000110100110000010000110011;
ROM[20893] <= 32'b00000000000001000010001110000011;
ROM[20894] <= 32'b00000000011100010010000000100011;
ROM[20895] <= 32'b00000000010000010000000100010011;
ROM[20896] <= 32'b11111111110000010000000100010011;
ROM[20897] <= 32'b00000000000000010010001110000011;
ROM[20898] <= 32'b00000000011100011010000000100011;
ROM[20899] <= 32'b11100011110111111111000011101111;
ROM[20900] <= 32'b00000000000000011010001110000011;
ROM[20901] <= 32'b00000000011100010010000000100011;
ROM[20902] <= 32'b00000000010000010000000100010011;
ROM[20903] <= 32'b00000001010000000000001110010011;
ROM[20904] <= 32'b01000000011100011000001110110011;
ROM[20905] <= 32'b00000000000000111010000010000011;
ROM[20906] <= 32'b11111111110000010000000100010011;
ROM[20907] <= 32'b00000000000000010010001110000011;
ROM[20908] <= 32'b00000000011100100010000000100011;
ROM[20909] <= 32'b00000000010000100000000100010011;
ROM[20910] <= 32'b00000001010000000000001110010011;
ROM[20911] <= 32'b01000000011100011000001110110011;
ROM[20912] <= 32'b00000000010000111010000110000011;
ROM[20913] <= 32'b00000000100000111010001000000011;
ROM[20914] <= 32'b00000000110000111010001010000011;
ROM[20915] <= 32'b00000001000000111010001100000011;
ROM[20916] <= 32'b00000000000000001000000011100111;
ROM[20917] <= 32'b00000000000000010010000000100011;
ROM[20918] <= 32'b00000000010000010000000100010011;
ROM[20919] <= 32'b00000000000000010010000000100011;
ROM[20920] <= 32'b00000000010000010000000100010011;
ROM[20921] <= 32'b00000000000000010010000000100011;
ROM[20922] <= 32'b00000000010000010000000100010011;
ROM[20923] <= 32'b00000000000000100010001110000011;
ROM[20924] <= 32'b00000000011100010010000000100011;
ROM[20925] <= 32'b00000000010000010000000100010011;
ROM[20926] <= 32'b00000000000000010100001110110111;
ROM[20927] <= 32'b01110100010000111000001110010011;
ROM[20928] <= 32'b00000000111000111000001110110011;
ROM[20929] <= 32'b00000000011100010010000000100011;
ROM[20930] <= 32'b00000000010000010000000100010011;
ROM[20931] <= 32'b00000000001100010010000000100011;
ROM[20932] <= 32'b00000000010000010000000100010011;
ROM[20933] <= 32'b00000000010000010010000000100011;
ROM[20934] <= 32'b00000000010000010000000100010011;
ROM[20935] <= 32'b00000000010100010010000000100011;
ROM[20936] <= 32'b00000000010000010000000100010011;
ROM[20937] <= 32'b00000000011000010010000000100011;
ROM[20938] <= 32'b00000000010000010000000100010011;
ROM[20939] <= 32'b00000001010000000000001110010011;
ROM[20940] <= 32'b00000000010000111000001110010011;
ROM[20941] <= 32'b01000000011100010000001110110011;
ROM[20942] <= 32'b00000000011100000000001000110011;
ROM[20943] <= 32'b00000000001000000000000110110011;
ROM[20944] <= 32'b11111111110111111110000011101111;
ROM[20945] <= 32'b11111111110000010000000100010011;
ROM[20946] <= 32'b00000000000000010010001110000011;
ROM[20947] <= 32'b00000000011100011010000000100011;
ROM[20948] <= 32'b00000000000000011010001110000011;
ROM[20949] <= 32'b00000000011100010010000000100011;
ROM[20950] <= 32'b00000000010000010000000100010011;
ROM[20951] <= 32'b00000000010000000000001110010011;
ROM[20952] <= 32'b00000000011100010010000000100011;
ROM[20953] <= 32'b00000000010000010000000100010011;
ROM[20954] <= 32'b11111111110000010000000100010011;
ROM[20955] <= 32'b00000000000000010010001110000011;
ROM[20956] <= 32'b11111111110000010000000100010011;
ROM[20957] <= 32'b00000000000000010010010000000011;
ROM[20958] <= 32'b00000000011101000000001110110011;
ROM[20959] <= 32'b00000000011100010010000000100011;
ROM[20960] <= 32'b00000000010000010000000100010011;
ROM[20961] <= 32'b11111111110000010000000100010011;
ROM[20962] <= 32'b00000000000000010010001110000011;
ROM[20963] <= 32'b00000000011100011010010000100011;
ROM[20964] <= 32'b00000000100000011010001110000011;
ROM[20965] <= 32'b00000000011100010010000000100011;
ROM[20966] <= 32'b00000000010000010000000100010011;
ROM[20967] <= 32'b11111111110000010000000100010011;
ROM[20968] <= 32'b00000000000000010010001110000011;
ROM[20969] <= 32'b00000110011101101010011000100011;
ROM[20970] <= 32'b00000000000000011010001110000011;
ROM[20971] <= 32'b00000000011100010010000000100011;
ROM[20972] <= 32'b00000000010000010000000100010011;
ROM[20973] <= 32'b00000000000000000000001110010011;
ROM[20974] <= 32'b00000000011100010010000000100011;
ROM[20975] <= 32'b00000000010000010000000100010011;
ROM[20976] <= 32'b11111111110000010000000100010011;
ROM[20977] <= 32'b00000000000000010010001110000011;
ROM[20978] <= 32'b11111111110000010000000100010011;
ROM[20979] <= 32'b00000000000000010010010000000011;
ROM[20980] <= 32'b00000000011101000010010010110011;
ROM[20981] <= 32'b00000000100000111010010100110011;
ROM[20982] <= 32'b00000000101001001000001110110011;
ROM[20983] <= 32'b00000000000100111000001110010011;
ROM[20984] <= 32'b00000000000100111111001110010011;
ROM[20985] <= 32'b00000000011100010010000000100011;
ROM[20986] <= 32'b00000000010000010000000100010011;
ROM[20987] <= 32'b11111111110000010000000100010011;
ROM[20988] <= 32'b00000000000000010010001110000011;
ROM[20989] <= 32'b01000000011100000000001110110011;
ROM[20990] <= 32'b00000000000100111000001110010011;
ROM[20991] <= 32'b00000000011100010010000000100011;
ROM[20992] <= 32'b00000000010000010000000100010011;
ROM[20993] <= 32'b11111111110000010000000100010011;
ROM[20994] <= 32'b00000000000000010010001110000011;
ROM[20995] <= 32'b00000000000000111000101001100011;
ROM[20996] <= 32'b00000000000000010101001110110111;
ROM[20997] <= 32'b10000010010000111000001110010011;
ROM[20998] <= 32'b00000000111000111000001110110011;
ROM[20999] <= 32'b00000000000000111000000011100111;
ROM[21000] <= 32'b01010001010000000000000011101111;
ROM[21001] <= 32'b00000000000000011010001110000011;
ROM[21002] <= 32'b00000000011100010010000000100011;
ROM[21003] <= 32'b00000000010000010000000100010011;
ROM[21004] <= 32'b00000110000001101010001110000011;
ROM[21005] <= 32'b00000000011100010010000000100011;
ROM[21006] <= 32'b00000000010000010000000100010011;
ROM[21007] <= 32'b11111111110000010000000100010011;
ROM[21008] <= 32'b00000000000000010010001110000011;
ROM[21009] <= 32'b11111111110000010000000100010011;
ROM[21010] <= 32'b00000000000000010010010000000011;
ROM[21011] <= 32'b00000000011101000000001110110011;
ROM[21012] <= 32'b00000000011100010010000000100011;
ROM[21013] <= 32'b00000000010000010000000100010011;
ROM[21014] <= 32'b11111111110000010000000100010011;
ROM[21015] <= 32'b00000000000000010010001110000011;
ROM[21016] <= 32'b00000000000000111000001100010011;
ROM[21017] <= 32'b00000000110100110000010000110011;
ROM[21018] <= 32'b00000000000001000010001110000011;
ROM[21019] <= 32'b00000000011100010010000000100011;
ROM[21020] <= 32'b00000000010000010000000100010011;
ROM[21021] <= 32'b00000000000000100010001110000011;
ROM[21022] <= 32'b00000000011100010010000000100011;
ROM[21023] <= 32'b00000000010000010000000100010011;
ROM[21024] <= 32'b00000000001100000000001110010011;
ROM[21025] <= 32'b00000000011100010010000000100011;
ROM[21026] <= 32'b00000000010000010000000100010011;
ROM[21027] <= 32'b11111111110000010000000100010011;
ROM[21028] <= 32'b00000000000000010010001110000011;
ROM[21029] <= 32'b11111111110000010000000100010011;
ROM[21030] <= 32'b00000000000000010010010000000011;
ROM[21031] <= 32'b00000000011101000000001110110011;
ROM[21032] <= 32'b00000000011100010010000000100011;
ROM[21033] <= 32'b00000000010000010000000100010011;
ROM[21034] <= 32'b11111111110000010000000100010011;
ROM[21035] <= 32'b00000000000000010010001110000011;
ROM[21036] <= 32'b11111111110000010000000100010011;
ROM[21037] <= 32'b00000000000000010010010000000011;
ROM[21038] <= 32'b00000000100000111010001110110011;
ROM[21039] <= 32'b00000000011100010010000000100011;
ROM[21040] <= 32'b00000000010000010000000100010011;
ROM[21041] <= 32'b11111111110000010000000100010011;
ROM[21042] <= 32'b00000000000000010010001110000011;
ROM[21043] <= 32'b00000000000000111000101001100011;
ROM[21044] <= 32'b00000000000000010101001110110111;
ROM[21045] <= 32'b10011111100000111000001110010011;
ROM[21046] <= 32'b00000000111000111000001110110011;
ROM[21047] <= 32'b00000000000000111000000011100111;
ROM[21048] <= 32'b00000000000000011010001110000011;
ROM[21049] <= 32'b00000000011100010010000000100011;
ROM[21050] <= 32'b00000000010000010000000100010011;
ROM[21051] <= 32'b00000110010001101010001110000011;
ROM[21052] <= 32'b00000000011100010010000000100011;
ROM[21053] <= 32'b00000000010000010000000100010011;
ROM[21054] <= 32'b11111111110000010000000100010011;
ROM[21055] <= 32'b00000000000000010010001110000011;
ROM[21056] <= 32'b11111111110000010000000100010011;
ROM[21057] <= 32'b00000000000000010010010000000011;
ROM[21058] <= 32'b00000000011101000000001110110011;
ROM[21059] <= 32'b00000000011100010010000000100011;
ROM[21060] <= 32'b00000000010000010000000100010011;
ROM[21061] <= 32'b11111111110000010000000100010011;
ROM[21062] <= 32'b00000000000000010010001110000011;
ROM[21063] <= 32'b00000000000000111000001100010011;
ROM[21064] <= 32'b00000000110100110000010000110011;
ROM[21065] <= 32'b00000000000001000010001110000011;
ROM[21066] <= 32'b00000000011100010010000000100011;
ROM[21067] <= 32'b00000000010000010000000100010011;
ROM[21068] <= 32'b11111111110000010000000100010011;
ROM[21069] <= 32'b00000000000000010010001110000011;
ROM[21070] <= 32'b00000000011100011010001000100011;
ROM[21071] <= 32'b00000000000000011010001110000011;
ROM[21072] <= 32'b00000000011100010010000000100011;
ROM[21073] <= 32'b00000000010000010000000100010011;
ROM[21074] <= 32'b00000110000001101010001110000011;
ROM[21075] <= 32'b00000000011100010010000000100011;
ROM[21076] <= 32'b00000000010000010000000100010011;
ROM[21077] <= 32'b11111111110000010000000100010011;
ROM[21078] <= 32'b00000000000000010010001110000011;
ROM[21079] <= 32'b11111111110000010000000100010011;
ROM[21080] <= 32'b00000000000000010010010000000011;
ROM[21081] <= 32'b00000000011101000000001110110011;
ROM[21082] <= 32'b00000000011100010010000000100011;
ROM[21083] <= 32'b00000000010000010000000100010011;
ROM[21084] <= 32'b11111111110000010000000100010011;
ROM[21085] <= 32'b00000000000000010010001110000011;
ROM[21086] <= 32'b00000000000000111000001100010011;
ROM[21087] <= 32'b00000000110100110000010000110011;
ROM[21088] <= 32'b00000000000001000010001110000011;
ROM[21089] <= 32'b00000000011100010010000000100011;
ROM[21090] <= 32'b00000000010000010000000100010011;
ROM[21091] <= 32'b00000000100000011010001110000011;
ROM[21092] <= 32'b00000000011100010010000000100011;
ROM[21093] <= 32'b00000000010000010000000100010011;
ROM[21094] <= 32'b00000110100001101010001110000011;
ROM[21095] <= 32'b00000000011100010010000000100011;
ROM[21096] <= 32'b00000000010000010000000100010011;
ROM[21097] <= 32'b11111111110000010000000100010011;
ROM[21098] <= 32'b00000000000000010010001110000011;
ROM[21099] <= 32'b11111111110000010000000100010011;
ROM[21100] <= 32'b00000000000000010010010000000011;
ROM[21101] <= 32'b00000000011101000000001110110011;
ROM[21102] <= 32'b00000000011100010010000000100011;
ROM[21103] <= 32'b00000000010000010000000100010011;
ROM[21104] <= 32'b11111111110000010000000100010011;
ROM[21105] <= 32'b00000000000000010010001110000011;
ROM[21106] <= 32'b00000000000000111000001100010011;
ROM[21107] <= 32'b11111111110000010000000100010011;
ROM[21108] <= 32'b00000000000000010010001110000011;
ROM[21109] <= 32'b00000000110100110000010000110011;
ROM[21110] <= 32'b00000000011101000010000000100011;
ROM[21111] <= 32'b00000000001000000000001110010011;
ROM[21112] <= 32'b00000000011100010010000000100011;
ROM[21113] <= 32'b00000000010000010000000100010011;
ROM[21114] <= 32'b11111111110000010000000100010011;
ROM[21115] <= 32'b00000000000000010010001110000011;
ROM[21116] <= 32'b00000110011101101010100000100011;
ROM[21117] <= 32'b00110100000000000000000011101111;
ROM[21118] <= 32'b00000000000000011010001110000011;
ROM[21119] <= 32'b00000000011100010010000000100011;
ROM[21120] <= 32'b00000000010000010000000100010011;
ROM[21121] <= 32'b00000000000000100010001110000011;
ROM[21122] <= 32'b00000000011100010010000000100011;
ROM[21123] <= 32'b00000000010000010000000100010011;
ROM[21124] <= 32'b11111111110000010000000100010011;
ROM[21125] <= 32'b00000000000000010010001110000011;
ROM[21126] <= 32'b11111111110000010000000100010011;
ROM[21127] <= 32'b00000000000000010010010000000011;
ROM[21128] <= 32'b00000000011101000000001110110011;
ROM[21129] <= 32'b00000000011100010010000000100011;
ROM[21130] <= 32'b00000000010000010000000100010011;
ROM[21131] <= 32'b00000000000000100010001110000011;
ROM[21132] <= 32'b00000000011100010010000000100011;
ROM[21133] <= 32'b00000000010000010000000100010011;
ROM[21134] <= 32'b11111111110000010000000100010011;
ROM[21135] <= 32'b00000000000000010010001110000011;
ROM[21136] <= 32'b11111111110000010000000100010011;
ROM[21137] <= 32'b00000000000000010010010000000011;
ROM[21138] <= 32'b00000000011101000000001110110011;
ROM[21139] <= 32'b00000000011100010010000000100011;
ROM[21140] <= 32'b00000000010000010000000100010011;
ROM[21141] <= 32'b00000000000000100010001110000011;
ROM[21142] <= 32'b00000000011100010010000000100011;
ROM[21143] <= 32'b00000000010000010000000100010011;
ROM[21144] <= 32'b11111111110000010000000100010011;
ROM[21145] <= 32'b00000000000000010010001110000011;
ROM[21146] <= 32'b11111111110000010000000100010011;
ROM[21147] <= 32'b00000000000000010010010000000011;
ROM[21148] <= 32'b00000000011101000000001110110011;
ROM[21149] <= 32'b00000000011100010010000000100011;
ROM[21150] <= 32'b00000000010000010000000100010011;
ROM[21151] <= 32'b00000000000000100010001110000011;
ROM[21152] <= 32'b00000000011100010010000000100011;
ROM[21153] <= 32'b00000000010000010000000100010011;
ROM[21154] <= 32'b11111111110000010000000100010011;
ROM[21155] <= 32'b00000000000000010010001110000011;
ROM[21156] <= 32'b11111111110000010000000100010011;
ROM[21157] <= 32'b00000000000000010010010000000011;
ROM[21158] <= 32'b00000000011101000000001110110011;
ROM[21159] <= 32'b00000000011100010010000000100011;
ROM[21160] <= 32'b00000000010000010000000100010011;
ROM[21161] <= 32'b00000000010000000000001110010011;
ROM[21162] <= 32'b00000000011100010010000000100011;
ROM[21163] <= 32'b00000000010000010000000100010011;
ROM[21164] <= 32'b11111111110000010000000100010011;
ROM[21165] <= 32'b00000000000000010010001110000011;
ROM[21166] <= 32'b11111111110000010000000100010011;
ROM[21167] <= 32'b00000000000000010010010000000011;
ROM[21168] <= 32'b00000000011101000000001110110011;
ROM[21169] <= 32'b00000000011100010010000000100011;
ROM[21170] <= 32'b00000000010000010000000100010011;
ROM[21171] <= 32'b11111111110000010000000100010011;
ROM[21172] <= 32'b00000000000000010010001110000011;
ROM[21173] <= 32'b00000000011100011010001000100011;
ROM[21174] <= 32'b00000000000000011010001110000011;
ROM[21175] <= 32'b00000000011100010010000000100011;
ROM[21176] <= 32'b00000000010000010000000100010011;
ROM[21177] <= 32'b00000110010001101010001110000011;
ROM[21178] <= 32'b00000000011100010010000000100011;
ROM[21179] <= 32'b00000000010000010000000100010011;
ROM[21180] <= 32'b11111111110000010000000100010011;
ROM[21181] <= 32'b00000000000000010010001110000011;
ROM[21182] <= 32'b11111111110000010000000100010011;
ROM[21183] <= 32'b00000000000000010010010000000011;
ROM[21184] <= 32'b00000000011101000000001110110011;
ROM[21185] <= 32'b00000000011100010010000000100011;
ROM[21186] <= 32'b00000000010000010000000100010011;
ROM[21187] <= 32'b11111111110000010000000100010011;
ROM[21188] <= 32'b00000000000000010010001110000011;
ROM[21189] <= 32'b00000000000000111000001100010011;
ROM[21190] <= 32'b00000000110100110000010000110011;
ROM[21191] <= 32'b00000000000001000010001110000011;
ROM[21192] <= 32'b00000000011100010010000000100011;
ROM[21193] <= 32'b00000000010000010000000100010011;
ROM[21194] <= 32'b00000000010000011010001110000011;
ROM[21195] <= 32'b00000000011100010010000000100011;
ROM[21196] <= 32'b00000000010000010000000100010011;
ROM[21197] <= 32'b00000110010001101010001110000011;
ROM[21198] <= 32'b00000000011100010010000000100011;
ROM[21199] <= 32'b00000000010000010000000100010011;
ROM[21200] <= 32'b11111111110000010000000100010011;
ROM[21201] <= 32'b00000000000000010010001110000011;
ROM[21202] <= 32'b11111111110000010000000100010011;
ROM[21203] <= 32'b00000000000000010010010000000011;
ROM[21204] <= 32'b00000000011101000000001110110011;
ROM[21205] <= 32'b00000000011100010010000000100011;
ROM[21206] <= 32'b00000000010000010000000100010011;
ROM[21207] <= 32'b11111111110000010000000100010011;
ROM[21208] <= 32'b00000000000000010010001110000011;
ROM[21209] <= 32'b00000000000000111000001100010011;
ROM[21210] <= 32'b11111111110000010000000100010011;
ROM[21211] <= 32'b00000000000000010010001110000011;
ROM[21212] <= 32'b00000000110100110000010000110011;
ROM[21213] <= 32'b00000000011101000010000000100011;
ROM[21214] <= 32'b00000000000000011010001110000011;
ROM[21215] <= 32'b00000000011100010010000000100011;
ROM[21216] <= 32'b00000000010000010000000100010011;
ROM[21217] <= 32'b00000110000001101010001110000011;
ROM[21218] <= 32'b00000000011100010010000000100011;
ROM[21219] <= 32'b00000000010000010000000100010011;
ROM[21220] <= 32'b11111111110000010000000100010011;
ROM[21221] <= 32'b00000000000000010010001110000011;
ROM[21222] <= 32'b11111111110000010000000100010011;
ROM[21223] <= 32'b00000000000000010010010000000011;
ROM[21224] <= 32'b00000000011101000000001110110011;
ROM[21225] <= 32'b00000000011100010010000000100011;
ROM[21226] <= 32'b00000000010000010000000100010011;
ROM[21227] <= 32'b11111111110000010000000100010011;
ROM[21228] <= 32'b00000000000000010010001110000011;
ROM[21229] <= 32'b00000000000000111000001100010011;
ROM[21230] <= 32'b00000000110100110000010000110011;
ROM[21231] <= 32'b00000000000001000010001110000011;
ROM[21232] <= 32'b00000000011100010010000000100011;
ROM[21233] <= 32'b00000000010000010000000100010011;
ROM[21234] <= 32'b00000000000000100010001110000011;
ROM[21235] <= 32'b00000000011100010010000000100011;
ROM[21236] <= 32'b00000000010000010000000100010011;
ROM[21237] <= 32'b11111111110000010000000100010011;
ROM[21238] <= 32'b00000000000000010010001110000011;
ROM[21239] <= 32'b11111111110000010000000100010011;
ROM[21240] <= 32'b00000000000000010010010000000011;
ROM[21241] <= 32'b01000000011101000000001110110011;
ROM[21242] <= 32'b00000000011100010010000000100011;
ROM[21243] <= 32'b00000000010000010000000100010011;
ROM[21244] <= 32'b00000000000100000000001110010011;
ROM[21245] <= 32'b00000000011100010010000000100011;
ROM[21246] <= 32'b00000000010000010000000100010011;
ROM[21247] <= 32'b11111111110000010000000100010011;
ROM[21248] <= 32'b00000000000000010010001110000011;
ROM[21249] <= 32'b11111111110000010000000100010011;
ROM[21250] <= 32'b00000000000000010010010000000011;
ROM[21251] <= 32'b01000000011101000000001110110011;
ROM[21252] <= 32'b00000000011100010010000000100011;
ROM[21253] <= 32'b00000000010000010000000100010011;
ROM[21254] <= 32'b00000000010000011010001110000011;
ROM[21255] <= 32'b00000000011100010010000000100011;
ROM[21256] <= 32'b00000000010000010000000100010011;
ROM[21257] <= 32'b00000110000001101010001110000011;
ROM[21258] <= 32'b00000000011100010010000000100011;
ROM[21259] <= 32'b00000000010000010000000100010011;
ROM[21260] <= 32'b11111111110000010000000100010011;
ROM[21261] <= 32'b00000000000000010010001110000011;
ROM[21262] <= 32'b11111111110000010000000100010011;
ROM[21263] <= 32'b00000000000000010010010000000011;
ROM[21264] <= 32'b00000000011101000000001110110011;
ROM[21265] <= 32'b00000000011100010010000000100011;
ROM[21266] <= 32'b00000000010000010000000100010011;
ROM[21267] <= 32'b11111111110000010000000100010011;
ROM[21268] <= 32'b00000000000000010010001110000011;
ROM[21269] <= 32'b00000000000000111000001100010011;
ROM[21270] <= 32'b11111111110000010000000100010011;
ROM[21271] <= 32'b00000000000000010010001110000011;
ROM[21272] <= 32'b00000000110100110000010000110011;
ROM[21273] <= 32'b00000000011101000010000000100011;
ROM[21274] <= 32'b00000000000000100010001110000011;
ROM[21275] <= 32'b00000000011100010010000000100011;
ROM[21276] <= 32'b00000000010000010000000100010011;
ROM[21277] <= 32'b00000000000100000000001110010011;
ROM[21278] <= 32'b00000000011100010010000000100011;
ROM[21279] <= 32'b00000000010000010000000100010011;
ROM[21280] <= 32'b11111111110000010000000100010011;
ROM[21281] <= 32'b00000000000000010010001110000011;
ROM[21282] <= 32'b11111111110000010000000100010011;
ROM[21283] <= 32'b00000000000000010010010000000011;
ROM[21284] <= 32'b00000000011101000000001110110011;
ROM[21285] <= 32'b00000000011100010010000000100011;
ROM[21286] <= 32'b00000000010000010000000100010011;
ROM[21287] <= 32'b00000000100000011010001110000011;
ROM[21288] <= 32'b00000000011100010010000000100011;
ROM[21289] <= 32'b00000000010000010000000100010011;
ROM[21290] <= 32'b00000110100001101010001110000011;
ROM[21291] <= 32'b00000000011100010010000000100011;
ROM[21292] <= 32'b00000000010000010000000100010011;
ROM[21293] <= 32'b11111111110000010000000100010011;
ROM[21294] <= 32'b00000000000000010010001110000011;
ROM[21295] <= 32'b11111111110000010000000100010011;
ROM[21296] <= 32'b00000000000000010010010000000011;
ROM[21297] <= 32'b00000000011101000000001110110011;
ROM[21298] <= 32'b00000000011100010010000000100011;
ROM[21299] <= 32'b00000000010000010000000100010011;
ROM[21300] <= 32'b11111111110000010000000100010011;
ROM[21301] <= 32'b00000000000000010010001110000011;
ROM[21302] <= 32'b00000000000000111000001100010011;
ROM[21303] <= 32'b11111111110000010000000100010011;
ROM[21304] <= 32'b00000000000000010010001110000011;
ROM[21305] <= 32'b00000000110100110000010000110011;
ROM[21306] <= 32'b00000000011101000010000000100011;
ROM[21307] <= 32'b00000000100000011010001110000011;
ROM[21308] <= 32'b00000000011100010010000000100011;
ROM[21309] <= 32'b00000000010000010000000100010011;
ROM[21310] <= 32'b11111111110000010000000100010011;
ROM[21311] <= 32'b00000000000000010010001110000011;
ROM[21312] <= 32'b00000110011101101010101000100011;
ROM[21313] <= 32'b00000000010000011010001110000011;
ROM[21314] <= 32'b00000000011100010010000000100011;
ROM[21315] <= 32'b00000000010000010000000100010011;
ROM[21316] <= 32'b11111111110000010000000100010011;
ROM[21317] <= 32'b00000000000000010010001110000011;
ROM[21318] <= 32'b00000100011101101010111000100011;
ROM[21319] <= 32'b00000000000100000000001110010011;
ROM[21320] <= 32'b00000000011100010010000000100011;
ROM[21321] <= 32'b00000000010000010000000100010011;
ROM[21322] <= 32'b11111111110000010000000100010011;
ROM[21323] <= 32'b00000000000000010010001110000011;
ROM[21324] <= 32'b00000110011101101010100000100011;
ROM[21325] <= 32'b00000000100000011010001110000011;
ROM[21326] <= 32'b00000000011100010010000000100011;
ROM[21327] <= 32'b00000000010000010000000100010011;
ROM[21328] <= 32'b00000001010000000000001110010011;
ROM[21329] <= 32'b01000000011100011000001110110011;
ROM[21330] <= 32'b00000000000000111010000010000011;
ROM[21331] <= 32'b11111111110000010000000100010011;
ROM[21332] <= 32'b00000000000000010010001110000011;
ROM[21333] <= 32'b00000000011100100010000000100011;
ROM[21334] <= 32'b00000000010000100000000100010011;
ROM[21335] <= 32'b00000001010000000000001110010011;
ROM[21336] <= 32'b01000000011100011000001110110011;
ROM[21337] <= 32'b00000000010000111010000110000011;
ROM[21338] <= 32'b00000000100000111010001000000011;
ROM[21339] <= 32'b00000000110000111010001010000011;
ROM[21340] <= 32'b00000001000000111010001100000011;
ROM[21341] <= 32'b00000000000000001000000011100111;
ROM[21342] <= 32'b00000000000000010010000000100011;
ROM[21343] <= 32'b00000000010000010000000100010011;
ROM[21344] <= 32'b00000000110000000000001110010011;
ROM[21345] <= 32'b00000000011100010010000000100011;
ROM[21346] <= 32'b00000000010000010000000100010011;
ROM[21347] <= 32'b00000000000000010101001110110111;
ROM[21348] <= 32'b11011101100000111000001110010011;
ROM[21349] <= 32'b00000000111000111000001110110011;
ROM[21350] <= 32'b00000000011100010010000000100011;
ROM[21351] <= 32'b00000000010000010000000100010011;
ROM[21352] <= 32'b00000000001100010010000000100011;
ROM[21353] <= 32'b00000000010000010000000100010011;
ROM[21354] <= 32'b00000000010000010010000000100011;
ROM[21355] <= 32'b00000000010000010000000100010011;
ROM[21356] <= 32'b00000000010100010010000000100011;
ROM[21357] <= 32'b00000000010000010000000100010011;
ROM[21358] <= 32'b00000000011000010010000000100011;
ROM[21359] <= 32'b00000000010000010000000100010011;
ROM[21360] <= 32'b00000001010000000000001110010011;
ROM[21361] <= 32'b00000000010000111000001110010011;
ROM[21362] <= 32'b01000000011100010000001110110011;
ROM[21363] <= 32'b00000000011100000000001000110011;
ROM[21364] <= 32'b00000000001000000000000110110011;
ROM[21365] <= 32'b10111001100011111110000011101111;
ROM[21366] <= 32'b11111111110000010000000100010011;
ROM[21367] <= 32'b00000000000000010010001110000011;
ROM[21368] <= 32'b00000000011100011010000000100011;
ROM[21369] <= 32'b00000010001000000000001110010011;
ROM[21370] <= 32'b00000000011100010010000000100011;
ROM[21371] <= 32'b00000000010000010000000100010011;
ROM[21372] <= 32'b00000000000000011010001110000011;
ROM[21373] <= 32'b00000000011100010010000000100011;
ROM[21374] <= 32'b00000000010000010000000100010011;
ROM[21375] <= 32'b00000000000000010101001110110111;
ROM[21376] <= 32'b11100100100000111000001110010011;
ROM[21377] <= 32'b00000000111000111000001110110011;
ROM[21378] <= 32'b00000000011100010010000000100011;
ROM[21379] <= 32'b00000000010000010000000100010011;
ROM[21380] <= 32'b00000000001100010010000000100011;
ROM[21381] <= 32'b00000000010000010000000100010011;
ROM[21382] <= 32'b00000000010000010010000000100011;
ROM[21383] <= 32'b00000000010000010000000100010011;
ROM[21384] <= 32'b00000000010100010010000000100011;
ROM[21385] <= 32'b00000000010000010000000100010011;
ROM[21386] <= 32'b00000000011000010010000000100011;
ROM[21387] <= 32'b00000000010000010000000100010011;
ROM[21388] <= 32'b00000001010000000000001110010011;
ROM[21389] <= 32'b00000000100000111000001110010011;
ROM[21390] <= 32'b01000000011100010000001110110011;
ROM[21391] <= 32'b00000000011100000000001000110011;
ROM[21392] <= 32'b00000000001000000000000110110011;
ROM[21393] <= 32'b10011110100111111100000011101111;
ROM[21394] <= 32'b11111111110000010000000100010011;
ROM[21395] <= 32'b00000000000000010010001110000011;
ROM[21396] <= 32'b00000000011100011010000000100011;
ROM[21397] <= 32'b00000000000000011010001110000011;
ROM[21398] <= 32'b00000000011100010010000000100011;
ROM[21399] <= 32'b00000000010000010000000100010011;
ROM[21400] <= 32'b01011000000000000000001110010011;
ROM[21401] <= 32'b00000000011100010010000000100011;
ROM[21402] <= 32'b00000000010000010000000100010011;
ROM[21403] <= 32'b11111111110000010000000100010011;
ROM[21404] <= 32'b00000000000000010010001110000011;
ROM[21405] <= 32'b11111111110000010000000100010011;
ROM[21406] <= 32'b00000000000000010010010000000011;
ROM[21407] <= 32'b00000000011101000000001110110011;
ROM[21408] <= 32'b00000000011100010010000000100011;
ROM[21409] <= 32'b00000000010000010000000100010011;
ROM[21410] <= 32'b11111111110000010000000100010011;
ROM[21411] <= 32'b00000000000000010010001110000011;
ROM[21412] <= 32'b00000000011100011010000000100011;
ROM[21413] <= 32'b00000000000000000000001110010011;
ROM[21414] <= 32'b00000000011100010010000000100011;
ROM[21415] <= 32'b00000000010000010000000100010011;
ROM[21416] <= 32'b00000000000000011010001110000011;
ROM[21417] <= 32'b00000000011100010010000000100011;
ROM[21418] <= 32'b00000000010000010000000100010011;
ROM[21419] <= 32'b11111111110000010000000100010011;
ROM[21420] <= 32'b00000000000000010010001110000011;
ROM[21421] <= 32'b11111111110000010000000100010011;
ROM[21422] <= 32'b00000000000000010010010000000011;
ROM[21423] <= 32'b01000000011101000000001110110011;
ROM[21424] <= 32'b00000000011100010010000000100011;
ROM[21425] <= 32'b00000000010000010000000100010011;
ROM[21426] <= 32'b11111111110000010000000100010011;
ROM[21427] <= 32'b00000000000000010010001110000011;
ROM[21428] <= 32'b00000110011101101010110000100011;
ROM[21429] <= 32'b00000000000000000100001110110111;
ROM[21430] <= 32'b00000000000000111000001110010011;
ROM[21431] <= 32'b00000000011100010010000000100011;
ROM[21432] <= 32'b00000000010000010000000100010011;
ROM[21433] <= 32'b11111111110000010000000100010011;
ROM[21434] <= 32'b00000000000000010010001110000011;
ROM[21435] <= 32'b00000110011101101010111000100011;
ROM[21436] <= 32'b00000000000000000000001110010011;
ROM[21437] <= 32'b00000000011100010010000000100011;
ROM[21438] <= 32'b00000000010000010000000100010011;
ROM[21439] <= 32'b11111111110000010000000100010011;
ROM[21440] <= 32'b00000000000000010010001110000011;
ROM[21441] <= 32'b00001000011101101010000000100011;
ROM[21442] <= 32'b00000000000000000000001110010011;
ROM[21443] <= 32'b00000000011100010010000000100011;
ROM[21444] <= 32'b00000000010000010000000100010011;
ROM[21445] <= 32'b11111111110000010000000100010011;
ROM[21446] <= 32'b00000000000000010010001110000011;
ROM[21447] <= 32'b00001000011101101010001000100011;
ROM[21448] <= 32'b00000000000000010101001110110111;
ROM[21449] <= 32'b11110110110000111000001110010011;
ROM[21450] <= 32'b00000000111000111000001110110011;
ROM[21451] <= 32'b00000000011100010010000000100011;
ROM[21452] <= 32'b00000000010000010000000100010011;
ROM[21453] <= 32'b00000000001100010010000000100011;
ROM[21454] <= 32'b00000000010000010000000100010011;
ROM[21455] <= 32'b00000000010000010010000000100011;
ROM[21456] <= 32'b00000000010000010000000100010011;
ROM[21457] <= 32'b00000000010100010010000000100011;
ROM[21458] <= 32'b00000000010000010000000100010011;
ROM[21459] <= 32'b00000000011000010010000000100011;
ROM[21460] <= 32'b00000000010000010000000100010011;
ROM[21461] <= 32'b00000001010000000000001110010011;
ROM[21462] <= 32'b00000000000000111000001110010011;
ROM[21463] <= 32'b01000000011100010000001110110011;
ROM[21464] <= 32'b00000000011100000000001000110011;
ROM[21465] <= 32'b00000000001000000000000110110011;
ROM[21466] <= 32'b00000101010000000000000011101111;
ROM[21467] <= 32'b11111111110000010000000100010011;
ROM[21468] <= 32'b00000000000000010010001110000011;
ROM[21469] <= 32'b00000000011101100010000000100011;
ROM[21470] <= 32'b00000000000000000000001110010011;
ROM[21471] <= 32'b00000000011100010010000000100011;
ROM[21472] <= 32'b00000000010000010000000100010011;
ROM[21473] <= 32'b00000001010000000000001110010011;
ROM[21474] <= 32'b01000000011100011000001110110011;
ROM[21475] <= 32'b00000000000000111010000010000011;
ROM[21476] <= 32'b11111111110000010000000100010011;
ROM[21477] <= 32'b00000000000000010010001110000011;
ROM[21478] <= 32'b00000000011100100010000000100011;
ROM[21479] <= 32'b00000000010000100000000100010011;
ROM[21480] <= 32'b00000001010000000000001110010011;
ROM[21481] <= 32'b01000000011100011000001110110011;
ROM[21482] <= 32'b00000000010000111010000110000011;
ROM[21483] <= 32'b00000000100000111010001000000011;
ROM[21484] <= 32'b00000000110000111010001010000011;
ROM[21485] <= 32'b00000001000000111010001100000011;
ROM[21486] <= 32'b00000000000000001000000011100111;
ROM[21487] <= 32'b00000000000000010010000000100011;
ROM[21488] <= 32'b00000000010000010000000100010011;
ROM[21489] <= 32'b00000111111100000000001110010011;
ROM[21490] <= 32'b00000000011100010010000000100011;
ROM[21491] <= 32'b00000000010000010000000100010011;
ROM[21492] <= 32'b00000000000000010101001110110111;
ROM[21493] <= 32'b00000001110000111000001110010011;
ROM[21494] <= 32'b00000000111000111000001110110011;
ROM[21495] <= 32'b00000000011100010010000000100011;
ROM[21496] <= 32'b00000000010000010000000100010011;
ROM[21497] <= 32'b00000000001100010010000000100011;
ROM[21498] <= 32'b00000000010000010000000100010011;
ROM[21499] <= 32'b00000000010000010010000000100011;
ROM[21500] <= 32'b00000000010000010000000100010011;
ROM[21501] <= 32'b00000000010100010010000000100011;
ROM[21502] <= 32'b00000000010000010000000100010011;
ROM[21503] <= 32'b00000000011000010010000000100011;
ROM[21504] <= 32'b00000000010000010000000100010011;
ROM[21505] <= 32'b00000001010000000000001110010011;
ROM[21506] <= 32'b00000000010000111000001110010011;
ROM[21507] <= 32'b01000000011100010000001110110011;
ROM[21508] <= 32'b00000000011100000000001000110011;
ROM[21509] <= 32'b00000000001000000000000110110011;
ROM[21510] <= 32'b10000110100011101011000011101111;
ROM[21511] <= 32'b11111111110000010000000100010011;
ROM[21512] <= 32'b00000000000000010010001110000011;
ROM[21513] <= 32'b00001000011101101010010000100011;
ROM[21514] <= 32'b00000000000000000000001110010011;
ROM[21515] <= 32'b00000000011100010010000000100011;
ROM[21516] <= 32'b00000000010000010000000100010011;
ROM[21517] <= 32'b00000011111100000000001110010011;
ROM[21518] <= 32'b00000000011100010010000000100011;
ROM[21519] <= 32'b00000000010000010000000100010011;
ROM[21520] <= 32'b00000011111100000000001110010011;
ROM[21521] <= 32'b00000000011100010010000000100011;
ROM[21522] <= 32'b00000000010000010000000100010011;
ROM[21523] <= 32'b00000011111100000000001110010011;
ROM[21524] <= 32'b00000000011100010010000000100011;
ROM[21525] <= 32'b00000000010000010000000100010011;
ROM[21526] <= 32'b00000011111100000000001110010011;
ROM[21527] <= 32'b00000000011100010010000000100011;
ROM[21528] <= 32'b00000000010000010000000100010011;
ROM[21529] <= 32'b00000011111100000000001110010011;
ROM[21530] <= 32'b00000000011100010010000000100011;
ROM[21531] <= 32'b00000000010000010000000100010011;
ROM[21532] <= 32'b00000011111100000000001110010011;
ROM[21533] <= 32'b00000000011100010010000000100011;
ROM[21534] <= 32'b00000000010000010000000100010011;
ROM[21535] <= 32'b00000000000000000000001110010011;
ROM[21536] <= 32'b00000000011100010010000000100011;
ROM[21537] <= 32'b00000000010000010000000100010011;
ROM[21538] <= 32'b00000000000000000000001110010011;
ROM[21539] <= 32'b00000000011100010010000000100011;
ROM[21540] <= 32'b00000000010000010000000100010011;
ROM[21541] <= 32'b00000000000000010101001110110111;
ROM[21542] <= 32'b00001110000000111000001110010011;
ROM[21543] <= 32'b00000000111000111000001110110011;
ROM[21544] <= 32'b00000000011100010010000000100011;
ROM[21545] <= 32'b00000000010000010000000100010011;
ROM[21546] <= 32'b00000000001100010010000000100011;
ROM[21547] <= 32'b00000000010000010000000100010011;
ROM[21548] <= 32'b00000000010000010010000000100011;
ROM[21549] <= 32'b00000000010000010000000100010011;
ROM[21550] <= 32'b00000000010100010010000000100011;
ROM[21551] <= 32'b00000000010000010000000100010011;
ROM[21552] <= 32'b00000000011000010010000000100011;
ROM[21553] <= 32'b00000000010000010000000100010011;
ROM[21554] <= 32'b00000001010000000000001110010011;
ROM[21555] <= 32'b00000010010000111000001110010011;
ROM[21556] <= 32'b01000000011100010000001110110011;
ROM[21557] <= 32'b00000000011100000000001000110011;
ROM[21558] <= 32'b00000000001000000000000110110011;
ROM[21559] <= 32'b01001110110000000000000011101111;
ROM[21560] <= 32'b11111111110000010000000100010011;
ROM[21561] <= 32'b00000000000000010010001110000011;
ROM[21562] <= 32'b00000000011101100010000000100011;
ROM[21563] <= 32'b00000100000100000000001110010011;
ROM[21564] <= 32'b00000000011100010010000000100011;
ROM[21565] <= 32'b00000000010000010000000100010011;
ROM[21566] <= 32'b00000000000000000000001110010011;
ROM[21567] <= 32'b00000000011100010010000000100011;
ROM[21568] <= 32'b00000000010000010000000100010011;
ROM[21569] <= 32'b00000000100000000000001110010011;
ROM[21570] <= 32'b00000000011100010010000000100011;
ROM[21571] <= 32'b00000000010000010000000100010011;
ROM[21572] <= 32'b00000001010000000000001110010011;
ROM[21573] <= 32'b00000000011100010010000000100011;
ROM[21574] <= 32'b00000000010000010000000100010011;
ROM[21575] <= 32'b00000010001000000000001110010011;
ROM[21576] <= 32'b00000000011100010010000000100011;
ROM[21577] <= 32'b00000000010000010000000100010011;
ROM[21578] <= 32'b00000011111000000000001110010011;
ROM[21579] <= 32'b00000000011100010010000000100011;
ROM[21580] <= 32'b00000000010000010000000100010011;
ROM[21581] <= 32'b00000010001000000000001110010011;
ROM[21582] <= 32'b00000000011100010010000000100011;
ROM[21583] <= 32'b00000000010000010000000100010011;
ROM[21584] <= 32'b00000010001000000000001110010011;
ROM[21585] <= 32'b00000000011100010010000000100011;
ROM[21586] <= 32'b00000000010000010000000100010011;
ROM[21587] <= 32'b00000000000000000000001110010011;
ROM[21588] <= 32'b00000000011100010010000000100011;
ROM[21589] <= 32'b00000000010000010000000100010011;
ROM[21590] <= 32'b00000000000000010101001110110111;
ROM[21591] <= 32'b00011010010000111000001110010011;
ROM[21592] <= 32'b00000000111000111000001110110011;
ROM[21593] <= 32'b00000000011100010010000000100011;
ROM[21594] <= 32'b00000000010000010000000100010011;
ROM[21595] <= 32'b00000000001100010010000000100011;
ROM[21596] <= 32'b00000000010000010000000100010011;
ROM[21597] <= 32'b00000000010000010010000000100011;
ROM[21598] <= 32'b00000000010000010000000100010011;
ROM[21599] <= 32'b00000000010100010010000000100011;
ROM[21600] <= 32'b00000000010000010000000100010011;
ROM[21601] <= 32'b00000000011000010010000000100011;
ROM[21602] <= 32'b00000000010000010000000100010011;
ROM[21603] <= 32'b00000001010000000000001110010011;
ROM[21604] <= 32'b00000010010000111000001110010011;
ROM[21605] <= 32'b01000000011100010000001110110011;
ROM[21606] <= 32'b00000000011100000000001000110011;
ROM[21607] <= 32'b00000000001000000000000110110011;
ROM[21608] <= 32'b01000010100000000000000011101111;
ROM[21609] <= 32'b11111111110000010000000100010011;
ROM[21610] <= 32'b00000000000000010010001110000011;
ROM[21611] <= 32'b00000000011101100010000000100011;
ROM[21612] <= 32'b00000100001000000000001110010011;
ROM[21613] <= 32'b00000000011100010010000000100011;
ROM[21614] <= 32'b00000000010000010000000100010011;
ROM[21615] <= 32'b00000001111000000000001110010011;
ROM[21616] <= 32'b00000000011100010010000000100011;
ROM[21617] <= 32'b00000000010000010000000100010011;
ROM[21618] <= 32'b00000010010000000000001110010011;
ROM[21619] <= 32'b00000000011100010010000000100011;
ROM[21620] <= 32'b00000000010000010000000100010011;
ROM[21621] <= 32'b00000010010000000000001110010011;
ROM[21622] <= 32'b00000000011100010010000000100011;
ROM[21623] <= 32'b00000000010000010000000100010011;
ROM[21624] <= 32'b00000011110000000000001110010011;
ROM[21625] <= 32'b00000000011100010010000000100011;
ROM[21626] <= 32'b00000000010000010000000100010011;
ROM[21627] <= 32'b00000010010000000000001110010011;
ROM[21628] <= 32'b00000000011100010010000000100011;
ROM[21629] <= 32'b00000000010000010000000100010011;
ROM[21630] <= 32'b00000010010000000000001110010011;
ROM[21631] <= 32'b00000000011100010010000000100011;
ROM[21632] <= 32'b00000000010000010000000100010011;
ROM[21633] <= 32'b00000001111000000000001110010011;
ROM[21634] <= 32'b00000000011100010010000000100011;
ROM[21635] <= 32'b00000000010000010000000100010011;
ROM[21636] <= 32'b00000000000000000000001110010011;
ROM[21637] <= 32'b00000000011100010010000000100011;
ROM[21638] <= 32'b00000000010000010000000100010011;
ROM[21639] <= 32'b00000000000000010101001110110111;
ROM[21640] <= 32'b00100110100000111000001110010011;
ROM[21641] <= 32'b00000000111000111000001110110011;
ROM[21642] <= 32'b00000000011100010010000000100011;
ROM[21643] <= 32'b00000000010000010000000100010011;
ROM[21644] <= 32'b00000000001100010010000000100011;
ROM[21645] <= 32'b00000000010000010000000100010011;
ROM[21646] <= 32'b00000000010000010010000000100011;
ROM[21647] <= 32'b00000000010000010000000100010011;
ROM[21648] <= 32'b00000000010100010010000000100011;
ROM[21649] <= 32'b00000000010000010000000100010011;
ROM[21650] <= 32'b00000000011000010010000000100011;
ROM[21651] <= 32'b00000000010000010000000100010011;
ROM[21652] <= 32'b00000001010000000000001110010011;
ROM[21653] <= 32'b00000010010000111000001110010011;
ROM[21654] <= 32'b01000000011100010000001110110011;
ROM[21655] <= 32'b00000000011100000000001000110011;
ROM[21656] <= 32'b00000000001000000000000110110011;
ROM[21657] <= 32'b00110110010000000000000011101111;
ROM[21658] <= 32'b11111111110000010000000100010011;
ROM[21659] <= 32'b00000000000000010010001110000011;
ROM[21660] <= 32'b00000000011101100010000000100011;
ROM[21661] <= 32'b00000100001100000000001110010011;
ROM[21662] <= 32'b00000000011100010010000000100011;
ROM[21663] <= 32'b00000000010000010000000100010011;
ROM[21664] <= 32'b00000000110000000000001110010011;
ROM[21665] <= 32'b00000000011100010010000000100011;
ROM[21666] <= 32'b00000000010000010000000100010011;
ROM[21667] <= 32'b00000001001000000000001110010011;
ROM[21668] <= 32'b00000000011100010010000000100011;
ROM[21669] <= 32'b00000000010000010000000100010011;
ROM[21670] <= 32'b00000010000000000000001110010011;
ROM[21671] <= 32'b00000000011100010010000000100011;
ROM[21672] <= 32'b00000000010000010000000100010011;
ROM[21673] <= 32'b00000010000000000000001110010011;
ROM[21674] <= 32'b00000000011100010010000000100011;
ROM[21675] <= 32'b00000000010000010000000100010011;
ROM[21676] <= 32'b00000010000000000000001110010011;
ROM[21677] <= 32'b00000000011100010010000000100011;
ROM[21678] <= 32'b00000000010000010000000100010011;
ROM[21679] <= 32'b00000001001000000000001110010011;
ROM[21680] <= 32'b00000000011100010010000000100011;
ROM[21681] <= 32'b00000000010000010000000100010011;
ROM[21682] <= 32'b00000000110000000000001110010011;
ROM[21683] <= 32'b00000000011100010010000000100011;
ROM[21684] <= 32'b00000000010000010000000100010011;
ROM[21685] <= 32'b00000000000000000000001110010011;
ROM[21686] <= 32'b00000000011100010010000000100011;
ROM[21687] <= 32'b00000000010000010000000100010011;
ROM[21688] <= 32'b00000000000000010101001110110111;
ROM[21689] <= 32'b00110010110000111000001110010011;
ROM[21690] <= 32'b00000000111000111000001110110011;
ROM[21691] <= 32'b00000000011100010010000000100011;
ROM[21692] <= 32'b00000000010000010000000100010011;
ROM[21693] <= 32'b00000000001100010010000000100011;
ROM[21694] <= 32'b00000000010000010000000100010011;
ROM[21695] <= 32'b00000000010000010010000000100011;
ROM[21696] <= 32'b00000000010000010000000100010011;
ROM[21697] <= 32'b00000000010100010010000000100011;
ROM[21698] <= 32'b00000000010000010000000100010011;
ROM[21699] <= 32'b00000000011000010010000000100011;
ROM[21700] <= 32'b00000000010000010000000100010011;
ROM[21701] <= 32'b00000001010000000000001110010011;
ROM[21702] <= 32'b00000010010000111000001110010011;
ROM[21703] <= 32'b01000000011100010000001110110011;
ROM[21704] <= 32'b00000000011100000000001000110011;
ROM[21705] <= 32'b00000000001000000000000110110011;
ROM[21706] <= 32'b00101010000000000000000011101111;
ROM[21707] <= 32'b11111111110000010000000100010011;
ROM[21708] <= 32'b00000000000000010010001110000011;
ROM[21709] <= 32'b00000000011101100010000000100011;
ROM[21710] <= 32'b00000100010000000000001110010011;
ROM[21711] <= 32'b00000000011100010010000000100011;
ROM[21712] <= 32'b00000000010000010000000100010011;
ROM[21713] <= 32'b00000001110000000000001110010011;
ROM[21714] <= 32'b00000000011100010010000000100011;
ROM[21715] <= 32'b00000000010000010000000100010011;
ROM[21716] <= 32'b00000010010000000000001110010011;
ROM[21717] <= 32'b00000000011100010010000000100011;
ROM[21718] <= 32'b00000000010000010000000100010011;
ROM[21719] <= 32'b00000010001000000000001110010011;
ROM[21720] <= 32'b00000000011100010010000000100011;
ROM[21721] <= 32'b00000000010000010000000100010011;
ROM[21722] <= 32'b00000010001000000000001110010011;
ROM[21723] <= 32'b00000000011100010010000000100011;
ROM[21724] <= 32'b00000000010000010000000100010011;
ROM[21725] <= 32'b00000010001000000000001110010011;
ROM[21726] <= 32'b00000000011100010010000000100011;
ROM[21727] <= 32'b00000000010000010000000100010011;
ROM[21728] <= 32'b00000010010000000000001110010011;
ROM[21729] <= 32'b00000000011100010010000000100011;
ROM[21730] <= 32'b00000000010000010000000100010011;
ROM[21731] <= 32'b00000001110000000000001110010011;
ROM[21732] <= 32'b00000000011100010010000000100011;
ROM[21733] <= 32'b00000000010000010000000100010011;
ROM[21734] <= 32'b00000000000000000000001110010011;
ROM[21735] <= 32'b00000000011100010010000000100011;
ROM[21736] <= 32'b00000000010000010000000100010011;
ROM[21737] <= 32'b00000000000000010101001110110111;
ROM[21738] <= 32'b00111111000000111000001110010011;
ROM[21739] <= 32'b00000000111000111000001110110011;
ROM[21740] <= 32'b00000000011100010010000000100011;
ROM[21741] <= 32'b00000000010000010000000100010011;
ROM[21742] <= 32'b00000000001100010010000000100011;
ROM[21743] <= 32'b00000000010000010000000100010011;
ROM[21744] <= 32'b00000000010000010010000000100011;
ROM[21745] <= 32'b00000000010000010000000100010011;
ROM[21746] <= 32'b00000000010100010010000000100011;
ROM[21747] <= 32'b00000000010000010000000100010011;
ROM[21748] <= 32'b00000000011000010010000000100011;
ROM[21749] <= 32'b00000000010000010000000100010011;
ROM[21750] <= 32'b00000001010000000000001110010011;
ROM[21751] <= 32'b00000010010000111000001110010011;
ROM[21752] <= 32'b01000000011100010000001110110011;
ROM[21753] <= 32'b00000000011100000000001000110011;
ROM[21754] <= 32'b00000000001000000000000110110011;
ROM[21755] <= 32'b00011101110000000000000011101111;
ROM[21756] <= 32'b11111111110000010000000100010011;
ROM[21757] <= 32'b00000000000000010010001110000011;
ROM[21758] <= 32'b00000000011101100010000000100011;
ROM[21759] <= 32'b00000100010100000000001110010011;
ROM[21760] <= 32'b00000000011100010010000000100011;
ROM[21761] <= 32'b00000000010000010000000100010011;
ROM[21762] <= 32'b00000011111000000000001110010011;
ROM[21763] <= 32'b00000000011100010010000000100011;
ROM[21764] <= 32'b00000000010000010000000100010011;
ROM[21765] <= 32'b00000010000000000000001110010011;
ROM[21766] <= 32'b00000000011100010010000000100011;
ROM[21767] <= 32'b00000000010000010000000100010011;
ROM[21768] <= 32'b00000010000000000000001110010011;
ROM[21769] <= 32'b00000000011100010010000000100011;
ROM[21770] <= 32'b00000000010000010000000100010011;
ROM[21771] <= 32'b00000011110000000000001110010011;
ROM[21772] <= 32'b00000000011100010010000000100011;
ROM[21773] <= 32'b00000000010000010000000100010011;
ROM[21774] <= 32'b00000010000000000000001110010011;
ROM[21775] <= 32'b00000000011100010010000000100011;
ROM[21776] <= 32'b00000000010000010000000100010011;
ROM[21777] <= 32'b00000010000000000000001110010011;
ROM[21778] <= 32'b00000000011100010010000000100011;
ROM[21779] <= 32'b00000000010000010000000100010011;
ROM[21780] <= 32'b00000011111000000000001110010011;
ROM[21781] <= 32'b00000000011100010010000000100011;
ROM[21782] <= 32'b00000000010000010000000100010011;
ROM[21783] <= 32'b00000000000000000000001110010011;
ROM[21784] <= 32'b00000000011100010010000000100011;
ROM[21785] <= 32'b00000000010000010000000100010011;
ROM[21786] <= 32'b00000000000000010101001110110111;
ROM[21787] <= 32'b01001011010000111000001110010011;
ROM[21788] <= 32'b00000000111000111000001110110011;
ROM[21789] <= 32'b00000000011100010010000000100011;
ROM[21790] <= 32'b00000000010000010000000100010011;
ROM[21791] <= 32'b00000000001100010010000000100011;
ROM[21792] <= 32'b00000000010000010000000100010011;
ROM[21793] <= 32'b00000000010000010010000000100011;
ROM[21794] <= 32'b00000000010000010000000100010011;
ROM[21795] <= 32'b00000000010100010010000000100011;
ROM[21796] <= 32'b00000000010000010000000100010011;
ROM[21797] <= 32'b00000000011000010010000000100011;
ROM[21798] <= 32'b00000000010000010000000100010011;
ROM[21799] <= 32'b00000001010000000000001110010011;
ROM[21800] <= 32'b00000010010000111000001110010011;
ROM[21801] <= 32'b01000000011100010000001110110011;
ROM[21802] <= 32'b00000000011100000000001000110011;
ROM[21803] <= 32'b00000000001000000000000110110011;
ROM[21804] <= 32'b00010001100000000000000011101111;
ROM[21805] <= 32'b11111111110000010000000100010011;
ROM[21806] <= 32'b00000000000000010010001110000011;
ROM[21807] <= 32'b00000000011101100010000000100011;
ROM[21808] <= 32'b00000100011000000000001110010011;
ROM[21809] <= 32'b00000000011100010010000000100011;
ROM[21810] <= 32'b00000000010000010000000100010011;
ROM[21811] <= 32'b00000011111000000000001110010011;
ROM[21812] <= 32'b00000000011100010010000000100011;
ROM[21813] <= 32'b00000000010000010000000100010011;
ROM[21814] <= 32'b00000010000000000000001110010011;
ROM[21815] <= 32'b00000000011100010010000000100011;
ROM[21816] <= 32'b00000000010000010000000100010011;
ROM[21817] <= 32'b00000010000000000000001110010011;
ROM[21818] <= 32'b00000000011100010010000000100011;
ROM[21819] <= 32'b00000000010000010000000100010011;
ROM[21820] <= 32'b00000011110000000000001110010011;
ROM[21821] <= 32'b00000000011100010010000000100011;
ROM[21822] <= 32'b00000000010000010000000100010011;
ROM[21823] <= 32'b00000010000000000000001110010011;
ROM[21824] <= 32'b00000000011100010010000000100011;
ROM[21825] <= 32'b00000000010000010000000100010011;
ROM[21826] <= 32'b00000010000000000000001110010011;
ROM[21827] <= 32'b00000000011100010010000000100011;
ROM[21828] <= 32'b00000000010000010000000100010011;
ROM[21829] <= 32'b00000010000000000000001110010011;
ROM[21830] <= 32'b00000000011100010010000000100011;
ROM[21831] <= 32'b00000000010000010000000100010011;
ROM[21832] <= 32'b00000000000000000000001110010011;
ROM[21833] <= 32'b00000000011100010010000000100011;
ROM[21834] <= 32'b00000000010000010000000100010011;
ROM[21835] <= 32'b00000000000000010101001110110111;
ROM[21836] <= 32'b01010111100000111000001110010011;
ROM[21837] <= 32'b00000000111000111000001110110011;
ROM[21838] <= 32'b00000000011100010010000000100011;
ROM[21839] <= 32'b00000000010000010000000100010011;
ROM[21840] <= 32'b00000000001100010010000000100011;
ROM[21841] <= 32'b00000000010000010000000100010011;
ROM[21842] <= 32'b00000000010000010010000000100011;
ROM[21843] <= 32'b00000000010000010000000100010011;
ROM[21844] <= 32'b00000000010100010010000000100011;
ROM[21845] <= 32'b00000000010000010000000100010011;
ROM[21846] <= 32'b00000000011000010010000000100011;
ROM[21847] <= 32'b00000000010000010000000100010011;
ROM[21848] <= 32'b00000001010000000000001110010011;
ROM[21849] <= 32'b00000010010000111000001110010011;
ROM[21850] <= 32'b01000000011100010000001110110011;
ROM[21851] <= 32'b00000000011100000000001000110011;
ROM[21852] <= 32'b00000000001000000000000110110011;
ROM[21853] <= 32'b00000101010000000000000011101111;
ROM[21854] <= 32'b11111111110000010000000100010011;
ROM[21855] <= 32'b00000000000000010010001110000011;
ROM[21856] <= 32'b00000000011101100010000000100011;
ROM[21857] <= 32'b00000000000000000000001110010011;
ROM[21858] <= 32'b00000000011100010010000000100011;
ROM[21859] <= 32'b00000000010000010000000100010011;
ROM[21860] <= 32'b00000001010000000000001110010011;
ROM[21861] <= 32'b01000000011100011000001110110011;
ROM[21862] <= 32'b00000000000000111010000010000011;
ROM[21863] <= 32'b11111111110000010000000100010011;
ROM[21864] <= 32'b00000000000000010010001110000011;
ROM[21865] <= 32'b00000000011100100010000000100011;
ROM[21866] <= 32'b00000000010000100000000100010011;
ROM[21867] <= 32'b00000001010000000000001110010011;
ROM[21868] <= 32'b01000000011100011000001110110011;
ROM[21869] <= 32'b00000000010000111010000110000011;
ROM[21870] <= 32'b00000000100000111010001000000011;
ROM[21871] <= 32'b00000000110000111010001010000011;
ROM[21872] <= 32'b00000001000000111010001100000011;
ROM[21873] <= 32'b00000000000000001000000011100111;
ROM[21874] <= 32'b00000000000000010010000000100011;
ROM[21875] <= 32'b00000000010000010000000100010011;
ROM[21876] <= 32'b00000000100000000000001110010011;
ROM[21877] <= 32'b00000000011100010010000000100011;
ROM[21878] <= 32'b00000000010000010000000100010011;
ROM[21879] <= 32'b00000000000000010101001110110111;
ROM[21880] <= 32'b01100010100000111000001110010011;
ROM[21881] <= 32'b00000000111000111000001110110011;
ROM[21882] <= 32'b00000000011100010010000000100011;
ROM[21883] <= 32'b00000000010000010000000100010011;
ROM[21884] <= 32'b00000000001100010010000000100011;
ROM[21885] <= 32'b00000000010000010000000100010011;
ROM[21886] <= 32'b00000000010000010010000000100011;
ROM[21887] <= 32'b00000000010000010000000100010011;
ROM[21888] <= 32'b00000000010100010010000000100011;
ROM[21889] <= 32'b00000000010000010000000100010011;
ROM[21890] <= 32'b00000000011000010010000000100011;
ROM[21891] <= 32'b00000000010000010000000100010011;
ROM[21892] <= 32'b00000001010000000000001110010011;
ROM[21893] <= 32'b00000000010000111000001110010011;
ROM[21894] <= 32'b01000000011100010000001110110011;
ROM[21895] <= 32'b00000000011100000000001000110011;
ROM[21896] <= 32'b00000000001000000000000110110011;
ROM[21897] <= 32'b10100101110111101010000011101111;
ROM[21898] <= 32'b11111111110000010000000100010011;
ROM[21899] <= 32'b00000000000000010010001110000011;
ROM[21900] <= 32'b00000000011100011010000000100011;
ROM[21901] <= 32'b00000000000000100010001110000011;
ROM[21902] <= 32'b00000000011100010010000000100011;
ROM[21903] <= 32'b00000000010000010000000100010011;
ROM[21904] <= 32'b00000000010000000000001110010011;
ROM[21905] <= 32'b00000000011100010010000000100011;
ROM[21906] <= 32'b00000000010000010000000100010011;
ROM[21907] <= 32'b00000000000000010101001110110111;
ROM[21908] <= 32'b01101001100000111000001110010011;
ROM[21909] <= 32'b00000000111000111000001110110011;
ROM[21910] <= 32'b00000000011100010010000000100011;
ROM[21911] <= 32'b00000000010000010000000100010011;
ROM[21912] <= 32'b00000000001100010010000000100011;
ROM[21913] <= 32'b00000000010000010000000100010011;
ROM[21914] <= 32'b00000000010000010010000000100011;
ROM[21915] <= 32'b00000000010000010000000100010011;
ROM[21916] <= 32'b00000000010100010010000000100011;
ROM[21917] <= 32'b00000000010000010000000100010011;
ROM[21918] <= 32'b00000000011000010010000000100011;
ROM[21919] <= 32'b00000000010000010000000100010011;
ROM[21920] <= 32'b00000001010000000000001110010011;
ROM[21921] <= 32'b00000000100000111000001110010011;
ROM[21922] <= 32'b01000000011100010000001110110011;
ROM[21923] <= 32'b00000000011100000000001000110011;
ROM[21924] <= 32'b00000000001000000000000110110011;
ROM[21925] <= 32'b10011001100011111100000011101111;
ROM[21926] <= 32'b11111111110000010000000100010011;
ROM[21927] <= 32'b00000000000000010010001110000011;
ROM[21928] <= 32'b00000000011100100010000000100011;
ROM[21929] <= 32'b00000000000000011010001110000011;
ROM[21930] <= 32'b00000000011100010010000000100011;
ROM[21931] <= 32'b00000000010000010000000100010011;
ROM[21932] <= 32'b00001000100001101010001110000011;
ROM[21933] <= 32'b00000000011100010010000000100011;
ROM[21934] <= 32'b00000000010000010000000100010011;
ROM[21935] <= 32'b00000000000000100010001110000011;
ROM[21936] <= 32'b00000000011100010010000000100011;
ROM[21937] <= 32'b00000000010000010000000100010011;
ROM[21938] <= 32'b11111111110000010000000100010011;
ROM[21939] <= 32'b00000000000000010010001110000011;
ROM[21940] <= 32'b11111111110000010000000100010011;
ROM[21941] <= 32'b00000000000000010010010000000011;
ROM[21942] <= 32'b00000000011101000000001110110011;
ROM[21943] <= 32'b00000000011100010010000000100011;
ROM[21944] <= 32'b00000000010000010000000100010011;
ROM[21945] <= 32'b11111111110000010000000100010011;
ROM[21946] <= 32'b00000000000000010010001110000011;
ROM[21947] <= 32'b00000000000000111000001100010011;
ROM[21948] <= 32'b11111111110000010000000100010011;
ROM[21949] <= 32'b00000000000000010010001110000011;
ROM[21950] <= 32'b00000000110100110000010000110011;
ROM[21951] <= 32'b00000000011101000010000000100011;
ROM[21952] <= 32'b00000000010000100010001110000011;
ROM[21953] <= 32'b00000000011100010010000000100011;
ROM[21954] <= 32'b00000000010000010000000100010011;
ROM[21955] <= 32'b00000000000000011010001110000011;
ROM[21956] <= 32'b00000000011100010010000000100011;
ROM[21957] <= 32'b00000000010000010000000100010011;
ROM[21958] <= 32'b00000000000000000000001110010011;
ROM[21959] <= 32'b00000000011100010010000000100011;
ROM[21960] <= 32'b00000000010000010000000100010011;
ROM[21961] <= 32'b11111111110000010000000100010011;
ROM[21962] <= 32'b00000000000000010010001110000011;
ROM[21963] <= 32'b11111111110000010000000100010011;
ROM[21964] <= 32'b00000000000000010010010000000011;
ROM[21965] <= 32'b00000000011101000000001110110011;
ROM[21966] <= 32'b00000000011100010010000000100011;
ROM[21967] <= 32'b00000000010000010000000100010011;
ROM[21968] <= 32'b11111111110000010000000100010011;
ROM[21969] <= 32'b00000000000000010010001110000011;
ROM[21970] <= 32'b00000000000000111000001100010011;
ROM[21971] <= 32'b11111111110000010000000100010011;
ROM[21972] <= 32'b00000000000000010010001110000011;
ROM[21973] <= 32'b00000000110100110000010000110011;
ROM[21974] <= 32'b00000000011101000010000000100011;
ROM[21975] <= 32'b00000000100000100010001110000011;
ROM[21976] <= 32'b00000000011100010010000000100011;
ROM[21977] <= 32'b00000000010000010000000100010011;
ROM[21978] <= 32'b00000000000000011010001110000011;
ROM[21979] <= 32'b00000000011100010010000000100011;
ROM[21980] <= 32'b00000000010000010000000100010011;
ROM[21981] <= 32'b00000000010000000000001110010011;
ROM[21982] <= 32'b00000000011100010010000000100011;
ROM[21983] <= 32'b00000000010000010000000100010011;
ROM[21984] <= 32'b11111111110000010000000100010011;
ROM[21985] <= 32'b00000000000000010010001110000011;
ROM[21986] <= 32'b11111111110000010000000100010011;
ROM[21987] <= 32'b00000000000000010010010000000011;
ROM[21988] <= 32'b00000000011101000000001110110011;
ROM[21989] <= 32'b00000000011100010010000000100011;
ROM[21990] <= 32'b00000000010000010000000100010011;
ROM[21991] <= 32'b11111111110000010000000100010011;
ROM[21992] <= 32'b00000000000000010010001110000011;
ROM[21993] <= 32'b00000000000000111000001100010011;
ROM[21994] <= 32'b11111111110000010000000100010011;
ROM[21995] <= 32'b00000000000000010010001110000011;
ROM[21996] <= 32'b00000000110100110000010000110011;
ROM[21997] <= 32'b00000000011101000010000000100011;
ROM[21998] <= 32'b00000000110000100010001110000011;
ROM[21999] <= 32'b00000000011100010010000000100011;
ROM[22000] <= 32'b00000000010000010000000100010011;
ROM[22001] <= 32'b00000000000000011010001110000011;
ROM[22002] <= 32'b00000000011100010010000000100011;
ROM[22003] <= 32'b00000000010000010000000100010011;
ROM[22004] <= 32'b00000000100000000000001110010011;
ROM[22005] <= 32'b00000000011100010010000000100011;
ROM[22006] <= 32'b00000000010000010000000100010011;
ROM[22007] <= 32'b11111111110000010000000100010011;
ROM[22008] <= 32'b00000000000000010010001110000011;
ROM[22009] <= 32'b11111111110000010000000100010011;
ROM[22010] <= 32'b00000000000000010010010000000011;
ROM[22011] <= 32'b00000000011101000000001110110011;
ROM[22012] <= 32'b00000000011100010010000000100011;
ROM[22013] <= 32'b00000000010000010000000100010011;
ROM[22014] <= 32'b11111111110000010000000100010011;
ROM[22015] <= 32'b00000000000000010010001110000011;
ROM[22016] <= 32'b00000000000000111000001100010011;
ROM[22017] <= 32'b11111111110000010000000100010011;
ROM[22018] <= 32'b00000000000000010010001110000011;
ROM[22019] <= 32'b00000000110100110000010000110011;
ROM[22020] <= 32'b00000000011101000010000000100011;
ROM[22021] <= 32'b00000001000000100010001110000011;
ROM[22022] <= 32'b00000000011100010010000000100011;
ROM[22023] <= 32'b00000000010000010000000100010011;
ROM[22024] <= 32'b00000000000000011010001110000011;
ROM[22025] <= 32'b00000000011100010010000000100011;
ROM[22026] <= 32'b00000000010000010000000100010011;
ROM[22027] <= 32'b00000000110000000000001110010011;
ROM[22028] <= 32'b00000000011100010010000000100011;
ROM[22029] <= 32'b00000000010000010000000100010011;
ROM[22030] <= 32'b11111111110000010000000100010011;
ROM[22031] <= 32'b00000000000000010010001110000011;
ROM[22032] <= 32'b11111111110000010000000100010011;
ROM[22033] <= 32'b00000000000000010010010000000011;
ROM[22034] <= 32'b00000000011101000000001110110011;
ROM[22035] <= 32'b00000000011100010010000000100011;
ROM[22036] <= 32'b00000000010000010000000100010011;
ROM[22037] <= 32'b11111111110000010000000100010011;
ROM[22038] <= 32'b00000000000000010010001110000011;
ROM[22039] <= 32'b00000000000000111000001100010011;
ROM[22040] <= 32'b11111111110000010000000100010011;
ROM[22041] <= 32'b00000000000000010010001110000011;
ROM[22042] <= 32'b00000000110100110000010000110011;
ROM[22043] <= 32'b00000000011101000010000000100011;
ROM[22044] <= 32'b00000001010000100010001110000011;
ROM[22045] <= 32'b00000000011100010010000000100011;
ROM[22046] <= 32'b00000000010000010000000100010011;
ROM[22047] <= 32'b00000000000000011010001110000011;
ROM[22048] <= 32'b00000000011100010010000000100011;
ROM[22049] <= 32'b00000000010000010000000100010011;
ROM[22050] <= 32'b00000001000000000000001110010011;
ROM[22051] <= 32'b00000000011100010010000000100011;
ROM[22052] <= 32'b00000000010000010000000100010011;
ROM[22053] <= 32'b11111111110000010000000100010011;
ROM[22054] <= 32'b00000000000000010010001110000011;
ROM[22055] <= 32'b11111111110000010000000100010011;
ROM[22056] <= 32'b00000000000000010010010000000011;
ROM[22057] <= 32'b00000000011101000000001110110011;
ROM[22058] <= 32'b00000000011100010010000000100011;
ROM[22059] <= 32'b00000000010000010000000100010011;
ROM[22060] <= 32'b11111111110000010000000100010011;
ROM[22061] <= 32'b00000000000000010010001110000011;
ROM[22062] <= 32'b00000000000000111000001100010011;
ROM[22063] <= 32'b11111111110000010000000100010011;
ROM[22064] <= 32'b00000000000000010010001110000011;
ROM[22065] <= 32'b00000000110100110000010000110011;
ROM[22066] <= 32'b00000000011101000010000000100011;
ROM[22067] <= 32'b00000001100000100010001110000011;
ROM[22068] <= 32'b00000000011100010010000000100011;
ROM[22069] <= 32'b00000000010000010000000100010011;
ROM[22070] <= 32'b00000000000000011010001110000011;
ROM[22071] <= 32'b00000000011100010010000000100011;
ROM[22072] <= 32'b00000000010000010000000100010011;
ROM[22073] <= 32'b00000001010000000000001110010011;
ROM[22074] <= 32'b00000000011100010010000000100011;
ROM[22075] <= 32'b00000000010000010000000100010011;
ROM[22076] <= 32'b11111111110000010000000100010011;
ROM[22077] <= 32'b00000000000000010010001110000011;
ROM[22078] <= 32'b11111111110000010000000100010011;
ROM[22079] <= 32'b00000000000000010010010000000011;
ROM[22080] <= 32'b00000000011101000000001110110011;
ROM[22081] <= 32'b00000000011100010010000000100011;
ROM[22082] <= 32'b00000000010000010000000100010011;
ROM[22083] <= 32'b11111111110000010000000100010011;
ROM[22084] <= 32'b00000000000000010010001110000011;
ROM[22085] <= 32'b00000000000000111000001100010011;
ROM[22086] <= 32'b11111111110000010000000100010011;
ROM[22087] <= 32'b00000000000000010010001110000011;
ROM[22088] <= 32'b00000000110100110000010000110011;
ROM[22089] <= 32'b00000000011101000010000000100011;
ROM[22090] <= 32'b00000001110000100010001110000011;
ROM[22091] <= 32'b00000000011100010010000000100011;
ROM[22092] <= 32'b00000000010000010000000100010011;
ROM[22093] <= 32'b00000000000000011010001110000011;
ROM[22094] <= 32'b00000000011100010010000000100011;
ROM[22095] <= 32'b00000000010000010000000100010011;
ROM[22096] <= 32'b00000001100000000000001110010011;
ROM[22097] <= 32'b00000000011100010010000000100011;
ROM[22098] <= 32'b00000000010000010000000100010011;
ROM[22099] <= 32'b11111111110000010000000100010011;
ROM[22100] <= 32'b00000000000000010010001110000011;
ROM[22101] <= 32'b11111111110000010000000100010011;
ROM[22102] <= 32'b00000000000000010010010000000011;
ROM[22103] <= 32'b00000000011101000000001110110011;
ROM[22104] <= 32'b00000000011100010010000000100011;
ROM[22105] <= 32'b00000000010000010000000100010011;
ROM[22106] <= 32'b11111111110000010000000100010011;
ROM[22107] <= 32'b00000000000000010010001110000011;
ROM[22108] <= 32'b00000000000000111000001100010011;
ROM[22109] <= 32'b11111111110000010000000100010011;
ROM[22110] <= 32'b00000000000000010010001110000011;
ROM[22111] <= 32'b00000000110100110000010000110011;
ROM[22112] <= 32'b00000000011101000010000000100011;
ROM[22113] <= 32'b00000010000000100010001110000011;
ROM[22114] <= 32'b00000000011100010010000000100011;
ROM[22115] <= 32'b00000000010000010000000100010011;
ROM[22116] <= 32'b00000000000000011010001110000011;
ROM[22117] <= 32'b00000000011100010010000000100011;
ROM[22118] <= 32'b00000000010000010000000100010011;
ROM[22119] <= 32'b00000001110000000000001110010011;
ROM[22120] <= 32'b00000000011100010010000000100011;
ROM[22121] <= 32'b00000000010000010000000100010011;
ROM[22122] <= 32'b11111111110000010000000100010011;
ROM[22123] <= 32'b00000000000000010010001110000011;
ROM[22124] <= 32'b11111111110000010000000100010011;
ROM[22125] <= 32'b00000000000000010010010000000011;
ROM[22126] <= 32'b00000000011101000000001110110011;
ROM[22127] <= 32'b00000000011100010010000000100011;
ROM[22128] <= 32'b00000000010000010000000100010011;
ROM[22129] <= 32'b11111111110000010000000100010011;
ROM[22130] <= 32'b00000000000000010010001110000011;
ROM[22131] <= 32'b00000000000000111000001100010011;
ROM[22132] <= 32'b11111111110000010000000100010011;
ROM[22133] <= 32'b00000000000000010010001110000011;
ROM[22134] <= 32'b00000000110100110000010000110011;
ROM[22135] <= 32'b00000000011101000010000000100011;
ROM[22136] <= 32'b00000000000000000000001110010011;
ROM[22137] <= 32'b00000000011100010010000000100011;
ROM[22138] <= 32'b00000000010000010000000100010011;
ROM[22139] <= 32'b00000001010000000000001110010011;
ROM[22140] <= 32'b01000000011100011000001110110011;
ROM[22141] <= 32'b00000000000000111010000010000011;
ROM[22142] <= 32'b11111111110000010000000100010011;
ROM[22143] <= 32'b00000000000000010010001110000011;
ROM[22144] <= 32'b00000000011100100010000000100011;
ROM[22145] <= 32'b00000000010000100000000100010011;
ROM[22146] <= 32'b00000001010000000000001110010011;
ROM[22147] <= 32'b01000000011100011000001110110011;
ROM[22148] <= 32'b00000000010000111010000110000011;
ROM[22149] <= 32'b00000000100000111010001000000011;
ROM[22150] <= 32'b00000000110000111010001010000011;
ROM[22151] <= 32'b00000001000000111010001100000011;
ROM[22152] <= 32'b00000000000000001000000011100111;
ROM[22153] <= 32'b00000000000000010010000000100011;
ROM[22154] <= 32'b00000000010000010000000100010011;
ROM[22155] <= 32'b00000000000000100010001110000011;
ROM[22156] <= 32'b00000000011100010010000000100011;
ROM[22157] <= 32'b00000000010000010000000100010011;
ROM[22158] <= 32'b00000010000000000000001110010011;
ROM[22159] <= 32'b00000000011100010010000000100011;
ROM[22160] <= 32'b00000000010000010000000100010011;
ROM[22161] <= 32'b11111111110000010000000100010011;
ROM[22162] <= 32'b00000000000000010010001110000011;
ROM[22163] <= 32'b11111111110000010000000100010011;
ROM[22164] <= 32'b00000000000000010010010000000011;
ROM[22165] <= 32'b00000000011101000010001110110011;
ROM[22166] <= 32'b00000000011100010010000000100011;
ROM[22167] <= 32'b00000000010000010000000100010011;
ROM[22168] <= 32'b00000000000000100010001110000011;
ROM[22169] <= 32'b00000000011100010010000000100011;
ROM[22170] <= 32'b00000000010000010000000100010011;
ROM[22171] <= 32'b00000111111000000000001110010011;
ROM[22172] <= 32'b00000000011100010010000000100011;
ROM[22173] <= 32'b00000000010000010000000100010011;
ROM[22174] <= 32'b11111111110000010000000100010011;
ROM[22175] <= 32'b00000000000000010010001110000011;
ROM[22176] <= 32'b11111111110000010000000100010011;
ROM[22177] <= 32'b00000000000000010010010000000011;
ROM[22178] <= 32'b00000000100000111010001110110011;
ROM[22179] <= 32'b00000000011100010010000000100011;
ROM[22180] <= 32'b00000000010000010000000100010011;
ROM[22181] <= 32'b11111111110000010000000100010011;
ROM[22182] <= 32'b00000000000000010010001110000011;
ROM[22183] <= 32'b11111111110000010000000100010011;
ROM[22184] <= 32'b00000000000000010010010000000011;
ROM[22185] <= 32'b00000000011101000110001110110011;
ROM[22186] <= 32'b00000000011100010010000000100011;
ROM[22187] <= 32'b00000000010000010000000100010011;
ROM[22188] <= 32'b11111111110000010000000100010011;
ROM[22189] <= 32'b00000000000000010010001110000011;
ROM[22190] <= 32'b00000000000000111000101001100011;
ROM[22191] <= 32'b00000000000000010110001110110111;
ROM[22192] <= 32'b10101101000000111000001110010011;
ROM[22193] <= 32'b00000000111000111000001110110011;
ROM[22194] <= 32'b00000000000000111000000011100111;
ROM[22195] <= 32'b00000001110000000000000011101111;
ROM[22196] <= 32'b00000000000000000000001110010011;
ROM[22197] <= 32'b00000000011100010010000000100011;
ROM[22198] <= 32'b00000000010000010000000100010011;
ROM[22199] <= 32'b11111111110000010000000100010011;
ROM[22200] <= 32'b00000000000000010010001110000011;
ROM[22201] <= 32'b00000000011100100010000000100011;
ROM[22202] <= 32'b00000000000000100010001110000011;
ROM[22203] <= 32'b00000000011100010010000000100011;
ROM[22204] <= 32'b00000000010000010000000100010011;
ROM[22205] <= 32'b00000000000000100010001110000011;
ROM[22206] <= 32'b00000000011100010010000000100011;
ROM[22207] <= 32'b00000000010000010000000100010011;
ROM[22208] <= 32'b11111111110000010000000100010011;
ROM[22209] <= 32'b00000000000000010010001110000011;
ROM[22210] <= 32'b11111111110000010000000100010011;
ROM[22211] <= 32'b00000000000000010010010000000011;
ROM[22212] <= 32'b00000000011101000000001110110011;
ROM[22213] <= 32'b00000000011100010010000000100011;
ROM[22214] <= 32'b00000000010000010000000100010011;
ROM[22215] <= 32'b00000000000000100010001110000011;
ROM[22216] <= 32'b00000000011100010010000000100011;
ROM[22217] <= 32'b00000000010000010000000100010011;
ROM[22218] <= 32'b11111111110000010000000100010011;
ROM[22219] <= 32'b00000000000000010010001110000011;
ROM[22220] <= 32'b11111111110000010000000100010011;
ROM[22221] <= 32'b00000000000000010010010000000011;
ROM[22222] <= 32'b00000000011101000000001110110011;
ROM[22223] <= 32'b00000000011100010010000000100011;
ROM[22224] <= 32'b00000000010000010000000100010011;
ROM[22225] <= 32'b00000000000000100010001110000011;
ROM[22226] <= 32'b00000000011100010010000000100011;
ROM[22227] <= 32'b00000000010000010000000100010011;
ROM[22228] <= 32'b11111111110000010000000100010011;
ROM[22229] <= 32'b00000000000000010010001110000011;
ROM[22230] <= 32'b11111111110000010000000100010011;
ROM[22231] <= 32'b00000000000000010010010000000011;
ROM[22232] <= 32'b00000000011101000000001110110011;
ROM[22233] <= 32'b00000000011100010010000000100011;
ROM[22234] <= 32'b00000000010000010000000100010011;
ROM[22235] <= 32'b11111111110000010000000100010011;
ROM[22236] <= 32'b00000000000000010010001110000011;
ROM[22237] <= 32'b00000000011100011010000000100011;
ROM[22238] <= 32'b00001000100001101010001110000011;
ROM[22239] <= 32'b00000000011100010010000000100011;
ROM[22240] <= 32'b00000000010000010000000100010011;
ROM[22241] <= 32'b00000000000000011010001110000011;
ROM[22242] <= 32'b00000000011100010010000000100011;
ROM[22243] <= 32'b00000000010000010000000100010011;
ROM[22244] <= 32'b11111111110000010000000100010011;
ROM[22245] <= 32'b00000000000000010010001110000011;
ROM[22246] <= 32'b11111111110000010000000100010011;
ROM[22247] <= 32'b00000000000000010010010000000011;
ROM[22248] <= 32'b00000000011101000000001110110011;
ROM[22249] <= 32'b00000000011100010010000000100011;
ROM[22250] <= 32'b00000000010000010000000100010011;
ROM[22251] <= 32'b11111111110000010000000100010011;
ROM[22252] <= 32'b00000000000000010010001110000011;
ROM[22253] <= 32'b00000000000000111000001100010011;
ROM[22254] <= 32'b00000000110100110000010000110011;
ROM[22255] <= 32'b00000000000001000010001110000011;
ROM[22256] <= 32'b00000000011100010010000000100011;
ROM[22257] <= 32'b00000000010000010000000100010011;
ROM[22258] <= 32'b00000001010000000000001110010011;
ROM[22259] <= 32'b01000000011100011000001110110011;
ROM[22260] <= 32'b00000000000000111010000010000011;
ROM[22261] <= 32'b11111111110000010000000100010011;
ROM[22262] <= 32'b00000000000000010010001110000011;
ROM[22263] <= 32'b00000000011100100010000000100011;
ROM[22264] <= 32'b00000000010000100000000100010011;
ROM[22265] <= 32'b00000001010000000000001110010011;
ROM[22266] <= 32'b01000000011100011000001110110011;
ROM[22267] <= 32'b00000000010000111010000110000011;
ROM[22268] <= 32'b00000000100000111010001000000011;
ROM[22269] <= 32'b00000000110000111010001010000011;
ROM[22270] <= 32'b00000001000000111010001100000011;
ROM[22271] <= 32'b00000000000000001000000011100111;
ROM[22272] <= 32'b00000000010000100010001110000011;
ROM[22273] <= 32'b00000000011100010010000000100011;
ROM[22274] <= 32'b00000000010000010000000100010011;
ROM[22275] <= 32'b11111111110000010000000100010011;
ROM[22276] <= 32'b00000000000000010010001110000011;
ROM[22277] <= 32'b00001000011101101010000000100011;
ROM[22278] <= 32'b00000000000000100010001110000011;
ROM[22279] <= 32'b00000000011100010010000000100011;
ROM[22280] <= 32'b00000000010000010000000100010011;
ROM[22281] <= 32'b11111111110000010000000100010011;
ROM[22282] <= 32'b00000000000000010010001110000011;
ROM[22283] <= 32'b00001000011101101010001000100011;
ROM[22284] <= 32'b00000000000000000000001110010011;
ROM[22285] <= 32'b00000000011100010010000000100011;
ROM[22286] <= 32'b00000000010000010000000100010011;
ROM[22287] <= 32'b00000001010000000000001110010011;
ROM[22288] <= 32'b01000000011100011000001110110011;
ROM[22289] <= 32'b00000000000000111010000010000011;
ROM[22290] <= 32'b11111111110000010000000100010011;
ROM[22291] <= 32'b00000000000000010010001110000011;
ROM[22292] <= 32'b00000000011100100010000000100011;
ROM[22293] <= 32'b00000000010000100000000100010011;
ROM[22294] <= 32'b00000001010000000000001110010011;
ROM[22295] <= 32'b01000000011100011000001110110011;
ROM[22296] <= 32'b00000000010000111010000110000011;
ROM[22297] <= 32'b00000000100000111010001000000011;
ROM[22298] <= 32'b00000000110000111010001010000011;
ROM[22299] <= 32'b00000001000000111010001100000011;
ROM[22300] <= 32'b00000000000000001000000011100111;
ROM[22301] <= 32'b00000000000000010010000000100011;
ROM[22302] <= 32'b00000000010000010000000100010011;
ROM[22303] <= 32'b00000000000000010010000000100011;
ROM[22304] <= 32'b00000000010000010000000100010011;
ROM[22305] <= 32'b00000000000000010010000000100011;
ROM[22306] <= 32'b00000000010000010000000100010011;
ROM[22307] <= 32'b00000000000000010010000000100011;
ROM[22308] <= 32'b00000000010000010000000100010011;
ROM[22309] <= 32'b00000000000000010010000000100011;
ROM[22310] <= 32'b00000000010000010000000100010011;
ROM[22311] <= 32'b00000000000000010010000000100011;
ROM[22312] <= 32'b00000000010000010000000100010011;
ROM[22313] <= 32'b00000000000000010010000000100011;
ROM[22314] <= 32'b00000000010000010000000100010011;
ROM[22315] <= 32'b00000000000000010010000000100011;
ROM[22316] <= 32'b00000000010000010000000100010011;
ROM[22317] <= 32'b00000000000000010010000000100011;
ROM[22318] <= 32'b00000000010000010000000100010011;
ROM[22319] <= 32'b00000000000000010010000000100011;
ROM[22320] <= 32'b00000000010000010000000100010011;
ROM[22321] <= 32'b00000000000000010010000000100011;
ROM[22322] <= 32'b00000000010000010000000100010011;
ROM[22323] <= 32'b00000000000000100010001110000011;
ROM[22324] <= 32'b00000000011100010010000000100011;
ROM[22325] <= 32'b00000000010000010000000100010011;
ROM[22326] <= 32'b00000000000000010110001110110111;
ROM[22327] <= 32'b11010010010000111000001110010011;
ROM[22328] <= 32'b00000000111000111000001110110011;
ROM[22329] <= 32'b00000000011100010010000000100011;
ROM[22330] <= 32'b00000000010000010000000100010011;
ROM[22331] <= 32'b00000000001100010010000000100011;
ROM[22332] <= 32'b00000000010000010000000100010011;
ROM[22333] <= 32'b00000000010000010010000000100011;
ROM[22334] <= 32'b00000000010000010000000100010011;
ROM[22335] <= 32'b00000000010100010010000000100011;
ROM[22336] <= 32'b00000000010000010000000100010011;
ROM[22337] <= 32'b00000000011000010010000000100011;
ROM[22338] <= 32'b00000000010000010000000100010011;
ROM[22339] <= 32'b00000001010000000000001110010011;
ROM[22340] <= 32'b00000000010000111000001110010011;
ROM[22341] <= 32'b01000000011100010000001110110011;
ROM[22342] <= 32'b00000000011100000000001000110011;
ROM[22343] <= 32'b00000000001000000000000110110011;
ROM[22344] <= 32'b11010000010111111111000011101111;
ROM[22345] <= 32'b11111111110000010000000100010011;
ROM[22346] <= 32'b00000000000000010010001110000011;
ROM[22347] <= 32'b00000000011100011010000000100011;
ROM[22348] <= 32'b00001000010001101010001110000011;
ROM[22349] <= 32'b00000000011100010010000000100011;
ROM[22350] <= 32'b00000000010000010000000100010011;
ROM[22351] <= 32'b00000000101000000000001110010011;
ROM[22352] <= 32'b00000000011100010010000000100011;
ROM[22353] <= 32'b00000000010000010000000100010011;
ROM[22354] <= 32'b00000000000000010110001110110111;
ROM[22355] <= 32'b11011001010000111000001110010011;
ROM[22356] <= 32'b00000000111000111000001110110011;
ROM[22357] <= 32'b00000000011100010010000000100011;
ROM[22358] <= 32'b00000000010000010000000100010011;
ROM[22359] <= 32'b00000000001100010010000000100011;
ROM[22360] <= 32'b00000000010000010000000100010011;
ROM[22361] <= 32'b00000000010000010010000000100011;
ROM[22362] <= 32'b00000000010000010000000100010011;
ROM[22363] <= 32'b00000000010100010010000000100011;
ROM[22364] <= 32'b00000000010000010000000100010011;
ROM[22365] <= 32'b00000000011000010010000000100011;
ROM[22366] <= 32'b00000000010000010000000100010011;
ROM[22367] <= 32'b00000001010000000000001110010011;
ROM[22368] <= 32'b00000000100000111000001110010011;
ROM[22369] <= 32'b01000000011100010000001110110011;
ROM[22370] <= 32'b00000000011100000000001000110011;
ROM[22371] <= 32'b00000000001000000000000110110011;
ROM[22372] <= 32'b10101001110111111011000011101111;
ROM[22373] <= 32'b00000000100000000000001110010011;
ROM[22374] <= 32'b00000000011100010010000000100011;
ROM[22375] <= 32'b00000000010000010000000100010011;
ROM[22376] <= 32'b00000000000000010110001110110111;
ROM[22377] <= 32'b11011110110000111000001110010011;
ROM[22378] <= 32'b00000000111000111000001110110011;
ROM[22379] <= 32'b00000000011100010010000000100011;
ROM[22380] <= 32'b00000000010000010000000100010011;
ROM[22381] <= 32'b00000000001100010010000000100011;
ROM[22382] <= 32'b00000000010000010000000100010011;
ROM[22383] <= 32'b00000000010000010010000000100011;
ROM[22384] <= 32'b00000000010000010000000100010011;
ROM[22385] <= 32'b00000000010100010010000000100011;
ROM[22386] <= 32'b00000000010000010000000100010011;
ROM[22387] <= 32'b00000000011000010010000000100011;
ROM[22388] <= 32'b00000000010000010000000100010011;
ROM[22389] <= 32'b00000001010000000000001110010011;
ROM[22390] <= 32'b00000000100000111000001110010011;
ROM[22391] <= 32'b01000000011100010000001110110011;
ROM[22392] <= 32'b00000000011100000000001000110011;
ROM[22393] <= 32'b00000000001000000000000110110011;
ROM[22394] <= 32'b10100100010111111011000011101111;
ROM[22395] <= 32'b00001000000001101010001110000011;
ROM[22396] <= 32'b00000000011100010010000000100011;
ROM[22397] <= 32'b00000000010000010000000100010011;
ROM[22398] <= 32'b00000000010000000000001110010011;
ROM[22399] <= 32'b00000000011100010010000000100011;
ROM[22400] <= 32'b00000000010000010000000100010011;
ROM[22401] <= 32'b00000000000000010110001110110111;
ROM[22402] <= 32'b11100101000000111000001110010011;
ROM[22403] <= 32'b00000000111000111000001110110011;
ROM[22404] <= 32'b00000000011100010010000000100011;
ROM[22405] <= 32'b00000000010000010000000100010011;
ROM[22406] <= 32'b00000000001100010010000000100011;
ROM[22407] <= 32'b00000000010000010000000100010011;
ROM[22408] <= 32'b00000000010000010010000000100011;
ROM[22409] <= 32'b00000000010000010000000100010011;
ROM[22410] <= 32'b00000000010100010010000000100011;
ROM[22411] <= 32'b00000000010000010000000100010011;
ROM[22412] <= 32'b00000000011000010010000000100011;
ROM[22413] <= 32'b00000000010000010000000100010011;
ROM[22414] <= 32'b00000001010000000000001110010011;
ROM[22415] <= 32'b00000000100000111000001110010011;
ROM[22416] <= 32'b01000000011100010000001110110011;
ROM[22417] <= 32'b00000000011100000000001000110011;
ROM[22418] <= 32'b00000000001000000000000110110011;
ROM[22419] <= 32'b11010101110111111011000011101111;
ROM[22420] <= 32'b11111111110000010000000100010011;
ROM[22421] <= 32'b00000000000000010010001110000011;
ROM[22422] <= 32'b11111111110000010000000100010011;
ROM[22423] <= 32'b00000000000000010010010000000011;
ROM[22424] <= 32'b00000000011101000000001110110011;
ROM[22425] <= 32'b00000000011100010010000000100011;
ROM[22426] <= 32'b00000000010000010000000100010011;
ROM[22427] <= 32'b11111111110000010000000100010011;
ROM[22428] <= 32'b00000000000000010010001110000011;
ROM[22429] <= 32'b00000000011100011010001000100011;
ROM[22430] <= 32'b00001000000001101010001110000011;
ROM[22431] <= 32'b00000000011100010010000000100011;
ROM[22432] <= 32'b00000000010000010000000100010011;
ROM[22433] <= 32'b00000000001100000000001110010011;
ROM[22434] <= 32'b00000000011100010010000000100011;
ROM[22435] <= 32'b00000000010000010000000100010011;
ROM[22436] <= 32'b11111111110000010000000100010011;
ROM[22437] <= 32'b00000000000000010010001110000011;
ROM[22438] <= 32'b11111111110000010000000100010011;
ROM[22439] <= 32'b00000000000000010010010000000011;
ROM[22440] <= 32'b00000000011101000111001110110011;
ROM[22441] <= 32'b00000000011100010010000000100011;
ROM[22442] <= 32'b00000000010000010000000100010011;
ROM[22443] <= 32'b11111111110000010000000100010011;
ROM[22444] <= 32'b00000000000000010010001110000011;
ROM[22445] <= 32'b00000000011100011010010000100011;
ROM[22446] <= 32'b00000000000000000000001110010011;
ROM[22447] <= 32'b00000000011100010010000000100011;
ROM[22448] <= 32'b00000000010000010000000100010011;
ROM[22449] <= 32'b11111111110000010000000100010011;
ROM[22450] <= 32'b00000000000000010010001110000011;
ROM[22451] <= 32'b00000000011100011010100000100011;
ROM[22452] <= 32'b00000001000000011010001110000011;
ROM[22453] <= 32'b00000000011100010010000000100011;
ROM[22454] <= 32'b00000000010000010000000100010011;
ROM[22455] <= 32'b00000000100000000000001110010011;
ROM[22456] <= 32'b00000000011100010010000000100011;
ROM[22457] <= 32'b00000000010000010000000100010011;
ROM[22458] <= 32'b11111111110000010000000100010011;
ROM[22459] <= 32'b00000000000000010010001110000011;
ROM[22460] <= 32'b11111111110000010000000100010011;
ROM[22461] <= 32'b00000000000000010010010000000011;
ROM[22462] <= 32'b00000000011101000010001110110011;
ROM[22463] <= 32'b00000000011100010010000000100011;
ROM[22464] <= 32'b00000000010000010000000100010011;
ROM[22465] <= 32'b11111111110000010000000100010011;
ROM[22466] <= 32'b00000000000000010010001110000011;
ROM[22467] <= 32'b01000000011100000000001110110011;
ROM[22468] <= 32'b00000000000100111000001110010011;
ROM[22469] <= 32'b00000000011100010010000000100011;
ROM[22470] <= 32'b00000000010000010000000100010011;
ROM[22471] <= 32'b11111111110000010000000100010011;
ROM[22472] <= 32'b00000000000000010010001110000011;
ROM[22473] <= 32'b00000000000000111000101001100011;
ROM[22474] <= 32'b00000000000000010111001110110111;
ROM[22475] <= 32'b11011101000000111000001110010011;
ROM[22476] <= 32'b00000000111000111000001110110011;
ROM[22477] <= 32'b00000000000000111000000011100111;
ROM[22478] <= 32'b00000001000000011010001110000011;
ROM[22479] <= 32'b00000000011100010010000000100011;
ROM[22480] <= 32'b00000000010000010000000100010011;
ROM[22481] <= 32'b00000000010000000000001110010011;
ROM[22482] <= 32'b00000000011100010010000000100011;
ROM[22483] <= 32'b00000000010000010000000100010011;
ROM[22484] <= 32'b00000000000000010110001110110111;
ROM[22485] <= 32'b11111001110000111000001110010011;
ROM[22486] <= 32'b00000000111000111000001110110011;
ROM[22487] <= 32'b00000000011100010010000000100011;
ROM[22488] <= 32'b00000000010000010000000100010011;
ROM[22489] <= 32'b00000000001100010010000000100011;
ROM[22490] <= 32'b00000000010000010000000100010011;
ROM[22491] <= 32'b00000000010000010010000000100011;
ROM[22492] <= 32'b00000000010000010000000100010011;
ROM[22493] <= 32'b00000000010100010010000000100011;
ROM[22494] <= 32'b00000000010000010000000100010011;
ROM[22495] <= 32'b00000000011000010010000000100011;
ROM[22496] <= 32'b00000000010000010000000100010011;
ROM[22497] <= 32'b00000001010000000000001110010011;
ROM[22498] <= 32'b00000000100000111000001110010011;
ROM[22499] <= 32'b01000000011100010000001110110011;
ROM[22500] <= 32'b00000000011100000000001000110011;
ROM[22501] <= 32'b00000000001000000000000110110011;
ROM[22502] <= 32'b10001001010111111011000011101111;
ROM[22503] <= 32'b11111111110000010000000100010011;
ROM[22504] <= 32'b00000000000000010010001110000011;
ROM[22505] <= 32'b00000000011100011010101000100011;
ROM[22506] <= 32'b00000000000000011010001110000011;
ROM[22507] <= 32'b00000000011100010010000000100011;
ROM[22508] <= 32'b00000000010000010000000100010011;
ROM[22509] <= 32'b00000001010000011010001110000011;
ROM[22510] <= 32'b00000000011100010010000000100011;
ROM[22511] <= 32'b00000000010000010000000100010011;
ROM[22512] <= 32'b11111111110000010000000100010011;
ROM[22513] <= 32'b00000000000000010010001110000011;
ROM[22514] <= 32'b11111111110000010000000100010011;
ROM[22515] <= 32'b00000000000000010010010000000011;
ROM[22516] <= 32'b00000000011101000000001110110011;
ROM[22517] <= 32'b00000000011100010010000000100011;
ROM[22518] <= 32'b00000000010000010000000100010011;
ROM[22519] <= 32'b11111111110000010000000100010011;
ROM[22520] <= 32'b00000000000000010010001110000011;
ROM[22521] <= 32'b00000000000000111000001100010011;
ROM[22522] <= 32'b00000000110100110000010000110011;
ROM[22523] <= 32'b00000000000001000010001110000011;
ROM[22524] <= 32'b00000000011100010010000000100011;
ROM[22525] <= 32'b00000000010000010000000100010011;
ROM[22526] <= 32'b11111111110000010000000100010011;
ROM[22527] <= 32'b00000000000000010010001110000011;
ROM[22528] <= 32'b00000000011100011010011000100011;
ROM[22529] <= 32'b00000000010000011010001110000011;
ROM[22530] <= 32'b00000000011100010010000000100011;
ROM[22531] <= 32'b00000000010000010000000100010011;
ROM[22532] <= 32'b00000000010000000000001110010011;
ROM[22533] <= 32'b00000000011100010010000000100011;
ROM[22534] <= 32'b00000000010000010000000100010011;
ROM[22535] <= 32'b00000000000000010110001110110111;
ROM[22536] <= 32'b00000110100000111000001110010011;
ROM[22537] <= 32'b00000000111000111000001110110011;
ROM[22538] <= 32'b00000000011100010010000000100011;
ROM[22539] <= 32'b00000000010000010000000100010011;
ROM[22540] <= 32'b00000000001100010010000000100011;
ROM[22541] <= 32'b00000000010000010000000100010011;
ROM[22542] <= 32'b00000000010000010010000000100011;
ROM[22543] <= 32'b00000000010000010000000100010011;
ROM[22544] <= 32'b00000000010100010010000000100011;
ROM[22545] <= 32'b00000000010000010000000100010011;
ROM[22546] <= 32'b00000000011000010010000000100011;
ROM[22547] <= 32'b00000000010000010000000100010011;
ROM[22548] <= 32'b00000001010000000000001110010011;
ROM[22549] <= 32'b00000000100000111000001110010011;
ROM[22550] <= 32'b01000000011100010000001110110011;
ROM[22551] <= 32'b00000000011100000000001000110011;
ROM[22552] <= 32'b00000000001000000000000110110011;
ROM[22553] <= 32'b11111100100011111011000011101111;
ROM[22554] <= 32'b11111111110000010000000100010011;
ROM[22555] <= 32'b00000000000000010010001110000011;
ROM[22556] <= 32'b00000000011100011010110000100011;
ROM[22557] <= 32'b00000000100000011010001110000011;
ROM[22558] <= 32'b00000000011100010010000000100011;
ROM[22559] <= 32'b00000000010000010000000100010011;
ROM[22560] <= 32'b00000000000000000000001110010011;
ROM[22561] <= 32'b00000000011100010010000000100011;
ROM[22562] <= 32'b00000000010000010000000100010011;
ROM[22563] <= 32'b11111111110000010000000100010011;
ROM[22564] <= 32'b00000000000000010010001110000011;
ROM[22565] <= 32'b11111111110000010000000100010011;
ROM[22566] <= 32'b00000000000000010010010000000011;
ROM[22567] <= 32'b00000000011101000010010010110011;
ROM[22568] <= 32'b00000000100000111010010100110011;
ROM[22569] <= 32'b00000000101001001000001110110011;
ROM[22570] <= 32'b00000000000100111000001110010011;
ROM[22571] <= 32'b00000000000100111111001110010011;
ROM[22572] <= 32'b00000000011100010010000000100011;
ROM[22573] <= 32'b00000000010000010000000100010011;
ROM[22574] <= 32'b11111111110000010000000100010011;
ROM[22575] <= 32'b00000000000000010010001110000011;
ROM[22576] <= 32'b00000000000000111000101001100011;
ROM[22577] <= 32'b00000000000000010111001110110111;
ROM[22578] <= 32'b10101000100000111000001110010011;
ROM[22579] <= 32'b00000000111000111000001110110011;
ROM[22580] <= 32'b00000000000000111000000011100111;
ROM[22581] <= 32'b00000000100000011010001110000011;
ROM[22582] <= 32'b00000000011100010010000000100011;
ROM[22583] <= 32'b00000000010000010000000100010011;
ROM[22584] <= 32'b00000000000100000000001110010011;
ROM[22585] <= 32'b00000000011100010010000000100011;
ROM[22586] <= 32'b00000000010000010000000100010011;
ROM[22587] <= 32'b11111111110000010000000100010011;
ROM[22588] <= 32'b00000000000000010010001110000011;
ROM[22589] <= 32'b11111111110000010000000100010011;
ROM[22590] <= 32'b00000000000000010010010000000011;
ROM[22591] <= 32'b00000000011101000010010010110011;
ROM[22592] <= 32'b00000000100000111010010100110011;
ROM[22593] <= 32'b00000000101001001000001110110011;
ROM[22594] <= 32'b00000000000100111000001110010011;
ROM[22595] <= 32'b00000000000100111111001110010011;
ROM[22596] <= 32'b00000000011100010010000000100011;
ROM[22597] <= 32'b00000000010000010000000100010011;
ROM[22598] <= 32'b11111111110000010000000100010011;
ROM[22599] <= 32'b00000000000000010010001110000011;
ROM[22600] <= 32'b00000000000000111000101001100011;
ROM[22601] <= 32'b00000000000000010110001110110111;
ROM[22602] <= 32'b01101100110000111000001110010011;
ROM[22603] <= 32'b00000000111000111000001110110011;
ROM[22604] <= 32'b00000000000000111000000011100111;
ROM[22605] <= 32'b00000000100000011010001110000011;
ROM[22606] <= 32'b00000000011100010010000000100011;
ROM[22607] <= 32'b00000000010000010000000100010011;
ROM[22608] <= 32'b00000000001000000000001110010011;
ROM[22609] <= 32'b00000000011100010010000000100011;
ROM[22610] <= 32'b00000000010000010000000100010011;
ROM[22611] <= 32'b11111111110000010000000100010011;
ROM[22612] <= 32'b00000000000000010010001110000011;
ROM[22613] <= 32'b11111111110000010000000100010011;
ROM[22614] <= 32'b00000000000000010010010000000011;
ROM[22615] <= 32'b00000000011101000010010010110011;
ROM[22616] <= 32'b00000000100000111010010100110011;
ROM[22617] <= 32'b00000000101001001000001110110011;
ROM[22618] <= 32'b00000000000100111000001110010011;
ROM[22619] <= 32'b00000000000100111111001110010011;
ROM[22620] <= 32'b00000000011100010010000000100011;
ROM[22621] <= 32'b00000000010000010000000100010011;
ROM[22622] <= 32'b11111111110000010000000100010011;
ROM[22623] <= 32'b00000000000000010010001110000011;
ROM[22624] <= 32'b00000000000000111000101001100011;
ROM[22625] <= 32'b00000000000000010110001110110111;
ROM[22626] <= 32'b00110001000000111000001110010011;
ROM[22627] <= 32'b00000000111000111000001110110011;
ROM[22628] <= 32'b00000000000000111000000011100111;
ROM[22629] <= 32'b00000111110001101010001110000011;
ROM[22630] <= 32'b00000000011100010010000000100011;
ROM[22631] <= 32'b00000000010000010000000100010011;
ROM[22632] <= 32'b00000001100000011010001110000011;
ROM[22633] <= 32'b00000000011100010010000000100011;
ROM[22634] <= 32'b00000000010000010000000100010011;
ROM[22635] <= 32'b11111111110000010000000100010011;
ROM[22636] <= 32'b00000000000000010010001110000011;
ROM[22637] <= 32'b11111111110000010000000100010011;
ROM[22638] <= 32'b00000000000000010010010000000011;
ROM[22639] <= 32'b00000000011101000000001110110011;
ROM[22640] <= 32'b00000000011100010010000000100011;
ROM[22641] <= 32'b00000000010000010000000100010011;
ROM[22642] <= 32'b11111111110000010000000100010011;
ROM[22643] <= 32'b00000000000000010010001110000011;
ROM[22644] <= 32'b00000000000000111000001100010011;
ROM[22645] <= 32'b00000000110100110000010000110011;
ROM[22646] <= 32'b00000000000001000010001110000011;
ROM[22647] <= 32'b00000000011100010010000000100011;
ROM[22648] <= 32'b00000000010000010000000100010011;
ROM[22649] <= 32'b00010000000000000000001110010011;
ROM[22650] <= 32'b00000000011100010010000000100011;
ROM[22651] <= 32'b00000000010000010000000100010011;
ROM[22652] <= 32'b11111111110000010000000100010011;
ROM[22653] <= 32'b00000000000000010010001110000011;
ROM[22654] <= 32'b01000000011100000000001110110011;
ROM[22655] <= 32'b00000000011100010010000000100011;
ROM[22656] <= 32'b00000000010000010000000100010011;
ROM[22657] <= 32'b11111111110000010000000100010011;
ROM[22658] <= 32'b00000000000000010010001110000011;
ROM[22659] <= 32'b11111111110000010000000100010011;
ROM[22660] <= 32'b00000000000000010010010000000011;
ROM[22661] <= 32'b00000000011101000111001110110011;
ROM[22662] <= 32'b00000000011100010010000000100011;
ROM[22663] <= 32'b00000000010000010000000100010011;
ROM[22664] <= 32'b00000000110000011010001110000011;
ROM[22665] <= 32'b00000000011100010010000000100011;
ROM[22666] <= 32'b00000000010000010000000100010011;
ROM[22667] <= 32'b11111111110000010000000100010011;
ROM[22668] <= 32'b00000000000000010010001110000011;
ROM[22669] <= 32'b11111111110000010000000100010011;
ROM[22670] <= 32'b00000000000000010010010000000011;
ROM[22671] <= 32'b00000000011101000110001110110011;
ROM[22672] <= 32'b00000000011100010010000000100011;
ROM[22673] <= 32'b00000000010000010000000100010011;
ROM[22674] <= 32'b11111111110000010000000100010011;
ROM[22675] <= 32'b00000000000000010010001110000011;
ROM[22676] <= 32'b00000010011100011010010000100011;
ROM[22677] <= 32'b00000010100000011010001110000011;
ROM[22678] <= 32'b00000000011100010010000000100011;
ROM[22679] <= 32'b00000000010000010000000100010011;
ROM[22680] <= 32'b00000111100001101010001110000011;
ROM[22681] <= 32'b00000000011100010010000000100011;
ROM[22682] <= 32'b00000000010000010000000100010011;
ROM[22683] <= 32'b00000001100000011010001110000011;
ROM[22684] <= 32'b00000000011100010010000000100011;
ROM[22685] <= 32'b00000000010000010000000100010011;
ROM[22686] <= 32'b11111111110000010000000100010011;
ROM[22687] <= 32'b00000000000000010010001110000011;
ROM[22688] <= 32'b11111111110000010000000100010011;
ROM[22689] <= 32'b00000000000000010010010000000011;
ROM[22690] <= 32'b00000000011101000000001110110011;
ROM[22691] <= 32'b00000000011100010010000000100011;
ROM[22692] <= 32'b00000000010000010000000100010011;
ROM[22693] <= 32'b11111111110000010000000100010011;
ROM[22694] <= 32'b00000000000000010010001110000011;
ROM[22695] <= 32'b00000000000000111000001100010011;
ROM[22696] <= 32'b11111111110000010000000100010011;
ROM[22697] <= 32'b00000000000000010010001110000011;
ROM[22698] <= 32'b00000000110100110000010000110011;
ROM[22699] <= 32'b00000000011101000010000000100011;
ROM[22700] <= 32'b00000010100000011010001110000011;
ROM[22701] <= 32'b00000000011100010010000000100011;
ROM[22702] <= 32'b00000000010000010000000100010011;
ROM[22703] <= 32'b00000111110001101010001110000011;
ROM[22704] <= 32'b00000000011100010010000000100011;
ROM[22705] <= 32'b00000000010000010000000100010011;
ROM[22706] <= 32'b00000001100000011010001110000011;
ROM[22707] <= 32'b00000000011100010010000000100011;
ROM[22708] <= 32'b00000000010000010000000100010011;
ROM[22709] <= 32'b11111111110000010000000100010011;
ROM[22710] <= 32'b00000000000000010010001110000011;
ROM[22711] <= 32'b11111111110000010000000100010011;
ROM[22712] <= 32'b00000000000000010010010000000011;
ROM[22713] <= 32'b00000000011101000000001110110011;
ROM[22714] <= 32'b00000000011100010010000000100011;
ROM[22715] <= 32'b00000000010000010000000100010011;
ROM[22716] <= 32'b11111111110000010000000100010011;
ROM[22717] <= 32'b00000000000000010010001110000011;
ROM[22718] <= 32'b00000000000000111000001100010011;
ROM[22719] <= 32'b11111111110000010000000100010011;
ROM[22720] <= 32'b00000000000000010010001110000011;
ROM[22721] <= 32'b00000000110100110000010000110011;
ROM[22722] <= 32'b00000000011101000010000000100011;
ROM[22723] <= 32'b00111011110000000000000011101111;
ROM[22724] <= 32'b00000001000000000000001110010011;
ROM[22725] <= 32'b00000000011100010010000000100011;
ROM[22726] <= 32'b00000000010000010000000100010011;
ROM[22727] <= 32'b00000000000000010110001110110111;
ROM[22728] <= 32'b00110110100000111000001110010011;
ROM[22729] <= 32'b00000000111000111000001110110011;
ROM[22730] <= 32'b00000000011100010010000000100011;
ROM[22731] <= 32'b00000000010000010000000100010011;
ROM[22732] <= 32'b00000000001100010010000000100011;
ROM[22733] <= 32'b00000000010000010000000100010011;
ROM[22734] <= 32'b00000000010000010010000000100011;
ROM[22735] <= 32'b00000000010000010000000100010011;
ROM[22736] <= 32'b00000000010100010010000000100011;
ROM[22737] <= 32'b00000000010000010000000100010011;
ROM[22738] <= 32'b00000000011000010010000000100011;
ROM[22739] <= 32'b00000000010000010000000100010011;
ROM[22740] <= 32'b00000001010000000000001110010011;
ROM[22741] <= 32'b00000000010000111000001110010011;
ROM[22742] <= 32'b01000000011100010000001110110011;
ROM[22743] <= 32'b00000000011100000000001000110011;
ROM[22744] <= 32'b00000000001000000000000110110011;
ROM[22745] <= 32'b11100000100111111100000011101111;
ROM[22746] <= 32'b00000000100000000000001110010011;
ROM[22747] <= 32'b00000000011100010010000000100011;
ROM[22748] <= 32'b00000000010000010000000100010011;
ROM[22749] <= 32'b00000000000000010110001110110111;
ROM[22750] <= 32'b00111100000000111000001110010011;
ROM[22751] <= 32'b00000000111000111000001110110011;
ROM[22752] <= 32'b00000000011100010010000000100011;
ROM[22753] <= 32'b00000000010000010000000100010011;
ROM[22754] <= 32'b00000000001100010010000000100011;
ROM[22755] <= 32'b00000000010000010000000100010011;
ROM[22756] <= 32'b00000000010000010010000000100011;
ROM[22757] <= 32'b00000000010000010000000100010011;
ROM[22758] <= 32'b00000000010100010010000000100011;
ROM[22759] <= 32'b00000000010000010000000100010011;
ROM[22760] <= 32'b00000000011000010010000000100011;
ROM[22761] <= 32'b00000000010000010000000100010011;
ROM[22762] <= 32'b00000001010000000000001110010011;
ROM[22763] <= 32'b00000000010000111000001110010011;
ROM[22764] <= 32'b01000000011100010000001110110011;
ROM[22765] <= 32'b00000000011100000000001000110011;
ROM[22766] <= 32'b00000000001000000000000110110011;
ROM[22767] <= 32'b11011011000111111100000011101111;
ROM[22768] <= 32'b11111111110000010000000100010011;
ROM[22769] <= 32'b00000000000000010010001110000011;
ROM[22770] <= 32'b11111111110000010000000100010011;
ROM[22771] <= 32'b00000000000000010010010000000011;
ROM[22772] <= 32'b01000000011101000000001110110011;
ROM[22773] <= 32'b00000000011100010010000000100011;
ROM[22774] <= 32'b00000000010000010000000100010011;
ROM[22775] <= 32'b11111111110000010000000100010011;
ROM[22776] <= 32'b00000000000000010010001110000011;
ROM[22777] <= 32'b00000010011100011010000000100011;
ROM[22778] <= 32'b00000000000000000000001110010011;
ROM[22779] <= 32'b00000000011100010010000000100011;
ROM[22780] <= 32'b00000000010000010000000100010011;
ROM[22781] <= 32'b00000010000000011010001110000011;
ROM[22782] <= 32'b00000000011100010010000000100011;
ROM[22783] <= 32'b00000000010000010000000100010011;
ROM[22784] <= 32'b11111111110000010000000100010011;
ROM[22785] <= 32'b00000000000000010010001110000011;
ROM[22786] <= 32'b11111111110000010000000100010011;
ROM[22787] <= 32'b00000000000000010010010000000011;
ROM[22788] <= 32'b01000000011101000000001110110011;
ROM[22789] <= 32'b00000000011100010010000000100011;
ROM[22790] <= 32'b00000000010000010000000100010011;
ROM[22791] <= 32'b11111111110000010000000100010011;
ROM[22792] <= 32'b00000000000000010010001110000011;
ROM[22793] <= 32'b00000010011100011010001000100011;
ROM[22794] <= 32'b00000010010000011010001110000011;
ROM[22795] <= 32'b00000000011100010010000000100011;
ROM[22796] <= 32'b00000000010000010000000100010011;
ROM[22797] <= 32'b00000000000100000000001110010011;
ROM[22798] <= 32'b00000000011100010010000000100011;
ROM[22799] <= 32'b00000000010000010000000100010011;
ROM[22800] <= 32'b11111111110000010000000100010011;
ROM[22801] <= 32'b00000000000000010010001110000011;
ROM[22802] <= 32'b11111111110000010000000100010011;
ROM[22803] <= 32'b00000000000000010010010000000011;
ROM[22804] <= 32'b01000000011101000000001110110011;
ROM[22805] <= 32'b00000000011100010010000000100011;
ROM[22806] <= 32'b00000000010000010000000100010011;
ROM[22807] <= 32'b11111111110000010000000100010011;
ROM[22808] <= 32'b00000000000000010010001110000011;
ROM[22809] <= 32'b00000010011100011010001000100011;
ROM[22810] <= 32'b00000000110000011010001110000011;
ROM[22811] <= 32'b00000000011100010010000000100011;
ROM[22812] <= 32'b00000000010000010000000100010011;
ROM[22813] <= 32'b00000000100000000000001110010011;
ROM[22814] <= 32'b00000000011100010010000000100011;
ROM[22815] <= 32'b00000000010000010000000100010011;
ROM[22816] <= 32'b00000000000000010110001110110111;
ROM[22817] <= 32'b01001100110000111000001110010011;
ROM[22818] <= 32'b00000000111000111000001110110011;
ROM[22819] <= 32'b00000000011100010010000000100011;
ROM[22820] <= 32'b00000000010000010000000100010011;
ROM[22821] <= 32'b00000000001100010010000000100011;
ROM[22822] <= 32'b00000000010000010000000100010011;
ROM[22823] <= 32'b00000000010000010010000000100011;
ROM[22824] <= 32'b00000000010000010000000100010011;
ROM[22825] <= 32'b00000000010100010010000000100011;
ROM[22826] <= 32'b00000000010000010000000100010011;
ROM[22827] <= 32'b00000000011000010010000000100011;
ROM[22828] <= 32'b00000000010000010000000100010011;
ROM[22829] <= 32'b00000001010000000000001110010011;
ROM[22830] <= 32'b00000000010000111000001110010011;
ROM[22831] <= 32'b01000000011100010000001110110011;
ROM[22832] <= 32'b00000000011100000000001000110011;
ROM[22833] <= 32'b00000000001000000000000110110011;
ROM[22834] <= 32'b11001010010111111100000011101111;
ROM[22835] <= 32'b00000000000000010110001110110111;
ROM[22836] <= 32'b01010001100000111000001110010011;
ROM[22837] <= 32'b00000000111000111000001110110011;
ROM[22838] <= 32'b00000000011100010010000000100011;
ROM[22839] <= 32'b00000000010000010000000100010011;
ROM[22840] <= 32'b00000000001100010010000000100011;
ROM[22841] <= 32'b00000000010000010000000100010011;
ROM[22842] <= 32'b00000000010000010010000000100011;
ROM[22843] <= 32'b00000000010000010000000100010011;
ROM[22844] <= 32'b00000000010100010010000000100011;
ROM[22845] <= 32'b00000000010000010000000100010011;
ROM[22846] <= 32'b00000000011000010010000000100011;
ROM[22847] <= 32'b00000000010000010000000100010011;
ROM[22848] <= 32'b00000001010000000000001110010011;
ROM[22849] <= 32'b00000000100000111000001110010011;
ROM[22850] <= 32'b01000000011100010000001110110011;
ROM[22851] <= 32'b00000000011100000000001000110011;
ROM[22852] <= 32'b00000000001000000000000110110011;
ROM[22853] <= 32'b10110001100011111011000011101111;
ROM[22854] <= 32'b11111111110000010000000100010011;
ROM[22855] <= 32'b00000000000000010010001110000011;
ROM[22856] <= 32'b00000000011100011010011000100011;
ROM[22857] <= 32'b00000000110000011010001110000011;
ROM[22858] <= 32'b00000000011100010010000000100011;
ROM[22859] <= 32'b00000000010000010000000100010011;
ROM[22860] <= 32'b00000010000000011010001110000011;
ROM[22861] <= 32'b00000000011100010010000000100011;
ROM[22862] <= 32'b00000000010000010000000100010011;
ROM[22863] <= 32'b11111111110000010000000100010011;
ROM[22864] <= 32'b00000000000000010010001110000011;
ROM[22865] <= 32'b11111111110000010000000100010011;
ROM[22866] <= 32'b00000000000000010010010000000011;
ROM[22867] <= 32'b00000000011101000111001110110011;
ROM[22868] <= 32'b00000000011100010010000000100011;
ROM[22869] <= 32'b00000000010000010000000100010011;
ROM[22870] <= 32'b11111111110000010000000100010011;
ROM[22871] <= 32'b00000000000000010010001110000011;
ROM[22872] <= 32'b00000000011100011010011000100011;
ROM[22873] <= 32'b00000111110001101010001110000011;
ROM[22874] <= 32'b00000000011100010010000000100011;
ROM[22875] <= 32'b00000000010000010000000100010011;
ROM[22876] <= 32'b00000001100000011010001110000011;
ROM[22877] <= 32'b00000000011100010010000000100011;
ROM[22878] <= 32'b00000000010000010000000100010011;
ROM[22879] <= 32'b11111111110000010000000100010011;
ROM[22880] <= 32'b00000000000000010010001110000011;
ROM[22881] <= 32'b11111111110000010000000100010011;
ROM[22882] <= 32'b00000000000000010010010000000011;
ROM[22883] <= 32'b00000000011101000000001110110011;
ROM[22884] <= 32'b00000000011100010010000000100011;
ROM[22885] <= 32'b00000000010000010000000100010011;
ROM[22886] <= 32'b11111111110000010000000100010011;
ROM[22887] <= 32'b00000000000000010010001110000011;
ROM[22888] <= 32'b00000000000000111000001100010011;
ROM[22889] <= 32'b00000000110100110000010000110011;
ROM[22890] <= 32'b00000000000001000010001110000011;
ROM[22891] <= 32'b00000000011100010010000000100011;
ROM[22892] <= 32'b00000000010000010000000100010011;
ROM[22893] <= 32'b00000010010000011010001110000011;
ROM[22894] <= 32'b00000000011100010010000000100011;
ROM[22895] <= 32'b00000000010000010000000100010011;
ROM[22896] <= 32'b11111111110000010000000100010011;
ROM[22897] <= 32'b00000000000000010010001110000011;
ROM[22898] <= 32'b11111111110000010000000100010011;
ROM[22899] <= 32'b00000000000000010010010000000011;
ROM[22900] <= 32'b00000000011101000111001110110011;
ROM[22901] <= 32'b00000000011100010010000000100011;
ROM[22902] <= 32'b00000000010000010000000100010011;
ROM[22903] <= 32'b00000000110000011010001110000011;
ROM[22904] <= 32'b00000000011100010010000000100011;
ROM[22905] <= 32'b00000000010000010000000100010011;
ROM[22906] <= 32'b11111111110000010000000100010011;
ROM[22907] <= 32'b00000000000000010010001110000011;
ROM[22908] <= 32'b11111111110000010000000100010011;
ROM[22909] <= 32'b00000000000000010010010000000011;
ROM[22910] <= 32'b00000000011101000110001110110011;
ROM[22911] <= 32'b00000000011100010010000000100011;
ROM[22912] <= 32'b00000000010000010000000100010011;
ROM[22913] <= 32'b11111111110000010000000100010011;
ROM[22914] <= 32'b00000000000000010010001110000011;
ROM[22915] <= 32'b00000010011100011010010000100011;
ROM[22916] <= 32'b00000010100000011010001110000011;
ROM[22917] <= 32'b00000000011100010010000000100011;
ROM[22918] <= 32'b00000000010000010000000100010011;
ROM[22919] <= 32'b00000111100001101010001110000011;
ROM[22920] <= 32'b00000000011100010010000000100011;
ROM[22921] <= 32'b00000000010000010000000100010011;
ROM[22922] <= 32'b00000001100000011010001110000011;
ROM[22923] <= 32'b00000000011100010010000000100011;
ROM[22924] <= 32'b00000000010000010000000100010011;
ROM[22925] <= 32'b11111111110000010000000100010011;
ROM[22926] <= 32'b00000000000000010010001110000011;
ROM[22927] <= 32'b11111111110000010000000100010011;
ROM[22928] <= 32'b00000000000000010010010000000011;
ROM[22929] <= 32'b00000000011101000000001110110011;
ROM[22930] <= 32'b00000000011100010010000000100011;
ROM[22931] <= 32'b00000000010000010000000100010011;
ROM[22932] <= 32'b11111111110000010000000100010011;
ROM[22933] <= 32'b00000000000000010010001110000011;
ROM[22934] <= 32'b00000000000000111000001100010011;
ROM[22935] <= 32'b11111111110000010000000100010011;
ROM[22936] <= 32'b00000000000000010010001110000011;
ROM[22937] <= 32'b00000000110100110000010000110011;
ROM[22938] <= 32'b00000000011101000010000000100011;
ROM[22939] <= 32'b00000010100000011010001110000011;
ROM[22940] <= 32'b00000000011100010010000000100011;
ROM[22941] <= 32'b00000000010000010000000100010011;
ROM[22942] <= 32'b00000111110001101010001110000011;
ROM[22943] <= 32'b00000000011100010010000000100011;
ROM[22944] <= 32'b00000000010000010000000100010011;
ROM[22945] <= 32'b00000001100000011010001110000011;
ROM[22946] <= 32'b00000000011100010010000000100011;
ROM[22947] <= 32'b00000000010000010000000100010011;
ROM[22948] <= 32'b11111111110000010000000100010011;
ROM[22949] <= 32'b00000000000000010010001110000011;
ROM[22950] <= 32'b11111111110000010000000100010011;
ROM[22951] <= 32'b00000000000000010010010000000011;
ROM[22952] <= 32'b00000000011101000000001110110011;
ROM[22953] <= 32'b00000000011100010010000000100011;
ROM[22954] <= 32'b00000000010000010000000100010011;
ROM[22955] <= 32'b11111111110000010000000100010011;
ROM[22956] <= 32'b00000000000000010010001110000011;
ROM[22957] <= 32'b00000000000000111000001100010011;
ROM[22958] <= 32'b11111111110000010000000100010011;
ROM[22959] <= 32'b00000000000000010010001110000011;
ROM[22960] <= 32'b00000000110100110000010000110011;
ROM[22961] <= 32'b00000000011101000010000000100011;
ROM[22962] <= 32'b00111011110000000000000011101111;
ROM[22963] <= 32'b00000001100000000000001110010011;
ROM[22964] <= 32'b00000000011100010010000000100011;
ROM[22965] <= 32'b00000000010000010000000100010011;
ROM[22966] <= 32'b00000000000000010110001110110111;
ROM[22967] <= 32'b01110010010000111000001110010011;
ROM[22968] <= 32'b00000000111000111000001110110011;
ROM[22969] <= 32'b00000000011100010010000000100011;
ROM[22970] <= 32'b00000000010000010000000100010011;
ROM[22971] <= 32'b00000000001100010010000000100011;
ROM[22972] <= 32'b00000000010000010000000100010011;
ROM[22973] <= 32'b00000000010000010010000000100011;
ROM[22974] <= 32'b00000000010000010000000100010011;
ROM[22975] <= 32'b00000000010100010010000000100011;
ROM[22976] <= 32'b00000000010000010000000100010011;
ROM[22977] <= 32'b00000000011000010010000000100011;
ROM[22978] <= 32'b00000000010000010000000100010011;
ROM[22979] <= 32'b00000001010000000000001110010011;
ROM[22980] <= 32'b00000000010000111000001110010011;
ROM[22981] <= 32'b01000000011100010000001110110011;
ROM[22982] <= 32'b00000000011100000000001000110011;
ROM[22983] <= 32'b00000000001000000000000110110011;
ROM[22984] <= 32'b10100100110111111100000011101111;
ROM[22985] <= 32'b00000001000000000000001110010011;
ROM[22986] <= 32'b00000000011100010010000000100011;
ROM[22987] <= 32'b00000000010000010000000100010011;
ROM[22988] <= 32'b00000000000000010110001110110111;
ROM[22989] <= 32'b01110111110000111000001110010011;
ROM[22990] <= 32'b00000000111000111000001110110011;
ROM[22991] <= 32'b00000000011100010010000000100011;
ROM[22992] <= 32'b00000000010000010000000100010011;
ROM[22993] <= 32'b00000000001100010010000000100011;
ROM[22994] <= 32'b00000000010000010000000100010011;
ROM[22995] <= 32'b00000000010000010010000000100011;
ROM[22996] <= 32'b00000000010000010000000100010011;
ROM[22997] <= 32'b00000000010100010010000000100011;
ROM[22998] <= 32'b00000000010000010000000100010011;
ROM[22999] <= 32'b00000000011000010010000000100011;
ROM[23000] <= 32'b00000000010000010000000100010011;
ROM[23001] <= 32'b00000001010000000000001110010011;
ROM[23002] <= 32'b00000000010000111000001110010011;
ROM[23003] <= 32'b01000000011100010000001110110011;
ROM[23004] <= 32'b00000000011100000000001000110011;
ROM[23005] <= 32'b00000000001000000000000110110011;
ROM[23006] <= 32'b10011111010111111100000011101111;
ROM[23007] <= 32'b11111111110000010000000100010011;
ROM[23008] <= 32'b00000000000000010010001110000011;
ROM[23009] <= 32'b11111111110000010000000100010011;
ROM[23010] <= 32'b00000000000000010010010000000011;
ROM[23011] <= 32'b01000000011101000000001110110011;
ROM[23012] <= 32'b00000000011100010010000000100011;
ROM[23013] <= 32'b00000000010000010000000100010011;
ROM[23014] <= 32'b11111111110000010000000100010011;
ROM[23015] <= 32'b00000000000000010010001110000011;
ROM[23016] <= 32'b00000000011100011010111000100011;
ROM[23017] <= 32'b00000000000000000000001110010011;
ROM[23018] <= 32'b00000000011100010010000000100011;
ROM[23019] <= 32'b00000000010000010000000100010011;
ROM[23020] <= 32'b00000001110000011010001110000011;
ROM[23021] <= 32'b00000000011100010010000000100011;
ROM[23022] <= 32'b00000000010000010000000100010011;
ROM[23023] <= 32'b11111111110000010000000100010011;
ROM[23024] <= 32'b00000000000000010010001110000011;
ROM[23025] <= 32'b11111111110000010000000100010011;
ROM[23026] <= 32'b00000000000000010010010000000011;
ROM[23027] <= 32'b01000000011101000000001110110011;
ROM[23028] <= 32'b00000000011100010010000000100011;
ROM[23029] <= 32'b00000000010000010000000100010011;
ROM[23030] <= 32'b11111111110000010000000100010011;
ROM[23031] <= 32'b00000000000000010010001110000011;
ROM[23032] <= 32'b00000010011100011010001000100011;
ROM[23033] <= 32'b00000010010000011010001110000011;
ROM[23034] <= 32'b00000000011100010010000000100011;
ROM[23035] <= 32'b00000000010000010000000100010011;
ROM[23036] <= 32'b00000000000100000000001110010011;
ROM[23037] <= 32'b00000000011100010010000000100011;
ROM[23038] <= 32'b00000000010000010000000100010011;
ROM[23039] <= 32'b11111111110000010000000100010011;
ROM[23040] <= 32'b00000000000000010010001110000011;
ROM[23041] <= 32'b11111111110000010000000100010011;
ROM[23042] <= 32'b00000000000000010010010000000011;
ROM[23043] <= 32'b01000000011101000000001110110011;
ROM[23044] <= 32'b00000000011100010010000000100011;
ROM[23045] <= 32'b00000000010000010000000100010011;
ROM[23046] <= 32'b11111111110000010000000100010011;
ROM[23047] <= 32'b00000000000000010010001110000011;
ROM[23048] <= 32'b00000010011100011010001000100011;
ROM[23049] <= 32'b00000000110000011010001110000011;
ROM[23050] <= 32'b00000000011100010010000000100011;
ROM[23051] <= 32'b00000000010000010000000100010011;
ROM[23052] <= 32'b00000001000000000000001110010011;
ROM[23053] <= 32'b00000000011100010010000000100011;
ROM[23054] <= 32'b00000000010000010000000100010011;
ROM[23055] <= 32'b00000000000000010111001110110111;
ROM[23056] <= 32'b10001000100000111000001110010011;
ROM[23057] <= 32'b00000000111000111000001110110011;
ROM[23058] <= 32'b00000000011100010010000000100011;
ROM[23059] <= 32'b00000000010000010000000100010011;
ROM[23060] <= 32'b00000000001100010010000000100011;
ROM[23061] <= 32'b00000000010000010000000100010011;
ROM[23062] <= 32'b00000000010000010010000000100011;
ROM[23063] <= 32'b00000000010000010000000100010011;
ROM[23064] <= 32'b00000000010100010010000000100011;
ROM[23065] <= 32'b00000000010000010000000100010011;
ROM[23066] <= 32'b00000000011000010010000000100011;
ROM[23067] <= 32'b00000000010000010000000100010011;
ROM[23068] <= 32'b00000001010000000000001110010011;
ROM[23069] <= 32'b00000000010000111000001110010011;
ROM[23070] <= 32'b01000000011100010000001110110011;
ROM[23071] <= 32'b00000000011100000000001000110011;
ROM[23072] <= 32'b00000000001000000000000110110011;
ROM[23073] <= 32'b10001110100111111100000011101111;
ROM[23074] <= 32'b00000000000000010111001110110111;
ROM[23075] <= 32'b10001101010000111000001110010011;
ROM[23076] <= 32'b00000000111000111000001110110011;
ROM[23077] <= 32'b00000000011100010010000000100011;
ROM[23078] <= 32'b00000000010000010000000100010011;
ROM[23079] <= 32'b00000000001100010010000000100011;
ROM[23080] <= 32'b00000000010000010000000100010011;
ROM[23081] <= 32'b00000000010000010010000000100011;
ROM[23082] <= 32'b00000000010000010000000100010011;
ROM[23083] <= 32'b00000000010100010010000000100011;
ROM[23084] <= 32'b00000000010000010000000100010011;
ROM[23085] <= 32'b00000000011000010010000000100011;
ROM[23086] <= 32'b00000000010000010000000100010011;
ROM[23087] <= 32'b00000001010000000000001110010011;
ROM[23088] <= 32'b00000000100000111000001110010011;
ROM[23089] <= 32'b01000000011100010000001110110011;
ROM[23090] <= 32'b00000000011100000000001000110011;
ROM[23091] <= 32'b00000000001000000000000110110011;
ROM[23092] <= 32'b11110101110111111010000011101111;
ROM[23093] <= 32'b11111111110000010000000100010011;
ROM[23094] <= 32'b00000000000000010010001110000011;
ROM[23095] <= 32'b00000000011100011010011000100011;
ROM[23096] <= 32'b00000000110000011010001110000011;
ROM[23097] <= 32'b00000000011100010010000000100011;
ROM[23098] <= 32'b00000000010000010000000100010011;
ROM[23099] <= 32'b00000001110000011010001110000011;
ROM[23100] <= 32'b00000000011100010010000000100011;
ROM[23101] <= 32'b00000000010000010000000100010011;
ROM[23102] <= 32'b11111111110000010000000100010011;
ROM[23103] <= 32'b00000000000000010010001110000011;
ROM[23104] <= 32'b11111111110000010000000100010011;
ROM[23105] <= 32'b00000000000000010010010000000011;
ROM[23106] <= 32'b00000000011101000111001110110011;
ROM[23107] <= 32'b00000000011100010010000000100011;
ROM[23108] <= 32'b00000000010000010000000100010011;
ROM[23109] <= 32'b11111111110000010000000100010011;
ROM[23110] <= 32'b00000000000000010010001110000011;
ROM[23111] <= 32'b00000000011100011010011000100011;
ROM[23112] <= 32'b00000111110001101010001110000011;
ROM[23113] <= 32'b00000000011100010010000000100011;
ROM[23114] <= 32'b00000000010000010000000100010011;
ROM[23115] <= 32'b00000001100000011010001110000011;
ROM[23116] <= 32'b00000000011100010010000000100011;
ROM[23117] <= 32'b00000000010000010000000100010011;
ROM[23118] <= 32'b11111111110000010000000100010011;
ROM[23119] <= 32'b00000000000000010010001110000011;
ROM[23120] <= 32'b11111111110000010000000100010011;
ROM[23121] <= 32'b00000000000000010010010000000011;
ROM[23122] <= 32'b00000000011101000000001110110011;
ROM[23123] <= 32'b00000000011100010010000000100011;
ROM[23124] <= 32'b00000000010000010000000100010011;
ROM[23125] <= 32'b11111111110000010000000100010011;
ROM[23126] <= 32'b00000000000000010010001110000011;
ROM[23127] <= 32'b00000000000000111000001100010011;
ROM[23128] <= 32'b00000000110100110000010000110011;
ROM[23129] <= 32'b00000000000001000010001110000011;
ROM[23130] <= 32'b00000000011100010010000000100011;
ROM[23131] <= 32'b00000000010000010000000100010011;
ROM[23132] <= 32'b00000010010000011010001110000011;
ROM[23133] <= 32'b00000000011100010010000000100011;
ROM[23134] <= 32'b00000000010000010000000100010011;
ROM[23135] <= 32'b11111111110000010000000100010011;
ROM[23136] <= 32'b00000000000000010010001110000011;
ROM[23137] <= 32'b11111111110000010000000100010011;
ROM[23138] <= 32'b00000000000000010010010000000011;
ROM[23139] <= 32'b00000000011101000111001110110011;
ROM[23140] <= 32'b00000000011100010010000000100011;
ROM[23141] <= 32'b00000000010000010000000100010011;
ROM[23142] <= 32'b00000000110000011010001110000011;
ROM[23143] <= 32'b00000000011100010010000000100011;
ROM[23144] <= 32'b00000000010000010000000100010011;
ROM[23145] <= 32'b11111111110000010000000100010011;
ROM[23146] <= 32'b00000000000000010010001110000011;
ROM[23147] <= 32'b11111111110000010000000100010011;
ROM[23148] <= 32'b00000000000000010010010000000011;
ROM[23149] <= 32'b00000000011101000110001110110011;
ROM[23150] <= 32'b00000000011100010010000000100011;
ROM[23151] <= 32'b00000000010000010000000100010011;
ROM[23152] <= 32'b11111111110000010000000100010011;
ROM[23153] <= 32'b00000000000000010010001110000011;
ROM[23154] <= 32'b00000010011100011010010000100011;
ROM[23155] <= 32'b00000010100000011010001110000011;
ROM[23156] <= 32'b00000000011100010010000000100011;
ROM[23157] <= 32'b00000000010000010000000100010011;
ROM[23158] <= 32'b00000111100001101010001110000011;
ROM[23159] <= 32'b00000000011100010010000000100011;
ROM[23160] <= 32'b00000000010000010000000100010011;
ROM[23161] <= 32'b00000001100000011010001110000011;
ROM[23162] <= 32'b00000000011100010010000000100011;
ROM[23163] <= 32'b00000000010000010000000100010011;
ROM[23164] <= 32'b11111111110000010000000100010011;
ROM[23165] <= 32'b00000000000000010010001110000011;
ROM[23166] <= 32'b11111111110000010000000100010011;
ROM[23167] <= 32'b00000000000000010010010000000011;
ROM[23168] <= 32'b00000000011101000000001110110011;
ROM[23169] <= 32'b00000000011100010010000000100011;
ROM[23170] <= 32'b00000000010000010000000100010011;
ROM[23171] <= 32'b11111111110000010000000100010011;
ROM[23172] <= 32'b00000000000000010010001110000011;
ROM[23173] <= 32'b00000000000000111000001100010011;
ROM[23174] <= 32'b11111111110000010000000100010011;
ROM[23175] <= 32'b00000000000000010010001110000011;
ROM[23176] <= 32'b00000000110100110000010000110011;
ROM[23177] <= 32'b00000000011101000010000000100011;
ROM[23178] <= 32'b00000010100000011010001110000011;
ROM[23179] <= 32'b00000000011100010010000000100011;
ROM[23180] <= 32'b00000000010000010000000100010011;
ROM[23181] <= 32'b00000111110001101010001110000011;
ROM[23182] <= 32'b00000000011100010010000000100011;
ROM[23183] <= 32'b00000000010000010000000100010011;
ROM[23184] <= 32'b00000001100000011010001110000011;
ROM[23185] <= 32'b00000000011100010010000000100011;
ROM[23186] <= 32'b00000000010000010000000100010011;
ROM[23187] <= 32'b11111111110000010000000100010011;
ROM[23188] <= 32'b00000000000000010010001110000011;
ROM[23189] <= 32'b11111111110000010000000100010011;
ROM[23190] <= 32'b00000000000000010010010000000011;
ROM[23191] <= 32'b00000000011101000000001110110011;
ROM[23192] <= 32'b00000000011100010010000000100011;
ROM[23193] <= 32'b00000000010000010000000100010011;
ROM[23194] <= 32'b11111111110000010000000100010011;
ROM[23195] <= 32'b00000000000000010010001110000011;
ROM[23196] <= 32'b00000000000000111000001100010011;
ROM[23197] <= 32'b11111111110000010000000100010011;
ROM[23198] <= 32'b00000000000000010010001110000011;
ROM[23199] <= 32'b00000000110100110000010000110011;
ROM[23200] <= 32'b00000000011101000010000000100011;
ROM[23201] <= 32'b00101100100000000000000011101111;
ROM[23202] <= 32'b00000001100000000000001110010011;
ROM[23203] <= 32'b00000000011100010010000000100011;
ROM[23204] <= 32'b00000000010000010000000100010011;
ROM[23205] <= 32'b00000000000000010111001110110111;
ROM[23206] <= 32'b10101110000000111000001110010011;
ROM[23207] <= 32'b00000000111000111000001110110011;
ROM[23208] <= 32'b00000000011100010010000000100011;
ROM[23209] <= 32'b00000000010000010000000100010011;
ROM[23210] <= 32'b00000000001100010010000000100011;
ROM[23211] <= 32'b00000000010000010000000100010011;
ROM[23212] <= 32'b00000000010000010010000000100011;
ROM[23213] <= 32'b00000000010000010000000100010011;
ROM[23214] <= 32'b00000000010100010010000000100011;
ROM[23215] <= 32'b00000000010000010000000100010011;
ROM[23216] <= 32'b00000000011000010010000000100011;
ROM[23217] <= 32'b00000000010000010000000100010011;
ROM[23218] <= 32'b00000001010000000000001110010011;
ROM[23219] <= 32'b00000000010000111000001110010011;
ROM[23220] <= 32'b01000000011100010000001110110011;
ROM[23221] <= 32'b00000000011100000000001000110011;
ROM[23222] <= 32'b00000000001000000000000110110011;
ROM[23223] <= 32'b11101001000011111100000011101111;
ROM[23224] <= 32'b11111111110000010000000100010011;
ROM[23225] <= 32'b00000000000000010010001110000011;
ROM[23226] <= 32'b00000010011100011010001000100011;
ROM[23227] <= 32'b00000000110000011010001110000011;
ROM[23228] <= 32'b00000000011100010010000000100011;
ROM[23229] <= 32'b00000000010000010000000100010011;
ROM[23230] <= 32'b00000001100000000000001110010011;
ROM[23231] <= 32'b00000000011100010010000000100011;
ROM[23232] <= 32'b00000000010000010000000100010011;
ROM[23233] <= 32'b00000000000000010111001110110111;
ROM[23234] <= 32'b10110101000000111000001110010011;
ROM[23235] <= 32'b00000000111000111000001110110011;
ROM[23236] <= 32'b00000000011100010010000000100011;
ROM[23237] <= 32'b00000000010000010000000100010011;
ROM[23238] <= 32'b00000000001100010010000000100011;
ROM[23239] <= 32'b00000000010000010000000100010011;
ROM[23240] <= 32'b00000000010000010010000000100011;
ROM[23241] <= 32'b00000000010000010000000100010011;
ROM[23242] <= 32'b00000000010100010010000000100011;
ROM[23243] <= 32'b00000000010000010000000100010011;
ROM[23244] <= 32'b00000000011000010010000000100011;
ROM[23245] <= 32'b00000000010000010000000100010011;
ROM[23246] <= 32'b00000001010000000000001110010011;
ROM[23247] <= 32'b00000000010000111000001110010011;
ROM[23248] <= 32'b01000000011100010000001110110011;
ROM[23249] <= 32'b00000000011100000000001000110011;
ROM[23250] <= 32'b00000000001000000000000110110011;
ROM[23251] <= 32'b11100010000011111100000011101111;
ROM[23252] <= 32'b00000000000000010111001110110111;
ROM[23253] <= 32'b10111001110000111000001110010011;
ROM[23254] <= 32'b00000000111000111000001110110011;
ROM[23255] <= 32'b00000000011100010010000000100011;
ROM[23256] <= 32'b00000000010000010000000100010011;
ROM[23257] <= 32'b00000000001100010010000000100011;
ROM[23258] <= 32'b00000000010000010000000100010011;
ROM[23259] <= 32'b00000000010000010010000000100011;
ROM[23260] <= 32'b00000000010000010000000100010011;
ROM[23261] <= 32'b00000000010100010010000000100011;
ROM[23262] <= 32'b00000000010000010000000100010011;
ROM[23263] <= 32'b00000000011000010010000000100011;
ROM[23264] <= 32'b00000000010000010000000100010011;
ROM[23265] <= 32'b00000001010000000000001110010011;
ROM[23266] <= 32'b00000000100000111000001110010011;
ROM[23267] <= 32'b01000000011100010000001110110011;
ROM[23268] <= 32'b00000000011100000000001000110011;
ROM[23269] <= 32'b00000000001000000000000110110011;
ROM[23270] <= 32'b11001001010111111010000011101111;
ROM[23271] <= 32'b11111111110000010000000100010011;
ROM[23272] <= 32'b00000000000000010010001110000011;
ROM[23273] <= 32'b00000000011100011010011000100011;
ROM[23274] <= 32'b00000010010000011010001110000011;
ROM[23275] <= 32'b00000000011100010010000000100011;
ROM[23276] <= 32'b00000000010000010000000100010011;
ROM[23277] <= 32'b00000000000100000000001110010011;
ROM[23278] <= 32'b00000000011100010010000000100011;
ROM[23279] <= 32'b00000000010000010000000100010011;
ROM[23280] <= 32'b11111111110000010000000100010011;
ROM[23281] <= 32'b00000000000000010010001110000011;
ROM[23282] <= 32'b11111111110000010000000100010011;
ROM[23283] <= 32'b00000000000000010010010000000011;
ROM[23284] <= 32'b01000000011101000000001110110011;
ROM[23285] <= 32'b00000000011100010010000000100011;
ROM[23286] <= 32'b00000000010000010000000100010011;
ROM[23287] <= 32'b11111111110000010000000100010011;
ROM[23288] <= 32'b00000000000000010010001110000011;
ROM[23289] <= 32'b00000010011100011010001000100011;
ROM[23290] <= 32'b00000111110001101010001110000011;
ROM[23291] <= 32'b00000000011100010010000000100011;
ROM[23292] <= 32'b00000000010000010000000100010011;
ROM[23293] <= 32'b00000001100000011010001110000011;
ROM[23294] <= 32'b00000000011100010010000000100011;
ROM[23295] <= 32'b00000000010000010000000100010011;
ROM[23296] <= 32'b11111111110000010000000100010011;
ROM[23297] <= 32'b00000000000000010010001110000011;
ROM[23298] <= 32'b11111111110000010000000100010011;
ROM[23299] <= 32'b00000000000000010010010000000011;
ROM[23300] <= 32'b00000000011101000000001110110011;
ROM[23301] <= 32'b00000000011100010010000000100011;
ROM[23302] <= 32'b00000000010000010000000100010011;
ROM[23303] <= 32'b11111111110000010000000100010011;
ROM[23304] <= 32'b00000000000000010010001110000011;
ROM[23305] <= 32'b00000000000000111000001100010011;
ROM[23306] <= 32'b00000000110100110000010000110011;
ROM[23307] <= 32'b00000000000001000010001110000011;
ROM[23308] <= 32'b00000000011100010010000000100011;
ROM[23309] <= 32'b00000000010000010000000100010011;
ROM[23310] <= 32'b00000010010000011010001110000011;
ROM[23311] <= 32'b00000000011100010010000000100011;
ROM[23312] <= 32'b00000000010000010000000100010011;
ROM[23313] <= 32'b11111111110000010000000100010011;
ROM[23314] <= 32'b00000000000000010010001110000011;
ROM[23315] <= 32'b11111111110000010000000100010011;
ROM[23316] <= 32'b00000000000000010010010000000011;
ROM[23317] <= 32'b00000000011101000111001110110011;
ROM[23318] <= 32'b00000000011100010010000000100011;
ROM[23319] <= 32'b00000000010000010000000100010011;
ROM[23320] <= 32'b00000000110000011010001110000011;
ROM[23321] <= 32'b00000000011100010010000000100011;
ROM[23322] <= 32'b00000000010000010000000100010011;
ROM[23323] <= 32'b11111111110000010000000100010011;
ROM[23324] <= 32'b00000000000000010010001110000011;
ROM[23325] <= 32'b11111111110000010000000100010011;
ROM[23326] <= 32'b00000000000000010010010000000011;
ROM[23327] <= 32'b00000000011101000110001110110011;
ROM[23328] <= 32'b00000000011100010010000000100011;
ROM[23329] <= 32'b00000000010000010000000100010011;
ROM[23330] <= 32'b11111111110000010000000100010011;
ROM[23331] <= 32'b00000000000000010010001110000011;
ROM[23332] <= 32'b00000010011100011010010000100011;
ROM[23333] <= 32'b00000010100000011010001110000011;
ROM[23334] <= 32'b00000000011100010010000000100011;
ROM[23335] <= 32'b00000000010000010000000100010011;
ROM[23336] <= 32'b00000111100001101010001110000011;
ROM[23337] <= 32'b00000000011100010010000000100011;
ROM[23338] <= 32'b00000000010000010000000100010011;
ROM[23339] <= 32'b00000001100000011010001110000011;
ROM[23340] <= 32'b00000000011100010010000000100011;
ROM[23341] <= 32'b00000000010000010000000100010011;
ROM[23342] <= 32'b11111111110000010000000100010011;
ROM[23343] <= 32'b00000000000000010010001110000011;
ROM[23344] <= 32'b11111111110000010000000100010011;
ROM[23345] <= 32'b00000000000000010010010000000011;
ROM[23346] <= 32'b00000000011101000000001110110011;
ROM[23347] <= 32'b00000000011100010010000000100011;
ROM[23348] <= 32'b00000000010000010000000100010011;
ROM[23349] <= 32'b11111111110000010000000100010011;
ROM[23350] <= 32'b00000000000000010010001110000011;
ROM[23351] <= 32'b00000000000000111000001100010011;
ROM[23352] <= 32'b11111111110000010000000100010011;
ROM[23353] <= 32'b00000000000000010010001110000011;
ROM[23354] <= 32'b00000000110100110000010000110011;
ROM[23355] <= 32'b00000000011101000010000000100011;
ROM[23356] <= 32'b00000010100000011010001110000011;
ROM[23357] <= 32'b00000000011100010010000000100011;
ROM[23358] <= 32'b00000000010000010000000100010011;
ROM[23359] <= 32'b00000111110001101010001110000011;
ROM[23360] <= 32'b00000000011100010010000000100011;
ROM[23361] <= 32'b00000000010000010000000100010011;
ROM[23362] <= 32'b00000001100000011010001110000011;
ROM[23363] <= 32'b00000000011100010010000000100011;
ROM[23364] <= 32'b00000000010000010000000100010011;
ROM[23365] <= 32'b11111111110000010000000100010011;
ROM[23366] <= 32'b00000000000000010010001110000011;
ROM[23367] <= 32'b11111111110000010000000100010011;
ROM[23368] <= 32'b00000000000000010010010000000011;
ROM[23369] <= 32'b00000000011101000000001110110011;
ROM[23370] <= 32'b00000000011100010010000000100011;
ROM[23371] <= 32'b00000000010000010000000100010011;
ROM[23372] <= 32'b11111111110000010000000100010011;
ROM[23373] <= 32'b00000000000000010010001110000011;
ROM[23374] <= 32'b00000000000000111000001100010011;
ROM[23375] <= 32'b11111111110000010000000100010011;
ROM[23376] <= 32'b00000000000000010010001110000011;
ROM[23377] <= 32'b00000000110100110000010000110011;
ROM[23378] <= 32'b00000000011101000010000000100011;
ROM[23379] <= 32'b00000000010000011010001110000011;
ROM[23380] <= 32'b00000000011100010010000000100011;
ROM[23381] <= 32'b00000000010000010000000100010011;
ROM[23382] <= 32'b00000000101000000000001110010011;
ROM[23383] <= 32'b00000000011100010010000000100011;
ROM[23384] <= 32'b00000000010000010000000100010011;
ROM[23385] <= 32'b11111111110000010000000100010011;
ROM[23386] <= 32'b00000000000000010010001110000011;
ROM[23387] <= 32'b11111111110000010000000100010011;
ROM[23388] <= 32'b00000000000000010010010000000011;
ROM[23389] <= 32'b00000000011101000000001110110011;
ROM[23390] <= 32'b00000000011100010010000000100011;
ROM[23391] <= 32'b00000000010000010000000100010011;
ROM[23392] <= 32'b11111111110000010000000100010011;
ROM[23393] <= 32'b00000000000000010010001110000011;
ROM[23394] <= 32'b00000000011100011010001000100011;
ROM[23395] <= 32'b00000001000000011010001110000011;
ROM[23396] <= 32'b00000000011100010010000000100011;
ROM[23397] <= 32'b00000000010000010000000100010011;
ROM[23398] <= 32'b00000000000100000000001110010011;
ROM[23399] <= 32'b00000000011100010010000000100011;
ROM[23400] <= 32'b00000000010000010000000100010011;
ROM[23401] <= 32'b11111111110000010000000100010011;
ROM[23402] <= 32'b00000000000000010010001110000011;
ROM[23403] <= 32'b11111111110000010000000100010011;
ROM[23404] <= 32'b00000000000000010010010000000011;
ROM[23405] <= 32'b00000000011101000000001110110011;
ROM[23406] <= 32'b00000000011100010010000000100011;
ROM[23407] <= 32'b00000000010000010000000100010011;
ROM[23408] <= 32'b11111111110000010000000100010011;
ROM[23409] <= 32'b00000000000000010010001110000011;
ROM[23410] <= 32'b00000000011100011010100000100011;
ROM[23411] <= 32'b10010000010011111111000011101111;
ROM[23412] <= 32'b00001000000001101010001110000011;
ROM[23413] <= 32'b00000000011100010010000000100011;
ROM[23414] <= 32'b00000000010000010000000100010011;
ROM[23415] <= 32'b00000010011100000000001110010011;
ROM[23416] <= 32'b00000000011100010010000000100011;
ROM[23417] <= 32'b00000000010000010000000100010011;
ROM[23418] <= 32'b11111111110000010000000100010011;
ROM[23419] <= 32'b00000000000000010010001110000011;
ROM[23420] <= 32'b11111111110000010000000100010011;
ROM[23421] <= 32'b00000000000000010010010000000011;
ROM[23422] <= 32'b00000000011101000010010010110011;
ROM[23423] <= 32'b00000000100000111010010100110011;
ROM[23424] <= 32'b00000000101001001000001110110011;
ROM[23425] <= 32'b00000000000100111000001110010011;
ROM[23426] <= 32'b00000000000100111111001110010011;
ROM[23427] <= 32'b00000000011100010010000000100011;
ROM[23428] <= 32'b00000000010000010000000100010011;
ROM[23429] <= 32'b11111111110000010000000100010011;
ROM[23430] <= 32'b00000000000000010010001110000011;
ROM[23431] <= 32'b00000000000000111000101001100011;
ROM[23432] <= 32'b00000000000000010111001110110111;
ROM[23433] <= 32'b11101100110000111000001110010011;
ROM[23434] <= 32'b00000000111000111000001110110011;
ROM[23435] <= 32'b00000000000000111000000011100111;
ROM[23436] <= 32'b00001000010001101010001110000011;
ROM[23437] <= 32'b00000000011100010010000000100011;
ROM[23438] <= 32'b00000000010000010000000100010011;
ROM[23439] <= 32'b00001000000001101010001110000011;
ROM[23440] <= 32'b00000000011100010010000000100011;
ROM[23441] <= 32'b00000000010000010000000100010011;
ROM[23442] <= 32'b00000000000100000000001110010011;
ROM[23443] <= 32'b00000000011100010010000000100011;
ROM[23444] <= 32'b00000000010000010000000100010011;
ROM[23445] <= 32'b11111111110000010000000100010011;
ROM[23446] <= 32'b00000000000000010010001110000011;
ROM[23447] <= 32'b11111111110000010000000100010011;
ROM[23448] <= 32'b00000000000000010010010000000011;
ROM[23449] <= 32'b00000000011101000000001110110011;
ROM[23450] <= 32'b00000000011100010010000000100011;
ROM[23451] <= 32'b00000000010000010000000100010011;
ROM[23452] <= 32'b00000000000000010111001110110111;
ROM[23453] <= 32'b11101011110000111000001110010011;
ROM[23454] <= 32'b00000000111000111000001110110011;
ROM[23455] <= 32'b00000000011100010010000000100011;
ROM[23456] <= 32'b00000000010000010000000100010011;
ROM[23457] <= 32'b00000000001100010010000000100011;
ROM[23458] <= 32'b00000000010000010000000100010011;
ROM[23459] <= 32'b00000000010000010010000000100011;
ROM[23460] <= 32'b00000000010000010000000100010011;
ROM[23461] <= 32'b00000000010100010010000000100011;
ROM[23462] <= 32'b00000000010000010000000100010011;
ROM[23463] <= 32'b00000000011000010010000000100011;
ROM[23464] <= 32'b00000000010000010000000100010011;
ROM[23465] <= 32'b00000001010000000000001110010011;
ROM[23466] <= 32'b00000000100000111000001110010011;
ROM[23467] <= 32'b01000000011100010000001110110011;
ROM[23468] <= 32'b00000000011100000000001000110011;
ROM[23469] <= 32'b00000000001000000000000110110011;
ROM[23470] <= 32'b11010100100111111110000011101111;
ROM[23471] <= 32'b11111111110000010000000100010011;
ROM[23472] <= 32'b00000000000000010010001110000011;
ROM[23473] <= 32'b00000000011101100010000000100011;
ROM[23474] <= 32'b00000101110000000000000011101111;
ROM[23475] <= 32'b00000000000000010111001110110111;
ROM[23476] <= 32'b11110001100000111000001110010011;
ROM[23477] <= 32'b00000000111000111000001110110011;
ROM[23478] <= 32'b00000000011100010010000000100011;
ROM[23479] <= 32'b00000000010000010000000100010011;
ROM[23480] <= 32'b00000000001100010010000000100011;
ROM[23481] <= 32'b00000000010000010000000100010011;
ROM[23482] <= 32'b00000000010000010010000000100011;
ROM[23483] <= 32'b00000000010000010000000100010011;
ROM[23484] <= 32'b00000000010100010010000000100011;
ROM[23485] <= 32'b00000000010000010000000100010011;
ROM[23486] <= 32'b00000000011000010010000000100011;
ROM[23487] <= 32'b00000000010000010000000100010011;
ROM[23488] <= 32'b00000001010000000000001110010011;
ROM[23489] <= 32'b00000000000000111000001110010011;
ROM[23490] <= 32'b01000000011100010000001110110011;
ROM[23491] <= 32'b00000000011100000000001000110011;
ROM[23492] <= 32'b00000000001000000000000110110011;
ROM[23493] <= 32'b01000101010000000000000011101111;
ROM[23494] <= 32'b11111111110000010000000100010011;
ROM[23495] <= 32'b00000000000000010010001110000011;
ROM[23496] <= 32'b00000000011101100010000000100011;
ROM[23497] <= 32'b00000000000000000000001110010011;
ROM[23498] <= 32'b00000000011100010010000000100011;
ROM[23499] <= 32'b00000000010000010000000100010011;
ROM[23500] <= 32'b00000001010000000000001110010011;
ROM[23501] <= 32'b01000000011100011000001110110011;
ROM[23502] <= 32'b00000000000000111010000010000011;
ROM[23503] <= 32'b11111111110000010000000100010011;
ROM[23504] <= 32'b00000000000000010010001110000011;
ROM[23505] <= 32'b00000000011100100010000000100011;
ROM[23506] <= 32'b00000000010000100000000100010011;
ROM[23507] <= 32'b00000001010000000000001110010011;
ROM[23508] <= 32'b01000000011100011000001110110011;
ROM[23509] <= 32'b00000000010000111010000110000011;
ROM[23510] <= 32'b00000000100000111010001000000011;
ROM[23511] <= 32'b00000000110000111010001010000011;
ROM[23512] <= 32'b00000001000000111010001100000011;
ROM[23513] <= 32'b00000000000000001000000011100111;
ROM[23514] <= 32'b00000000000000010010000000100011;
ROM[23515] <= 32'b00000000010000010000000100010011;
ROM[23516] <= 32'b00000000000000000000001110010011;
ROM[23517] <= 32'b00000000011100010010000000100011;
ROM[23518] <= 32'b00000000010000010000000100010011;
ROM[23519] <= 32'b11111111110000010000000100010011;
ROM[23520] <= 32'b00000000000000010010001110000011;
ROM[23521] <= 32'b00000000011100011010000000100011;
ROM[23522] <= 32'b00000000000000011010001110000011;
ROM[23523] <= 32'b00000000011100010010000000100011;
ROM[23524] <= 32'b00000000010000010000000100010011;
ROM[23525] <= 32'b00000000000000100010001110000011;
ROM[23526] <= 32'b00000000011100010010000000100011;
ROM[23527] <= 32'b00000000010000010000000100010011;
ROM[23528] <= 32'b00000000000000010111001110110111;
ROM[23529] <= 32'b11111110110000111000001110010011;
ROM[23530] <= 32'b00000000111000111000001110110011;
ROM[23531] <= 32'b00000000011100010010000000100011;
ROM[23532] <= 32'b00000000010000010000000100010011;
ROM[23533] <= 32'b00000000001100010010000000100011;
ROM[23534] <= 32'b00000000010000010000000100010011;
ROM[23535] <= 32'b00000000010000010010000000100011;
ROM[23536] <= 32'b00000000010000010000000100010011;
ROM[23537] <= 32'b00000000010100010010000000100011;
ROM[23538] <= 32'b00000000010000010000000100010011;
ROM[23539] <= 32'b00000000011000010010000000100011;
ROM[23540] <= 32'b00000000010000010000000100010011;
ROM[23541] <= 32'b00000001010000000000001110010011;
ROM[23542] <= 32'b00000000010000111000001110010011;
ROM[23543] <= 32'b01000000011100010000001110110011;
ROM[23544] <= 32'b00000000011100000000001000110011;
ROM[23545] <= 32'b00000000001000000000000110110011;
ROM[23546] <= 32'b00010001010100010010000011101111;
ROM[23547] <= 32'b11111111110000010000000100010011;
ROM[23548] <= 32'b00000000000000010010001110000011;
ROM[23549] <= 32'b11111111110000010000000100010011;
ROM[23550] <= 32'b00000000000000010010010000000011;
ROM[23551] <= 32'b00000000011101000010001110110011;
ROM[23552] <= 32'b00000000011100010010000000100011;
ROM[23553] <= 32'b00000000010000010000000100010011;
ROM[23554] <= 32'b11111111110000010000000100010011;
ROM[23555] <= 32'b00000000000000010010001110000011;
ROM[23556] <= 32'b01000000011100000000001110110011;
ROM[23557] <= 32'b00000000000100111000001110010011;
ROM[23558] <= 32'b00000000011100010010000000100011;
ROM[23559] <= 32'b00000000010000010000000100010011;
ROM[23560] <= 32'b11111111110000010000000100010011;
ROM[23561] <= 32'b00000000000000010010001110000011;
ROM[23562] <= 32'b00000000000000111000101001100011;
ROM[23563] <= 32'b00000000000000010111001110110111;
ROM[23564] <= 32'b00010011110000111000001110010011;
ROM[23565] <= 32'b00000000111000111000001110110011;
ROM[23566] <= 32'b00000000000000111000000011100111;
ROM[23567] <= 32'b00000000000000100010001110000011;
ROM[23568] <= 32'b00000000011100010010000000100011;
ROM[23569] <= 32'b00000000010000010000000100010011;
ROM[23570] <= 32'b00000000000000011010001110000011;
ROM[23571] <= 32'b00000000011100010010000000100011;
ROM[23572] <= 32'b00000000010000010000000100010011;
ROM[23573] <= 32'b00000000000000010111001110110111;
ROM[23574] <= 32'b00001010000000111000001110010011;
ROM[23575] <= 32'b00000000111000111000001110110011;
ROM[23576] <= 32'b00000000011100010010000000100011;
ROM[23577] <= 32'b00000000010000010000000100010011;
ROM[23578] <= 32'b00000000001100010010000000100011;
ROM[23579] <= 32'b00000000010000010000000100010011;
ROM[23580] <= 32'b00000000010000010010000000100011;
ROM[23581] <= 32'b00000000010000010000000100010011;
ROM[23582] <= 32'b00000000010100010010000000100011;
ROM[23583] <= 32'b00000000010000010000000100010011;
ROM[23584] <= 32'b00000000011000010010000000100011;
ROM[23585] <= 32'b00000000010000010000000100010011;
ROM[23586] <= 32'b00000001010000000000001110010011;
ROM[23587] <= 32'b00000000100000111000001110010011;
ROM[23588] <= 32'b01000000011100010000001110110011;
ROM[23589] <= 32'b00000000011100000000001000110011;
ROM[23590] <= 32'b00000000001000000000000110110011;
ROM[23591] <= 32'b00001100000100010010000011101111;
ROM[23592] <= 32'b00000000000000010111001110110111;
ROM[23593] <= 32'b00001110110000111000001110010011;
ROM[23594] <= 32'b00000000111000111000001110110011;
ROM[23595] <= 32'b00000000011100010010000000100011;
ROM[23596] <= 32'b00000000010000010000000100010011;
ROM[23597] <= 32'b00000000001100010010000000100011;
ROM[23598] <= 32'b00000000010000010000000100010011;
ROM[23599] <= 32'b00000000010000010010000000100011;
ROM[23600] <= 32'b00000000010000010000000100010011;
ROM[23601] <= 32'b00000000010100010010000000100011;
ROM[23602] <= 32'b00000000010000010000000100010011;
ROM[23603] <= 32'b00000000011000010010000000100011;
ROM[23604] <= 32'b00000000010000010000000100010011;
ROM[23605] <= 32'b00000001010000000000001110010011;
ROM[23606] <= 32'b00000000010000111000001110010011;
ROM[23607] <= 32'b01000000011100010000001110110011;
ROM[23608] <= 32'b00000000011100000000001000110011;
ROM[23609] <= 32'b00000000001000000000000110110011;
ROM[23610] <= 32'b10111000110111111110000011101111;
ROM[23611] <= 32'b11111111110000010000000100010011;
ROM[23612] <= 32'b00000000000000010010001110000011;
ROM[23613] <= 32'b00000000011101100010000000100011;
ROM[23614] <= 32'b00000000000000011010001110000011;
ROM[23615] <= 32'b00000000011100010010000000100011;
ROM[23616] <= 32'b00000000010000010000000100010011;
ROM[23617] <= 32'b00000000000100000000001110010011;
ROM[23618] <= 32'b00000000011100010010000000100011;
ROM[23619] <= 32'b00000000010000010000000100010011;
ROM[23620] <= 32'b11111111110000010000000100010011;
ROM[23621] <= 32'b00000000000000010010001110000011;
ROM[23622] <= 32'b11111111110000010000000100010011;
ROM[23623] <= 32'b00000000000000010010010000000011;
ROM[23624] <= 32'b00000000011101000000001110110011;
ROM[23625] <= 32'b00000000011100010010000000100011;
ROM[23626] <= 32'b00000000010000010000000100010011;
ROM[23627] <= 32'b11111111110000010000000100010011;
ROM[23628] <= 32'b00000000000000010010001110000011;
ROM[23629] <= 32'b00000000011100011010000000100011;
ROM[23630] <= 32'b11100101000111111111000011101111;
ROM[23631] <= 32'b00000000000000000000001110010011;
ROM[23632] <= 32'b00000000011100010010000000100011;
ROM[23633] <= 32'b00000000010000010000000100010011;
ROM[23634] <= 32'b00000001010000000000001110010011;
ROM[23635] <= 32'b01000000011100011000001110110011;
ROM[23636] <= 32'b00000000000000111010000010000011;
ROM[23637] <= 32'b11111111110000010000000100010011;
ROM[23638] <= 32'b00000000000000010010001110000011;
ROM[23639] <= 32'b00000000011100100010000000100011;
ROM[23640] <= 32'b00000000010000100000000100010011;
ROM[23641] <= 32'b00000001010000000000001110010011;
ROM[23642] <= 32'b01000000011100011000001110110011;
ROM[23643] <= 32'b00000000010000111010000110000011;
ROM[23644] <= 32'b00000000100000111010001000000011;
ROM[23645] <= 32'b00000000110000111010001010000011;
ROM[23646] <= 32'b00000001000000111010001100000011;
ROM[23647] <= 32'b00000000000000001000000011100111;
ROM[23648] <= 32'b00000000000000010010000000100011;
ROM[23649] <= 32'b00000000010000010000000100010011;
ROM[23650] <= 32'b00000000101000000000001110010011;
ROM[23651] <= 32'b00000000011100010010000000100011;
ROM[23652] <= 32'b00000000010000010000000100010011;
ROM[23653] <= 32'b00000000000000010111001110110111;
ROM[23654] <= 32'b00011110000000111000001110010011;
ROM[23655] <= 32'b00000000111000111000001110110011;
ROM[23656] <= 32'b00000000011100010010000000100011;
ROM[23657] <= 32'b00000000010000010000000100010011;
ROM[23658] <= 32'b00000000001100010010000000100011;
ROM[23659] <= 32'b00000000010000010000000100010011;
ROM[23660] <= 32'b00000000010000010010000000100011;
ROM[23661] <= 32'b00000000010000010000000100010011;
ROM[23662] <= 32'b00000000010100010010000000100011;
ROM[23663] <= 32'b00000000010000010000000100010011;
ROM[23664] <= 32'b00000000011000010010000000100011;
ROM[23665] <= 32'b00000000010000010000000100010011;
ROM[23666] <= 32'b00000001010000000000001110010011;
ROM[23667] <= 32'b00000000010000111000001110010011;
ROM[23668] <= 32'b01000000011100010000001110110011;
ROM[23669] <= 32'b00000000011100000000001000110011;
ROM[23670] <= 32'b00000000001000000000000110110011;
ROM[23671] <= 32'b01010110000000010010000011101111;
ROM[23672] <= 32'b11111111110000010000000100010011;
ROM[23673] <= 32'b00000000000000010010001110000011;
ROM[23674] <= 32'b00000000011100011010000000100011;
ROM[23675] <= 32'b00000000000000011010001110000011;
ROM[23676] <= 32'b00000000011100010010000000100011;
ROM[23677] <= 32'b00000000010000010000000100010011;
ROM[23678] <= 32'b00000000000000100010001110000011;
ROM[23679] <= 32'b00000000011100010010000000100011;
ROM[23680] <= 32'b00000000010000010000000100010011;
ROM[23681] <= 32'b00000000000000010111001110110111;
ROM[23682] <= 32'b00100101000000111000001110010011;
ROM[23683] <= 32'b00000000111000111000001110110011;
ROM[23684] <= 32'b00000000011100010010000000100011;
ROM[23685] <= 32'b00000000010000010000000100010011;
ROM[23686] <= 32'b00000000001100010010000000100011;
ROM[23687] <= 32'b00000000010000010000000100010011;
ROM[23688] <= 32'b00000000010000010010000000100011;
ROM[23689] <= 32'b00000000010000010000000100010011;
ROM[23690] <= 32'b00000000010100010010000000100011;
ROM[23691] <= 32'b00000000010000010000000100010011;
ROM[23692] <= 32'b00000000011000010010000000100011;
ROM[23693] <= 32'b00000000010000010000000100010011;
ROM[23694] <= 32'b00000001010000000000001110010011;
ROM[23695] <= 32'b00000000100000111000001110010011;
ROM[23696] <= 32'b01000000011100010000001110110011;
ROM[23697] <= 32'b00000000011100000000001000110011;
ROM[23698] <= 32'b00000000001000000000000110110011;
ROM[23699] <= 32'b01000100010000010011000011101111;
ROM[23700] <= 32'b11111111110000010000000100010011;
ROM[23701] <= 32'b00000000000000010010001110000011;
ROM[23702] <= 32'b00000000011101100010000000100011;
ROM[23703] <= 32'b00000000000000011010001110000011;
ROM[23704] <= 32'b00000000011100010010000000100011;
ROM[23705] <= 32'b00000000010000010000000100010011;
ROM[23706] <= 32'b00000000000000010111001110110111;
ROM[23707] <= 32'b00101011010000111000001110010011;
ROM[23708] <= 32'b00000000111000111000001110110011;
ROM[23709] <= 32'b00000000011100010010000000100011;
ROM[23710] <= 32'b00000000010000010000000100010011;
ROM[23711] <= 32'b00000000001100010010000000100011;
ROM[23712] <= 32'b00000000010000010000000100010011;
ROM[23713] <= 32'b00000000010000010010000000100011;
ROM[23714] <= 32'b00000000010000010000000100010011;
ROM[23715] <= 32'b00000000010100010010000000100011;
ROM[23716] <= 32'b00000000010000010000000100010011;
ROM[23717] <= 32'b00000000011000010010000000100011;
ROM[23718] <= 32'b00000000010000010000000100010011;
ROM[23719] <= 32'b00000001010000000000001110010011;
ROM[23720] <= 32'b00000000010000111000001110010011;
ROM[23721] <= 32'b01000000011100010000001110110011;
ROM[23722] <= 32'b00000000011100000000001000110011;
ROM[23723] <= 32'b00000000001000000000000110110011;
ROM[23724] <= 32'b11001011100111111111000011101111;
ROM[23725] <= 32'b11111111110000010000000100010011;
ROM[23726] <= 32'b00000000000000010010001110000011;
ROM[23727] <= 32'b00000000011101100010000000100011;
ROM[23728] <= 32'b00000000000000011010001110000011;
ROM[23729] <= 32'b00000000011100010010000000100011;
ROM[23730] <= 32'b00000000010000010000000100010011;
ROM[23731] <= 32'b00000000000000010111001110110111;
ROM[23732] <= 32'b00110001100000111000001110010011;
ROM[23733] <= 32'b00000000111000111000001110110011;
ROM[23734] <= 32'b00000000011100010010000000100011;
ROM[23735] <= 32'b00000000010000010000000100010011;
ROM[23736] <= 32'b00000000001100010010000000100011;
ROM[23737] <= 32'b00000000010000010000000100010011;
ROM[23738] <= 32'b00000000010000010010000000100011;
ROM[23739] <= 32'b00000000010000010000000100010011;
ROM[23740] <= 32'b00000000010100010010000000100011;
ROM[23741] <= 32'b00000000010000010000000100010011;
ROM[23742] <= 32'b00000000011000010010000000100011;
ROM[23743] <= 32'b00000000010000010000000100010011;
ROM[23744] <= 32'b00000001010000000000001110010011;
ROM[23745] <= 32'b00000000010000111000001110010011;
ROM[23746] <= 32'b01000000011100010000001110110011;
ROM[23747] <= 32'b00000000011100000000001000110011;
ROM[23748] <= 32'b00000000001000000000000110110011;
ROM[23749] <= 32'b00011111110100010011000011101111;
ROM[23750] <= 32'b11111111110000010000000100010011;
ROM[23751] <= 32'b00000000000000010010001110000011;
ROM[23752] <= 32'b00000000011101100010000000100011;
ROM[23753] <= 32'b00000000000000000000001110010011;
ROM[23754] <= 32'b00000000011100010010000000100011;
ROM[23755] <= 32'b00000000010000010000000100010011;
ROM[23756] <= 32'b00000001010000000000001110010011;
ROM[23757] <= 32'b01000000011100011000001110110011;
ROM[23758] <= 32'b00000000000000111010000010000011;
ROM[23759] <= 32'b11111111110000010000000100010011;
ROM[23760] <= 32'b00000000000000010010001110000011;
ROM[23761] <= 32'b00000000011100100010000000100011;
ROM[23762] <= 32'b00000000010000100000000100010011;
ROM[23763] <= 32'b00000001010000000000001110010011;
ROM[23764] <= 32'b01000000011100011000001110110011;
ROM[23765] <= 32'b00000000010000111010000110000011;
ROM[23766] <= 32'b00000000100000111010001000000011;
ROM[23767] <= 32'b00000000110000111010001010000011;
ROM[23768] <= 32'b00000001000000111010001100000011;
ROM[23769] <= 32'b00000000000000001000000011100111;
ROM[23770] <= 32'b00001000010001101010001110000011;
ROM[23771] <= 32'b00000000011100010010000000100011;
ROM[23772] <= 32'b00000000010000010000000100010011;
ROM[23773] <= 32'b00000001110100000000001110010011;
ROM[23774] <= 32'b00000000011100010010000000100011;
ROM[23775] <= 32'b00000000010000010000000100010011;
ROM[23776] <= 32'b11111111110000010000000100010011;
ROM[23777] <= 32'b00000000000000010010001110000011;
ROM[23778] <= 32'b11111111110000010000000100010011;
ROM[23779] <= 32'b00000000000000010010010000000011;
ROM[23780] <= 32'b00000000011101000010001110110011;
ROM[23781] <= 32'b00000000011100010010000000100011;
ROM[23782] <= 32'b00000000010000010000000100010011;
ROM[23783] <= 32'b11111111110000010000000100010011;
ROM[23784] <= 32'b00000000000000010010001110000011;
ROM[23785] <= 32'b00000000000000111000101001100011;
ROM[23786] <= 32'b00000000000000010111001110110111;
ROM[23787] <= 32'b01000010110000111000001110010011;
ROM[23788] <= 32'b00000000111000111000001110110011;
ROM[23789] <= 32'b00000000000000111000000011100111;
ROM[23790] <= 32'b00000000000000000000001110010011;
ROM[23791] <= 32'b00000000011100010010000000100011;
ROM[23792] <= 32'b00000000010000010000000100010011;
ROM[23793] <= 32'b00000000000000000000001110010011;
ROM[23794] <= 32'b00000000011100010010000000100011;
ROM[23795] <= 32'b00000000010000010000000100010011;
ROM[23796] <= 32'b00000000000000010111001110110111;
ROM[23797] <= 32'b01000001110000111000001110010011;
ROM[23798] <= 32'b00000000111000111000001110110011;
ROM[23799] <= 32'b00000000011100010010000000100011;
ROM[23800] <= 32'b00000000010000010000000100010011;
ROM[23801] <= 32'b00000000001100010010000000100011;
ROM[23802] <= 32'b00000000010000010000000100010011;
ROM[23803] <= 32'b00000000010000010010000000100011;
ROM[23804] <= 32'b00000000010000010000000100010011;
ROM[23805] <= 32'b00000000010100010010000000100011;
ROM[23806] <= 32'b00000000010000010000000100010011;
ROM[23807] <= 32'b00000000011000010010000000100011;
ROM[23808] <= 32'b00000000010000010000000100010011;
ROM[23809] <= 32'b00000001010000000000001110010011;
ROM[23810] <= 32'b00000000100000111000001110010011;
ROM[23811] <= 32'b01000000011100010000001110110011;
ROM[23812] <= 32'b00000000011100000000001000110011;
ROM[23813] <= 32'b00000000001000000000000110110011;
ROM[23814] <= 32'b11111110100011111110000011101111;
ROM[23815] <= 32'b11111111110000010000000100010011;
ROM[23816] <= 32'b00000000000000010010001110000011;
ROM[23817] <= 32'b00000000011101100010000000100011;
ROM[23818] <= 32'b00001001110000000000000011101111;
ROM[23819] <= 32'b00001000010001101010001110000011;
ROM[23820] <= 32'b00000000011100010010000000100011;
ROM[23821] <= 32'b00000000010000010000000100010011;
ROM[23822] <= 32'b00000000000100000000001110010011;
ROM[23823] <= 32'b00000000011100010010000000100011;
ROM[23824] <= 32'b00000000010000010000000100010011;
ROM[23825] <= 32'b11111111110000010000000100010011;
ROM[23826] <= 32'b00000000000000010010001110000011;
ROM[23827] <= 32'b11111111110000010000000100010011;
ROM[23828] <= 32'b00000000000000010010010000000011;
ROM[23829] <= 32'b00000000011101000000001110110011;
ROM[23830] <= 32'b00000000011100010010000000100011;
ROM[23831] <= 32'b00000000010000010000000100010011;
ROM[23832] <= 32'b00000000000000000000001110010011;
ROM[23833] <= 32'b00000000011100010010000000100011;
ROM[23834] <= 32'b00000000010000010000000100010011;
ROM[23835] <= 32'b00000000000000010111001110110111;
ROM[23836] <= 32'b01001011100000111000001110010011;
ROM[23837] <= 32'b00000000111000111000001110110011;
ROM[23838] <= 32'b00000000011100010010000000100011;
ROM[23839] <= 32'b00000000010000010000000100010011;
ROM[23840] <= 32'b00000000001100010010000000100011;
ROM[23841] <= 32'b00000000010000010000000100010011;
ROM[23842] <= 32'b00000000010000010010000000100011;
ROM[23843] <= 32'b00000000010000010000000100010011;
ROM[23844] <= 32'b00000000010100010010000000100011;
ROM[23845] <= 32'b00000000010000010000000100010011;
ROM[23846] <= 32'b00000000011000010010000000100011;
ROM[23847] <= 32'b00000000010000010000000100010011;
ROM[23848] <= 32'b00000001010000000000001110010011;
ROM[23849] <= 32'b00000000100000111000001110010011;
ROM[23850] <= 32'b01000000011100010000001110110011;
ROM[23851] <= 32'b00000000011100000000001000110011;
ROM[23852] <= 32'b00000000001000000000000110110011;
ROM[23853] <= 32'b11110100110011111110000011101111;
ROM[23854] <= 32'b11111111110000010000000100010011;
ROM[23855] <= 32'b00000000000000010010001110000011;
ROM[23856] <= 32'b00000000011101100010000000100011;
ROM[23857] <= 32'b00000000000000000000001110010011;
ROM[23858] <= 32'b00000000011100010010000000100011;
ROM[23859] <= 32'b00000000010000010000000100010011;
ROM[23860] <= 32'b00000001010000000000001110010011;
ROM[23861] <= 32'b01000000011100011000001110110011;
ROM[23862] <= 32'b00000000000000111010000010000011;
ROM[23863] <= 32'b11111111110000010000000100010011;
ROM[23864] <= 32'b00000000000000010010001110000011;
ROM[23865] <= 32'b00000000011100100010000000100011;
ROM[23866] <= 32'b00000000010000100000000100010011;
ROM[23867] <= 32'b00000001010000000000001110010011;
ROM[23868] <= 32'b01000000011100011000001110110011;
ROM[23869] <= 32'b00000000010000111010000110000011;
ROM[23870] <= 32'b00000000100000111010001000000011;
ROM[23871] <= 32'b00000000110000111010001010000011;
ROM[23872] <= 32'b00000001000000111010001100000011;
ROM[23873] <= 32'b00000000000000001000000011100111;
ROM[23874] <= 32'b00000000000000010010000000100011;
ROM[23875] <= 32'b00000000010000010000000100010011;
ROM[23876] <= 32'b00000000000000010010000000100011;
ROM[23877] <= 32'b00000000010000010000000100010011;
ROM[23878] <= 32'b00000000000000010010000000100011;
ROM[23879] <= 32'b00000000010000010000000100010011;
ROM[23880] <= 32'b00000000000000010010000000100011;
ROM[23881] <= 32'b00000000010000010000000100010011;
ROM[23882] <= 32'b00000000000000010010000000100011;
ROM[23883] <= 32'b00000000010000010000000100010011;
ROM[23884] <= 32'b00000000000000010010000000100011;
ROM[23885] <= 32'b00000000010000010000000100010011;
ROM[23886] <= 32'b00000000000000010010000000100011;
ROM[23887] <= 32'b00000000010000010000000100010011;
ROM[23888] <= 32'b00000000000000010010000000100011;
ROM[23889] <= 32'b00000000010000010000000100010011;
ROM[23890] <= 32'b00000000000000010010000000100011;
ROM[23891] <= 32'b00000000010000010000000100010011;
ROM[23892] <= 32'b00001000000001101010001110000011;
ROM[23893] <= 32'b00000000011100010010000000100011;
ROM[23894] <= 32'b00000000010000010000000100010011;
ROM[23895] <= 32'b00000000000000000000001110010011;
ROM[23896] <= 32'b00000000011100010010000000100011;
ROM[23897] <= 32'b00000000010000010000000100010011;
ROM[23898] <= 32'b11111111110000010000000100010011;
ROM[23899] <= 32'b00000000000000010010001110000011;
ROM[23900] <= 32'b11111111110000010000000100010011;
ROM[23901] <= 32'b00000000000000010010010000000011;
ROM[23902] <= 32'b00000000011101000010010010110011;
ROM[23903] <= 32'b00000000100000111010010100110011;
ROM[23904] <= 32'b00000000101001001000001110110011;
ROM[23905] <= 32'b00000000000100111000001110010011;
ROM[23906] <= 32'b00000000000100111111001110010011;
ROM[23907] <= 32'b00000000011100010010000000100011;
ROM[23908] <= 32'b00000000010000010000000100010011;
ROM[23909] <= 32'b11111111110000010000000100010011;
ROM[23910] <= 32'b00000000000000010010001110000011;
ROM[23911] <= 32'b00000000000000111000101001100011;
ROM[23912] <= 32'b00000000000000010111001110110111;
ROM[23913] <= 32'b01100100110000111000001110010011;
ROM[23914] <= 32'b00000000111000111000001110110011;
ROM[23915] <= 32'b00000000000000111000000011100111;
ROM[23916] <= 32'b00001000010001101010001110000011;
ROM[23917] <= 32'b00000000011100010010000000100011;
ROM[23918] <= 32'b00000000010000010000000100010011;
ROM[23919] <= 32'b00001000000001101010001110000011;
ROM[23920] <= 32'b00000000011100010010000000100011;
ROM[23921] <= 32'b00000000010000010000000100010011;
ROM[23922] <= 32'b00000000000100000000001110010011;
ROM[23923] <= 32'b00000000011100010010000000100011;
ROM[23924] <= 32'b00000000010000010000000100010011;
ROM[23925] <= 32'b11111111110000010000000100010011;
ROM[23926] <= 32'b00000000000000010010001110000011;
ROM[23927] <= 32'b11111111110000010000000100010011;
ROM[23928] <= 32'b00000000000000010010010000000011;
ROM[23929] <= 32'b01000000011101000000001110110011;
ROM[23930] <= 32'b00000000011100010010000000100011;
ROM[23931] <= 32'b00000000010000010000000100010011;
ROM[23932] <= 32'b00000000000000010111001110110111;
ROM[23933] <= 32'b01100011110000111000001110010011;
ROM[23934] <= 32'b00000000111000111000001110110011;
ROM[23935] <= 32'b00000000011100010010000000100011;
ROM[23936] <= 32'b00000000010000010000000100010011;
ROM[23937] <= 32'b00000000001100010010000000100011;
ROM[23938] <= 32'b00000000010000010000000100010011;
ROM[23939] <= 32'b00000000010000010010000000100011;
ROM[23940] <= 32'b00000000010000010000000100010011;
ROM[23941] <= 32'b00000000010100010010000000100011;
ROM[23942] <= 32'b00000000010000010000000100010011;
ROM[23943] <= 32'b00000000011000010010000000100011;
ROM[23944] <= 32'b00000000010000010000000100010011;
ROM[23945] <= 32'b00000001010000000000001110010011;
ROM[23946] <= 32'b00000000100000111000001110010011;
ROM[23947] <= 32'b01000000011100010000001110110011;
ROM[23948] <= 32'b00000000011100000000001000110011;
ROM[23949] <= 32'b00000000001000000000000110110011;
ROM[23950] <= 32'b11011100100011111110000011101111;
ROM[23951] <= 32'b11111111110000010000000100010011;
ROM[23952] <= 32'b00000000000000010010001110000011;
ROM[23953] <= 32'b00000000011101100010000000100011;
ROM[23954] <= 32'b00010001100000000000000011101111;
ROM[23955] <= 32'b00001000010001101010001110000011;
ROM[23956] <= 32'b00000000011100010010000000100011;
ROM[23957] <= 32'b00000000010000010000000100010011;
ROM[23958] <= 32'b00000000000000000000001110010011;
ROM[23959] <= 32'b00000000011100010010000000100011;
ROM[23960] <= 32'b00000000010000010000000100010011;
ROM[23961] <= 32'b11111111110000010000000100010011;
ROM[23962] <= 32'b00000000000000010010001110000011;
ROM[23963] <= 32'b11111111110000010000000100010011;
ROM[23964] <= 32'b00000000000000010010010000000011;
ROM[23965] <= 32'b00000000011101000010010010110011;
ROM[23966] <= 32'b00000000100000111010010100110011;
ROM[23967] <= 32'b00000000101001001000001110110011;
ROM[23968] <= 32'b00000000000100111000001110010011;
ROM[23969] <= 32'b00000000000100111111001110010011;
ROM[23970] <= 32'b00000000011100010010000000100011;
ROM[23971] <= 32'b00000000010000010000000100010011;
ROM[23972] <= 32'b11111111110000010000000100010011;
ROM[23973] <= 32'b00000000000000010010001110000011;
ROM[23974] <= 32'b01000000011100000000001110110011;
ROM[23975] <= 32'b00000000000100111000001110010011;
ROM[23976] <= 32'b00000000011100010010000000100011;
ROM[23977] <= 32'b00000000010000010000000100010011;
ROM[23978] <= 32'b11111111110000010000000100010011;
ROM[23979] <= 32'b00000000000000010010001110000011;
ROM[23980] <= 32'b00000000000000111000101001100011;
ROM[23981] <= 32'b00000000000000010111001110110111;
ROM[23982] <= 32'b01101100100000111000001110010011;
ROM[23983] <= 32'b00000000111000111000001110110011;
ROM[23984] <= 32'b00000000000000111000000011100111;
ROM[23985] <= 32'b00001001110000000000000011101111;
ROM[23986] <= 32'b00001000010001101010001110000011;
ROM[23987] <= 32'b00000000011100010010000000100011;
ROM[23988] <= 32'b00000000010000010000000100010011;
ROM[23989] <= 32'b00000000000100000000001110010011;
ROM[23990] <= 32'b00000000011100010010000000100011;
ROM[23991] <= 32'b00000000010000010000000100010011;
ROM[23992] <= 32'b11111111110000010000000100010011;
ROM[23993] <= 32'b00000000000000010010001110000011;
ROM[23994] <= 32'b11111111110000010000000100010011;
ROM[23995] <= 32'b00000000000000010010010000000011;
ROM[23996] <= 32'b01000000011101000000001110110011;
ROM[23997] <= 32'b00000000011100010010000000100011;
ROM[23998] <= 32'b00000000010000010000000100010011;
ROM[23999] <= 32'b00000010011100000000001110010011;
ROM[24000] <= 32'b00000000011100010010000000100011;
ROM[24001] <= 32'b00000000010000010000000100010011;
ROM[24002] <= 32'b00000000000000010111001110110111;
ROM[24003] <= 32'b01110101010000111000001110010011;
ROM[24004] <= 32'b00000000111000111000001110110011;
ROM[24005] <= 32'b00000000011100010010000000100011;
ROM[24006] <= 32'b00000000010000010000000100010011;
ROM[24007] <= 32'b00000000001100010010000000100011;
ROM[24008] <= 32'b00000000010000010000000100010011;
ROM[24009] <= 32'b00000000010000010010000000100011;
ROM[24010] <= 32'b00000000010000010000000100010011;
ROM[24011] <= 32'b00000000010100010010000000100011;
ROM[24012] <= 32'b00000000010000010000000100010011;
ROM[24013] <= 32'b00000000011000010010000000100011;
ROM[24014] <= 32'b00000000010000010000000100010011;
ROM[24015] <= 32'b00000001010000000000001110010011;
ROM[24016] <= 32'b00000000100000111000001110010011;
ROM[24017] <= 32'b01000000011100010000001110110011;
ROM[24018] <= 32'b00000000011100000000001000110011;
ROM[24019] <= 32'b00000000001000000000000110110011;
ROM[24020] <= 32'b11001011000011111110000011101111;
ROM[24021] <= 32'b11111111110000010000000100010011;
ROM[24022] <= 32'b00000000000000010010001110000011;
ROM[24023] <= 32'b00000000011101100010000000100011;
ROM[24024] <= 32'b00001000010001101010001110000011;
ROM[24025] <= 32'b00000000011100010010000000100011;
ROM[24026] <= 32'b00000000010000010000000100010011;
ROM[24027] <= 32'b00000000101000000000001110010011;
ROM[24028] <= 32'b00000000011100010010000000100011;
ROM[24029] <= 32'b00000000010000010000000100010011;
ROM[24030] <= 32'b00000000000000010111001110110111;
ROM[24031] <= 32'b01111100010000111000001110010011;
ROM[24032] <= 32'b00000000111000111000001110110011;
ROM[24033] <= 32'b00000000011100010010000000100011;
ROM[24034] <= 32'b00000000010000010000000100010011;
ROM[24035] <= 32'b00000000001100010010000000100011;
ROM[24036] <= 32'b00000000010000010000000100010011;
ROM[24037] <= 32'b00000000010000010010000000100011;
ROM[24038] <= 32'b00000000010000010000000100010011;
ROM[24039] <= 32'b00000000010100010010000000100011;
ROM[24040] <= 32'b00000000010000010000000100010011;
ROM[24041] <= 32'b00000000011000010010000000100011;
ROM[24042] <= 32'b00000000010000010000000100010011;
ROM[24043] <= 32'b00000001010000000000001110010011;
ROM[24044] <= 32'b00000000100000111000001110010011;
ROM[24045] <= 32'b01000000011100010000001110110011;
ROM[24046] <= 32'b00000000011100000000001000110011;
ROM[24047] <= 32'b00000000001000000000000110110011;
ROM[24048] <= 32'b10000110110011111010000011101111;
ROM[24049] <= 32'b00000000100000000000001110010011;
ROM[24050] <= 32'b00000000011100010010000000100011;
ROM[24051] <= 32'b00000000010000010000000100010011;
ROM[24052] <= 32'b00000000000000011000001110110111;
ROM[24053] <= 32'b10000001110000111000001110010011;
ROM[24054] <= 32'b00000000111000111000001110110011;
ROM[24055] <= 32'b00000000011100010010000000100011;
ROM[24056] <= 32'b00000000010000010000000100010011;
ROM[24057] <= 32'b00000000001100010010000000100011;
ROM[24058] <= 32'b00000000010000010000000100010011;
ROM[24059] <= 32'b00000000010000010010000000100011;
ROM[24060] <= 32'b00000000010000010000000100010011;
ROM[24061] <= 32'b00000000010100010010000000100011;
ROM[24062] <= 32'b00000000010000010000000100010011;
ROM[24063] <= 32'b00000000011000010010000000100011;
ROM[24064] <= 32'b00000000010000010000000100010011;
ROM[24065] <= 32'b00000001010000000000001110010011;
ROM[24066] <= 32'b00000000100000111000001110010011;
ROM[24067] <= 32'b01000000011100010000001110110011;
ROM[24068] <= 32'b00000000011100000000001000110011;
ROM[24069] <= 32'b00000000001000000000000110110011;
ROM[24070] <= 32'b10000001010011111010000011101111;
ROM[24071] <= 32'b00001000000001101010001110000011;
ROM[24072] <= 32'b00000000011100010010000000100011;
ROM[24073] <= 32'b00000000010000010000000100010011;
ROM[24074] <= 32'b00000000010000000000001110010011;
ROM[24075] <= 32'b00000000011100010010000000100011;
ROM[24076] <= 32'b00000000010000010000000100010011;
ROM[24077] <= 32'b00000000000000011000001110110111;
ROM[24078] <= 32'b10001000000000111000001110010011;
ROM[24079] <= 32'b00000000111000111000001110110011;
ROM[24080] <= 32'b00000000011100010010000000100011;
ROM[24081] <= 32'b00000000010000010000000100010011;
ROM[24082] <= 32'b00000000001100010010000000100011;
ROM[24083] <= 32'b00000000010000010000000100010011;
ROM[24084] <= 32'b00000000010000010010000000100011;
ROM[24085] <= 32'b00000000010000010000000100010011;
ROM[24086] <= 32'b00000000010100010010000000100011;
ROM[24087] <= 32'b00000000010000010000000100010011;
ROM[24088] <= 32'b00000000011000010010000000100011;
ROM[24089] <= 32'b00000000010000010000000100010011;
ROM[24090] <= 32'b00000001010000000000001110010011;
ROM[24091] <= 32'b00000000100000111000001110010011;
ROM[24092] <= 32'b01000000011100010000001110110011;
ROM[24093] <= 32'b00000000011100000000001000110011;
ROM[24094] <= 32'b00000000001000000000000110110011;
ROM[24095] <= 32'b10110010110011111010000011101111;
ROM[24096] <= 32'b11111111110000010000000100010011;
ROM[24097] <= 32'b00000000000000010010001110000011;
ROM[24098] <= 32'b11111111110000010000000100010011;
ROM[24099] <= 32'b00000000000000010010010000000011;
ROM[24100] <= 32'b00000000011101000000001110110011;
ROM[24101] <= 32'b00000000011100010010000000100011;
ROM[24102] <= 32'b00000000010000010000000100010011;
ROM[24103] <= 32'b11111111110000010000000100010011;
ROM[24104] <= 32'b00000000000000010010001110000011;
ROM[24105] <= 32'b00000000011100011010000000100011;
ROM[24106] <= 32'b00001000000001101010001110000011;
ROM[24107] <= 32'b00000000011100010010000000100011;
ROM[24108] <= 32'b00000000010000010000000100010011;
ROM[24109] <= 32'b00000000001100000000001110010011;
ROM[24110] <= 32'b00000000011100010010000000100011;
ROM[24111] <= 32'b00000000010000010000000100010011;
ROM[24112] <= 32'b11111111110000010000000100010011;
ROM[24113] <= 32'b00000000000000010010001110000011;
ROM[24114] <= 32'b11111111110000010000000100010011;
ROM[24115] <= 32'b00000000000000010010010000000011;
ROM[24116] <= 32'b00000000011101000111001110110011;
ROM[24117] <= 32'b00000000011100010010000000100011;
ROM[24118] <= 32'b00000000010000010000000100010011;
ROM[24119] <= 32'b11111111110000010000000100010011;
ROM[24120] <= 32'b00000000000000010010001110000011;
ROM[24121] <= 32'b00000000011100011010010000100011;
ROM[24122] <= 32'b00000000000000000000001110010011;
ROM[24123] <= 32'b00000000011100010010000000100011;
ROM[24124] <= 32'b00000000010000010000000100010011;
ROM[24125] <= 32'b11111111110000010000000100010011;
ROM[24126] <= 32'b00000000000000010010001110000011;
ROM[24127] <= 32'b00000000011100011010001000100011;
ROM[24128] <= 32'b00000000010000011010001110000011;
ROM[24129] <= 32'b00000000011100010010000000100011;
ROM[24130] <= 32'b00000000010000010000000100010011;
ROM[24131] <= 32'b00000000100000000000001110010011;
ROM[24132] <= 32'b00000000011100010010000000100011;
ROM[24133] <= 32'b00000000010000010000000100010011;
ROM[24134] <= 32'b11111111110000010000000100010011;
ROM[24135] <= 32'b00000000000000010010001110000011;
ROM[24136] <= 32'b11111111110000010000000100010011;
ROM[24137] <= 32'b00000000000000010010010000000011;
ROM[24138] <= 32'b00000000011101000010001110110011;
ROM[24139] <= 32'b00000000011100010010000000100011;
ROM[24140] <= 32'b00000000010000010000000100010011;
ROM[24141] <= 32'b11111111110000010000000100010011;
ROM[24142] <= 32'b00000000000000010010001110000011;
ROM[24143] <= 32'b01000000011100000000001110110011;
ROM[24144] <= 32'b00000000000100111000001110010011;
ROM[24145] <= 32'b00000000011100010010000000100011;
ROM[24146] <= 32'b00000000010000010000000100010011;
ROM[24147] <= 32'b11111111110000010000000100010011;
ROM[24148] <= 32'b00000000000000010010001110000011;
ROM[24149] <= 32'b00000000000000111000101001100011;
ROM[24150] <= 32'b00000000000000011000001110110111;
ROM[24151] <= 32'b00111111100000111000001110010011;
ROM[24152] <= 32'b00000000111000111000001110110011;
ROM[24153] <= 32'b00000000000000111000000011100111;
ROM[24154] <= 32'b00000000010000011010001110000011;
ROM[24155] <= 32'b00000000011100010010000000100011;
ROM[24156] <= 32'b00000000010000010000000100010011;
ROM[24157] <= 32'b00000000010000000000001110010011;
ROM[24158] <= 32'b00000000011100010010000000100011;
ROM[24159] <= 32'b00000000010000010000000100010011;
ROM[24160] <= 32'b00000000000000011000001110110111;
ROM[24161] <= 32'b10011100110000111000001110010011;
ROM[24162] <= 32'b00000000111000111000001110110011;
ROM[24163] <= 32'b00000000011100010010000000100011;
ROM[24164] <= 32'b00000000010000010000000100010011;
ROM[24165] <= 32'b00000000001100010010000000100011;
ROM[24166] <= 32'b00000000010000010000000100010011;
ROM[24167] <= 32'b00000000010000010010000000100011;
ROM[24168] <= 32'b00000000010000010000000100010011;
ROM[24169] <= 32'b00000000010100010010000000100011;
ROM[24170] <= 32'b00000000010000010000000100010011;
ROM[24171] <= 32'b00000000011000010010000000100011;
ROM[24172] <= 32'b00000000010000010000000100010011;
ROM[24173] <= 32'b00000001010000000000001110010011;
ROM[24174] <= 32'b00000000100000111000001110010011;
ROM[24175] <= 32'b01000000011100010000001110110011;
ROM[24176] <= 32'b00000000011100000000001000110011;
ROM[24177] <= 32'b00000000001000000000000110110011;
ROM[24178] <= 32'b11100110010111111001000011101111;
ROM[24179] <= 32'b11111111110000010000000100010011;
ROM[24180] <= 32'b00000000000000010010001110000011;
ROM[24181] <= 32'b00000000011100011010011000100011;
ROM[24182] <= 32'b00000000000000011010001110000011;
ROM[24183] <= 32'b00000000011100010010000000100011;
ROM[24184] <= 32'b00000000010000010000000100010011;
ROM[24185] <= 32'b00000000010000000000001110010011;
ROM[24186] <= 32'b00000000011100010010000000100011;
ROM[24187] <= 32'b00000000010000010000000100010011;
ROM[24188] <= 32'b00000000000000011000001110110111;
ROM[24189] <= 32'b10100011110000111000001110010011;
ROM[24190] <= 32'b00000000111000111000001110110011;
ROM[24191] <= 32'b00000000011100010010000000100011;
ROM[24192] <= 32'b00000000010000010000000100010011;
ROM[24193] <= 32'b00000000001100010010000000100011;
ROM[24194] <= 32'b00000000010000010000000100010011;
ROM[24195] <= 32'b00000000010000010010000000100011;
ROM[24196] <= 32'b00000000010000010000000100010011;
ROM[24197] <= 32'b00000000010100010010000000100011;
ROM[24198] <= 32'b00000000010000010000000100010011;
ROM[24199] <= 32'b00000000011000010010000000100011;
ROM[24200] <= 32'b00000000010000010000000100010011;
ROM[24201] <= 32'b00000001010000000000001110010011;
ROM[24202] <= 32'b00000000100000111000001110010011;
ROM[24203] <= 32'b01000000011100010000001110110011;
ROM[24204] <= 32'b00000000011100000000001000110011;
ROM[24205] <= 32'b00000000001000000000000110110011;
ROM[24206] <= 32'b11011111010111111001000011101111;
ROM[24207] <= 32'b11111111110000010000000100010011;
ROM[24208] <= 32'b00000000000000010010001110000011;
ROM[24209] <= 32'b00000000011100011010100000100011;
ROM[24210] <= 32'b00000000100000011010001110000011;
ROM[24211] <= 32'b00000000011100010010000000100011;
ROM[24212] <= 32'b00000000010000010000000100010011;
ROM[24213] <= 32'b00000000000000000000001110010011;
ROM[24214] <= 32'b00000000011100010010000000100011;
ROM[24215] <= 32'b00000000010000010000000100010011;
ROM[24216] <= 32'b11111111110000010000000100010011;
ROM[24217] <= 32'b00000000000000010010001110000011;
ROM[24218] <= 32'b11111111110000010000000100010011;
ROM[24219] <= 32'b00000000000000010010010000000011;
ROM[24220] <= 32'b00000000011101000010010010110011;
ROM[24221] <= 32'b00000000100000111010010100110011;
ROM[24222] <= 32'b00000000101001001000001110110011;
ROM[24223] <= 32'b00000000000100111000001110010011;
ROM[24224] <= 32'b00000000000100111111001110010011;
ROM[24225] <= 32'b00000000011100010010000000100011;
ROM[24226] <= 32'b00000000010000010000000100010011;
ROM[24227] <= 32'b11111111110000010000000100010011;
ROM[24228] <= 32'b00000000000000010010001110000011;
ROM[24229] <= 32'b00000000000000111000101001100011;
ROM[24230] <= 32'b00000000000000011000001110110111;
ROM[24231] <= 32'b00011110110000111000001110010011;
ROM[24232] <= 32'b00000000111000111000001110110011;
ROM[24233] <= 32'b00000000000000111000000011100111;
ROM[24234] <= 32'b00000000100000011010001110000011;
ROM[24235] <= 32'b00000000011100010010000000100011;
ROM[24236] <= 32'b00000000010000010000000100010011;
ROM[24237] <= 32'b00000000000100000000001110010011;
ROM[24238] <= 32'b00000000011100010010000000100011;
ROM[24239] <= 32'b00000000010000010000000100010011;
ROM[24240] <= 32'b11111111110000010000000100010011;
ROM[24241] <= 32'b00000000000000010010001110000011;
ROM[24242] <= 32'b11111111110000010000000100010011;
ROM[24243] <= 32'b00000000000000010010010000000011;
ROM[24244] <= 32'b00000000011101000010010010110011;
ROM[24245] <= 32'b00000000100000111010010100110011;
ROM[24246] <= 32'b00000000101001001000001110110011;
ROM[24247] <= 32'b00000000000100111000001110010011;
ROM[24248] <= 32'b00000000000100111111001110010011;
ROM[24249] <= 32'b00000000011100010010000000100011;
ROM[24250] <= 32'b00000000010000010000000100010011;
ROM[24251] <= 32'b11111111110000010000000100010011;
ROM[24252] <= 32'b00000000000000010010001110000011;
ROM[24253] <= 32'b00000000000000111000101001100011;
ROM[24254] <= 32'b00000000000000011000001110110111;
ROM[24255] <= 32'b11110101010000111000001110010011;
ROM[24256] <= 32'b00000000111000111000001110110011;
ROM[24257] <= 32'b00000000000000111000000011100111;
ROM[24258] <= 32'b00000000100000011010001110000011;
ROM[24259] <= 32'b00000000011100010010000000100011;
ROM[24260] <= 32'b00000000010000010000000100010011;
ROM[24261] <= 32'b00000000001000000000001110010011;
ROM[24262] <= 32'b00000000011100010010000000100011;
ROM[24263] <= 32'b00000000010000010000000100010011;
ROM[24264] <= 32'b11111111110000010000000100010011;
ROM[24265] <= 32'b00000000000000010010001110000011;
ROM[24266] <= 32'b11111111110000010000000100010011;
ROM[24267] <= 32'b00000000000000010010010000000011;
ROM[24268] <= 32'b00000000011101000010010010110011;
ROM[24269] <= 32'b00000000100000111010010100110011;
ROM[24270] <= 32'b00000000101001001000001110110011;
ROM[24271] <= 32'b00000000000100111000001110010011;
ROM[24272] <= 32'b00000000000100111111001110010011;
ROM[24273] <= 32'b00000000011100010010000000100011;
ROM[24274] <= 32'b00000000010000010000000100010011;
ROM[24275] <= 32'b11111111110000010000000100010011;
ROM[24276] <= 32'b00000000000000010010001110000011;
ROM[24277] <= 32'b00000000000000111000101001100011;
ROM[24278] <= 32'b00000000000000011000001110110111;
ROM[24279] <= 32'b11001011110000111000001110010011;
ROM[24280] <= 32'b00000000111000111000001110110011;
ROM[24281] <= 32'b00000000000000111000000011100111;
ROM[24282] <= 32'b00000111110001101010001110000011;
ROM[24283] <= 32'b00000000011100010010000000100011;
ROM[24284] <= 32'b00000000010000010000000100010011;
ROM[24285] <= 32'b00000001000000011010001110000011;
ROM[24286] <= 32'b00000000011100010010000000100011;
ROM[24287] <= 32'b00000000010000010000000100010011;
ROM[24288] <= 32'b11111111110000010000000100010011;
ROM[24289] <= 32'b00000000000000010010001110000011;
ROM[24290] <= 32'b11111111110000010000000100010011;
ROM[24291] <= 32'b00000000000000010010010000000011;
ROM[24292] <= 32'b00000000011101000000001110110011;
ROM[24293] <= 32'b00000000011100010010000000100011;
ROM[24294] <= 32'b00000000010000010000000100010011;
ROM[24295] <= 32'b11111111110000010000000100010011;
ROM[24296] <= 32'b00000000000000010010001110000011;
ROM[24297] <= 32'b00000000000000111000001100010011;
ROM[24298] <= 32'b00000000110100110000010000110011;
ROM[24299] <= 32'b00000000000001000010001110000011;
ROM[24300] <= 32'b00000000011100010010000000100011;
ROM[24301] <= 32'b00000000010000010000000100010011;
ROM[24302] <= 32'b00010000000000000000001110010011;
ROM[24303] <= 32'b00000000011100010010000000100011;
ROM[24304] <= 32'b00000000010000010000000100010011;
ROM[24305] <= 32'b11111111110000010000000100010011;
ROM[24306] <= 32'b00000000000000010010001110000011;
ROM[24307] <= 32'b01000000011100000000001110110011;
ROM[24308] <= 32'b00000000011100010010000000100011;
ROM[24309] <= 32'b00000000010000010000000100010011;
ROM[24310] <= 32'b11111111110000010000000100010011;
ROM[24311] <= 32'b00000000000000010010001110000011;
ROM[24312] <= 32'b11111111110000010000000100010011;
ROM[24313] <= 32'b00000000000000010010010000000011;
ROM[24314] <= 32'b00000000011101000111001110110011;
ROM[24315] <= 32'b00000000011100010010000000100011;
ROM[24316] <= 32'b00000000010000010000000100010011;
ROM[24317] <= 32'b11111111110000010000000100010011;
ROM[24318] <= 32'b00000000000000010010001110000011;
ROM[24319] <= 32'b00000010011100011010000000100011;
ROM[24320] <= 32'b00000010000000011010001110000011;
ROM[24321] <= 32'b00000000011100010010000000100011;
ROM[24322] <= 32'b00000000010000010000000100010011;
ROM[24323] <= 32'b00000111100001101010001110000011;
ROM[24324] <= 32'b00000000011100010010000000100011;
ROM[24325] <= 32'b00000000010000010000000100010011;
ROM[24326] <= 32'b00000001000000011010001110000011;
ROM[24327] <= 32'b00000000011100010010000000100011;
ROM[24328] <= 32'b00000000010000010000000100010011;
ROM[24329] <= 32'b11111111110000010000000100010011;
ROM[24330] <= 32'b00000000000000010010001110000011;
ROM[24331] <= 32'b11111111110000010000000100010011;
ROM[24332] <= 32'b00000000000000010010010000000011;
ROM[24333] <= 32'b00000000011101000000001110110011;
ROM[24334] <= 32'b00000000011100010010000000100011;
ROM[24335] <= 32'b00000000010000010000000100010011;
ROM[24336] <= 32'b11111111110000010000000100010011;
ROM[24337] <= 32'b00000000000000010010001110000011;
ROM[24338] <= 32'b00000000000000111000001100010011;
ROM[24339] <= 32'b11111111110000010000000100010011;
ROM[24340] <= 32'b00000000000000010010001110000011;
ROM[24341] <= 32'b00000000110100110000010000110011;
ROM[24342] <= 32'b00000000011101000010000000100011;
ROM[24343] <= 32'b00000010000000011010001110000011;
ROM[24344] <= 32'b00000000011100010010000000100011;
ROM[24345] <= 32'b00000000010000010000000100010011;
ROM[24346] <= 32'b00000111110001101010001110000011;
ROM[24347] <= 32'b00000000011100010010000000100011;
ROM[24348] <= 32'b00000000010000010000000100010011;
ROM[24349] <= 32'b00000001000000011010001110000011;
ROM[24350] <= 32'b00000000011100010010000000100011;
ROM[24351] <= 32'b00000000010000010000000100010011;
ROM[24352] <= 32'b11111111110000010000000100010011;
ROM[24353] <= 32'b00000000000000010010001110000011;
ROM[24354] <= 32'b11111111110000010000000100010011;
ROM[24355] <= 32'b00000000000000010010010000000011;
ROM[24356] <= 32'b00000000011101000000001110110011;
ROM[24357] <= 32'b00000000011100010010000000100011;
ROM[24358] <= 32'b00000000010000010000000100010011;
ROM[24359] <= 32'b11111111110000010000000100010011;
ROM[24360] <= 32'b00000000000000010010001110000011;
ROM[24361] <= 32'b00000000000000111000001100010011;
ROM[24362] <= 32'b11111111110000010000000100010011;
ROM[24363] <= 32'b00000000000000010010001110000011;
ROM[24364] <= 32'b00000000110100110000010000110011;
ROM[24365] <= 32'b00000000011101000010000000100011;
ROM[24366] <= 32'b00101001100000000000000011101111;
ROM[24367] <= 32'b00000001000000000000001110010011;
ROM[24368] <= 32'b00000000011100010010000000100011;
ROM[24369] <= 32'b00000000010000010000000100010011;
ROM[24370] <= 32'b00000000000000011000001110110111;
ROM[24371] <= 32'b11010001010000111000001110010011;
ROM[24372] <= 32'b00000000111000111000001110110011;
ROM[24373] <= 32'b00000000011100010010000000100011;
ROM[24374] <= 32'b00000000010000010000000100010011;
ROM[24375] <= 32'b00000000001100010010000000100011;
ROM[24376] <= 32'b00000000010000010000000100010011;
ROM[24377] <= 32'b00000000010000010010000000100011;
ROM[24378] <= 32'b00000000010000010000000100010011;
ROM[24379] <= 32'b00000000010100010010000000100011;
ROM[24380] <= 32'b00000000010000010000000100010011;
ROM[24381] <= 32'b00000000011000010010000000100011;
ROM[24382] <= 32'b00000000010000010000000100010011;
ROM[24383] <= 32'b00000001010000000000001110010011;
ROM[24384] <= 32'b00000000010000111000001110010011;
ROM[24385] <= 32'b01000000011100010000001110110011;
ROM[24386] <= 32'b00000000011100000000001000110011;
ROM[24387] <= 32'b00000000001000000000000110110011;
ROM[24388] <= 32'b11000101110011111011000011101111;
ROM[24389] <= 32'b00000000100000000000001110010011;
ROM[24390] <= 32'b00000000011100010010000000100011;
ROM[24391] <= 32'b00000000010000010000000100010011;
ROM[24392] <= 32'b00000000000000011000001110110111;
ROM[24393] <= 32'b11010110110000111000001110010011;
ROM[24394] <= 32'b00000000111000111000001110110011;
ROM[24395] <= 32'b00000000011100010010000000100011;
ROM[24396] <= 32'b00000000010000010000000100010011;
ROM[24397] <= 32'b00000000001100010010000000100011;
ROM[24398] <= 32'b00000000010000010000000100010011;
ROM[24399] <= 32'b00000000010000010010000000100011;
ROM[24400] <= 32'b00000000010000010000000100010011;
ROM[24401] <= 32'b00000000010100010010000000100011;
ROM[24402] <= 32'b00000000010000010000000100010011;
ROM[24403] <= 32'b00000000011000010010000000100011;
ROM[24404] <= 32'b00000000010000010000000100010011;
ROM[24405] <= 32'b00000001010000000000001110010011;
ROM[24406] <= 32'b00000000010000111000001110010011;
ROM[24407] <= 32'b01000000011100010000001110110011;
ROM[24408] <= 32'b00000000011100000000001000110011;
ROM[24409] <= 32'b00000000001000000000000110110011;
ROM[24410] <= 32'b11000000010011111011000011101111;
ROM[24411] <= 32'b11111111110000010000000100010011;
ROM[24412] <= 32'b00000000000000010010001110000011;
ROM[24413] <= 32'b11111111110000010000000100010011;
ROM[24414] <= 32'b00000000000000010010010000000011;
ROM[24415] <= 32'b01000000011101000000001110110011;
ROM[24416] <= 32'b00000000011100010010000000100011;
ROM[24417] <= 32'b00000000010000010000000100010011;
ROM[24418] <= 32'b11111111110000010000000100010011;
ROM[24419] <= 32'b00000000000000010010001110000011;
ROM[24420] <= 32'b00000000011100011010110000100011;
ROM[24421] <= 32'b00000000000000000000001110010011;
ROM[24422] <= 32'b00000000011100010010000000100011;
ROM[24423] <= 32'b00000000010000010000000100010011;
ROM[24424] <= 32'b00000001100000011010001110000011;
ROM[24425] <= 32'b00000000011100010010000000100011;
ROM[24426] <= 32'b00000000010000010000000100010011;
ROM[24427] <= 32'b11111111110000010000000100010011;
ROM[24428] <= 32'b00000000000000010010001110000011;
ROM[24429] <= 32'b11111111110000010000000100010011;
ROM[24430] <= 32'b00000000000000010010010000000011;
ROM[24431] <= 32'b01000000011101000000001110110011;
ROM[24432] <= 32'b00000000011100010010000000100011;
ROM[24433] <= 32'b00000000010000010000000100010011;
ROM[24434] <= 32'b11111111110000010000000100010011;
ROM[24435] <= 32'b00000000000000010010001110000011;
ROM[24436] <= 32'b00000000011100011010111000100011;
ROM[24437] <= 32'b00000001110000011010001110000011;
ROM[24438] <= 32'b00000000011100010010000000100011;
ROM[24439] <= 32'b00000000010000010000000100010011;
ROM[24440] <= 32'b00000000000100000000001110010011;
ROM[24441] <= 32'b00000000011100010010000000100011;
ROM[24442] <= 32'b00000000010000010000000100010011;
ROM[24443] <= 32'b11111111110000010000000100010011;
ROM[24444] <= 32'b00000000000000010010001110000011;
ROM[24445] <= 32'b11111111110000010000000100010011;
ROM[24446] <= 32'b00000000000000010010010000000011;
ROM[24447] <= 32'b01000000011101000000001110110011;
ROM[24448] <= 32'b00000000011100010010000000100011;
ROM[24449] <= 32'b00000000010000010000000100010011;
ROM[24450] <= 32'b11111111110000010000000100010011;
ROM[24451] <= 32'b00000000000000010010001110000011;
ROM[24452] <= 32'b00000000011100011010111000100011;
ROM[24453] <= 32'b00000111110001101010001110000011;
ROM[24454] <= 32'b00000000011100010010000000100011;
ROM[24455] <= 32'b00000000010000010000000100010011;
ROM[24456] <= 32'b00000001000000011010001110000011;
ROM[24457] <= 32'b00000000011100010010000000100011;
ROM[24458] <= 32'b00000000010000010000000100010011;
ROM[24459] <= 32'b11111111110000010000000100010011;
ROM[24460] <= 32'b00000000000000010010001110000011;
ROM[24461] <= 32'b11111111110000010000000100010011;
ROM[24462] <= 32'b00000000000000010010010000000011;
ROM[24463] <= 32'b00000000011101000000001110110011;
ROM[24464] <= 32'b00000000011100010010000000100011;
ROM[24465] <= 32'b00000000010000010000000100010011;
ROM[24466] <= 32'b11111111110000010000000100010011;
ROM[24467] <= 32'b00000000000000010010001110000011;
ROM[24468] <= 32'b00000000000000111000001100010011;
ROM[24469] <= 32'b00000000110100110000010000110011;
ROM[24470] <= 32'b00000000000001000010001110000011;
ROM[24471] <= 32'b00000000011100010010000000100011;
ROM[24472] <= 32'b00000000010000010000000100010011;
ROM[24473] <= 32'b00000001110000011010001110000011;
ROM[24474] <= 32'b00000000011100010010000000100011;
ROM[24475] <= 32'b00000000010000010000000100010011;
ROM[24476] <= 32'b11111111110000010000000100010011;
ROM[24477] <= 32'b00000000000000010010001110000011;
ROM[24478] <= 32'b11111111110000010000000100010011;
ROM[24479] <= 32'b00000000000000010010010000000011;
ROM[24480] <= 32'b00000000011101000111001110110011;
ROM[24481] <= 32'b00000000011100010010000000100011;
ROM[24482] <= 32'b00000000010000010000000100010011;
ROM[24483] <= 32'b11111111110000010000000100010011;
ROM[24484] <= 32'b00000000000000010010001110000011;
ROM[24485] <= 32'b00000010011100011010000000100011;
ROM[24486] <= 32'b00000010000000011010001110000011;
ROM[24487] <= 32'b00000000011100010010000000100011;
ROM[24488] <= 32'b00000000010000010000000100010011;
ROM[24489] <= 32'b00000111100001101010001110000011;
ROM[24490] <= 32'b00000000011100010010000000100011;
ROM[24491] <= 32'b00000000010000010000000100010011;
ROM[24492] <= 32'b00000001000000011010001110000011;
ROM[24493] <= 32'b00000000011100010010000000100011;
ROM[24494] <= 32'b00000000010000010000000100010011;
ROM[24495] <= 32'b11111111110000010000000100010011;
ROM[24496] <= 32'b00000000000000010010001110000011;
ROM[24497] <= 32'b11111111110000010000000100010011;
ROM[24498] <= 32'b00000000000000010010010000000011;
ROM[24499] <= 32'b00000000011101000000001110110011;
ROM[24500] <= 32'b00000000011100010010000000100011;
ROM[24501] <= 32'b00000000010000010000000100010011;
ROM[24502] <= 32'b11111111110000010000000100010011;
ROM[24503] <= 32'b00000000000000010010001110000011;
ROM[24504] <= 32'b00000000000000111000001100010011;
ROM[24505] <= 32'b11111111110000010000000100010011;
ROM[24506] <= 32'b00000000000000010010001110000011;
ROM[24507] <= 32'b00000000110100110000010000110011;
ROM[24508] <= 32'b00000000011101000010000000100011;
ROM[24509] <= 32'b00000010000000011010001110000011;
ROM[24510] <= 32'b00000000011100010010000000100011;
ROM[24511] <= 32'b00000000010000010000000100010011;
ROM[24512] <= 32'b00000111110001101010001110000011;
ROM[24513] <= 32'b00000000011100010010000000100011;
ROM[24514] <= 32'b00000000010000010000000100010011;
ROM[24515] <= 32'b00000001000000011010001110000011;
ROM[24516] <= 32'b00000000011100010010000000100011;
ROM[24517] <= 32'b00000000010000010000000100010011;
ROM[24518] <= 32'b11111111110000010000000100010011;
ROM[24519] <= 32'b00000000000000010010001110000011;
ROM[24520] <= 32'b11111111110000010000000100010011;
ROM[24521] <= 32'b00000000000000010010010000000011;
ROM[24522] <= 32'b00000000011101000000001110110011;
ROM[24523] <= 32'b00000000011100010010000000100011;
ROM[24524] <= 32'b00000000010000010000000100010011;
ROM[24525] <= 32'b11111111110000010000000100010011;
ROM[24526] <= 32'b00000000000000010010001110000011;
ROM[24527] <= 32'b00000000000000111000001100010011;
ROM[24528] <= 32'b11111111110000010000000100010011;
ROM[24529] <= 32'b00000000000000010010001110000011;
ROM[24530] <= 32'b00000000110100110000010000110011;
ROM[24531] <= 32'b00000000011101000010000000100011;
ROM[24532] <= 32'b00101001100000000000000011101111;
ROM[24533] <= 32'b00000001100000000000001110010011;
ROM[24534] <= 32'b00000000011100010010000000100011;
ROM[24535] <= 32'b00000000010000010000000100010011;
ROM[24536] <= 32'b00000000000000011000001110110111;
ROM[24537] <= 32'b11111010110000111000001110010011;
ROM[24538] <= 32'b00000000111000111000001110110011;
ROM[24539] <= 32'b00000000011100010010000000100011;
ROM[24540] <= 32'b00000000010000010000000100010011;
ROM[24541] <= 32'b00000000001100010010000000100011;
ROM[24542] <= 32'b00000000010000010000000100010011;
ROM[24543] <= 32'b00000000010000010010000000100011;
ROM[24544] <= 32'b00000000010000010000000100010011;
ROM[24545] <= 32'b00000000010100010010000000100011;
ROM[24546] <= 32'b00000000010000010000000100010011;
ROM[24547] <= 32'b00000000011000010010000000100011;
ROM[24548] <= 32'b00000000010000010000000100010011;
ROM[24549] <= 32'b00000001010000000000001110010011;
ROM[24550] <= 32'b00000000010000111000001110010011;
ROM[24551] <= 32'b01000000011100010000001110110011;
ROM[24552] <= 32'b00000000011100000000001000110011;
ROM[24553] <= 32'b00000000001000000000000110110011;
ROM[24554] <= 32'b10011100010011111011000011101111;
ROM[24555] <= 32'b00000001000000000000001110010011;
ROM[24556] <= 32'b00000000011100010010000000100011;
ROM[24557] <= 32'b00000000010000010000000100010011;
ROM[24558] <= 32'b00000000000000011000001110110111;
ROM[24559] <= 32'b00000000010000111000001110010011;
ROM[24560] <= 32'b00000000111000111000001110110011;
ROM[24561] <= 32'b00000000011100010010000000100011;
ROM[24562] <= 32'b00000000010000010000000100010011;
ROM[24563] <= 32'b00000000001100010010000000100011;
ROM[24564] <= 32'b00000000010000010000000100010011;
ROM[24565] <= 32'b00000000010000010010000000100011;
ROM[24566] <= 32'b00000000010000010000000100010011;
ROM[24567] <= 32'b00000000010100010010000000100011;
ROM[24568] <= 32'b00000000010000010000000100010011;
ROM[24569] <= 32'b00000000011000010010000000100011;
ROM[24570] <= 32'b00000000010000010000000100010011;
ROM[24571] <= 32'b00000001010000000000001110010011;
ROM[24572] <= 32'b00000000010000111000001110010011;
ROM[24573] <= 32'b01000000011100010000001110110011;
ROM[24574] <= 32'b00000000011100000000001000110011;
ROM[24575] <= 32'b00000000001000000000000110110011;
ROM[24576] <= 32'b10010110110011111011000011101111;
ROM[24577] <= 32'b11111111110000010000000100010011;
ROM[24578] <= 32'b00000000000000010010001110000011;
ROM[24579] <= 32'b11111111110000010000000100010011;
ROM[24580] <= 32'b00000000000000010010010000000011;
ROM[24581] <= 32'b01000000011101000000001110110011;
ROM[24582] <= 32'b00000000011100010010000000100011;
ROM[24583] <= 32'b00000000010000010000000100010011;
ROM[24584] <= 32'b11111111110000010000000100010011;
ROM[24585] <= 32'b00000000000000010010001110000011;
ROM[24586] <= 32'b00000000011100011010101000100011;
ROM[24587] <= 32'b00000000000000000000001110010011;
ROM[24588] <= 32'b00000000011100010010000000100011;
ROM[24589] <= 32'b00000000010000010000000100010011;
ROM[24590] <= 32'b00000001010000011010001110000011;
ROM[24591] <= 32'b00000000011100010010000000100011;
ROM[24592] <= 32'b00000000010000010000000100010011;
ROM[24593] <= 32'b11111111110000010000000100010011;
ROM[24594] <= 32'b00000000000000010010001110000011;
ROM[24595] <= 32'b11111111110000010000000100010011;
ROM[24596] <= 32'b00000000000000010010010000000011;
ROM[24597] <= 32'b01000000011101000000001110110011;
ROM[24598] <= 32'b00000000011100010010000000100011;
ROM[24599] <= 32'b00000000010000010000000100010011;
ROM[24600] <= 32'b11111111110000010000000100010011;
ROM[24601] <= 32'b00000000000000010010001110000011;
ROM[24602] <= 32'b00000000011100011010111000100011;
ROM[24603] <= 32'b00000001110000011010001110000011;
ROM[24604] <= 32'b00000000011100010010000000100011;
ROM[24605] <= 32'b00000000010000010000000100010011;
ROM[24606] <= 32'b00000000000100000000001110010011;
ROM[24607] <= 32'b00000000011100010010000000100011;
ROM[24608] <= 32'b00000000010000010000000100010011;
ROM[24609] <= 32'b11111111110000010000000100010011;
ROM[24610] <= 32'b00000000000000010010001110000011;
ROM[24611] <= 32'b11111111110000010000000100010011;
ROM[24612] <= 32'b00000000000000010010010000000011;
ROM[24613] <= 32'b01000000011101000000001110110011;
ROM[24614] <= 32'b00000000011100010010000000100011;
ROM[24615] <= 32'b00000000010000010000000100010011;
ROM[24616] <= 32'b11111111110000010000000100010011;
ROM[24617] <= 32'b00000000000000010010001110000011;
ROM[24618] <= 32'b00000000011100011010111000100011;
ROM[24619] <= 32'b00000111110001101010001110000011;
ROM[24620] <= 32'b00000000011100010010000000100011;
ROM[24621] <= 32'b00000000010000010000000100010011;
ROM[24622] <= 32'b00000001000000011010001110000011;
ROM[24623] <= 32'b00000000011100010010000000100011;
ROM[24624] <= 32'b00000000010000010000000100010011;
ROM[24625] <= 32'b11111111110000010000000100010011;
ROM[24626] <= 32'b00000000000000010010001110000011;
ROM[24627] <= 32'b11111111110000010000000100010011;
ROM[24628] <= 32'b00000000000000010010010000000011;
ROM[24629] <= 32'b00000000011101000000001110110011;
ROM[24630] <= 32'b00000000011100010010000000100011;
ROM[24631] <= 32'b00000000010000010000000100010011;
ROM[24632] <= 32'b11111111110000010000000100010011;
ROM[24633] <= 32'b00000000000000010010001110000011;
ROM[24634] <= 32'b00000000000000111000001100010011;
ROM[24635] <= 32'b00000000110100110000010000110011;
ROM[24636] <= 32'b00000000000001000010001110000011;
ROM[24637] <= 32'b00000000011100010010000000100011;
ROM[24638] <= 32'b00000000010000010000000100010011;
ROM[24639] <= 32'b00000001110000011010001110000011;
ROM[24640] <= 32'b00000000011100010010000000100011;
ROM[24641] <= 32'b00000000010000010000000100010011;
ROM[24642] <= 32'b11111111110000010000000100010011;
ROM[24643] <= 32'b00000000000000010010001110000011;
ROM[24644] <= 32'b11111111110000010000000100010011;
ROM[24645] <= 32'b00000000000000010010010000000011;
ROM[24646] <= 32'b00000000011101000111001110110011;
ROM[24647] <= 32'b00000000011100010010000000100011;
ROM[24648] <= 32'b00000000010000010000000100010011;
ROM[24649] <= 32'b11111111110000010000000100010011;
ROM[24650] <= 32'b00000000000000010010001110000011;
ROM[24651] <= 32'b00000010011100011010000000100011;
ROM[24652] <= 32'b00000010000000011010001110000011;
ROM[24653] <= 32'b00000000011100010010000000100011;
ROM[24654] <= 32'b00000000010000010000000100010011;
ROM[24655] <= 32'b00000111100001101010001110000011;
ROM[24656] <= 32'b00000000011100010010000000100011;
ROM[24657] <= 32'b00000000010000010000000100010011;
ROM[24658] <= 32'b00000001000000011010001110000011;
ROM[24659] <= 32'b00000000011100010010000000100011;
ROM[24660] <= 32'b00000000010000010000000100010011;
ROM[24661] <= 32'b11111111110000010000000100010011;
ROM[24662] <= 32'b00000000000000010010001110000011;
ROM[24663] <= 32'b11111111110000010000000100010011;
ROM[24664] <= 32'b00000000000000010010010000000011;
ROM[24665] <= 32'b00000000011101000000001110110011;
ROM[24666] <= 32'b00000000011100010010000000100011;
ROM[24667] <= 32'b00000000010000010000000100010011;
ROM[24668] <= 32'b11111111110000010000000100010011;
ROM[24669] <= 32'b00000000000000010010001110000011;
ROM[24670] <= 32'b00000000000000111000001100010011;
ROM[24671] <= 32'b11111111110000010000000100010011;
ROM[24672] <= 32'b00000000000000010010001110000011;
ROM[24673] <= 32'b00000000110100110000010000110011;
ROM[24674] <= 32'b00000000011101000010000000100011;
ROM[24675] <= 32'b00000010000000011010001110000011;
ROM[24676] <= 32'b00000000011100010010000000100011;
ROM[24677] <= 32'b00000000010000010000000100010011;
ROM[24678] <= 32'b00000111110001101010001110000011;
ROM[24679] <= 32'b00000000011100010010000000100011;
ROM[24680] <= 32'b00000000010000010000000100010011;
ROM[24681] <= 32'b00000001000000011010001110000011;
ROM[24682] <= 32'b00000000011100010010000000100011;
ROM[24683] <= 32'b00000000010000010000000100010011;
ROM[24684] <= 32'b11111111110000010000000100010011;
ROM[24685] <= 32'b00000000000000010010001110000011;
ROM[24686] <= 32'b11111111110000010000000100010011;
ROM[24687] <= 32'b00000000000000010010010000000011;
ROM[24688] <= 32'b00000000011101000000001110110011;
ROM[24689] <= 32'b00000000011100010010000000100011;
ROM[24690] <= 32'b00000000010000010000000100010011;
ROM[24691] <= 32'b11111111110000010000000100010011;
ROM[24692] <= 32'b00000000000000010010001110000011;
ROM[24693] <= 32'b00000000000000111000001100010011;
ROM[24694] <= 32'b11111111110000010000000100010011;
ROM[24695] <= 32'b00000000000000010010001110000011;
ROM[24696] <= 32'b00000000110100110000010000110011;
ROM[24697] <= 32'b00000000011101000010000000100011;
ROM[24698] <= 32'b00011100110000000000000011101111;
ROM[24699] <= 32'b00000001100000000000001110010011;
ROM[24700] <= 32'b00000000011100010010000000100011;
ROM[24701] <= 32'b00000000010000010000000100010011;
ROM[24702] <= 32'b00000000000000011000001110110111;
ROM[24703] <= 32'b00100100010000111000001110010011;
ROM[24704] <= 32'b00000000111000111000001110110011;
ROM[24705] <= 32'b00000000011100010010000000100011;
ROM[24706] <= 32'b00000000010000010000000100010011;
ROM[24707] <= 32'b00000000001100010010000000100011;
ROM[24708] <= 32'b00000000010000010000000100010011;
ROM[24709] <= 32'b00000000010000010010000000100011;
ROM[24710] <= 32'b00000000010000010000000100010011;
ROM[24711] <= 32'b00000000010100010010000000100011;
ROM[24712] <= 32'b00000000010000010000000100010011;
ROM[24713] <= 32'b00000000011000010010000000100011;
ROM[24714] <= 32'b00000000010000010000000100010011;
ROM[24715] <= 32'b00000001010000000000001110010011;
ROM[24716] <= 32'b00000000010000111000001110010011;
ROM[24717] <= 32'b01000000011100010000001110110011;
ROM[24718] <= 32'b00000000011100000000001000110011;
ROM[24719] <= 32'b00000000001000000000000110110011;
ROM[24720] <= 32'b11110010110111111010000011101111;
ROM[24721] <= 32'b00000000000100000000001110010011;
ROM[24722] <= 32'b00000000011100010010000000100011;
ROM[24723] <= 32'b00000000010000010000000100010011;
ROM[24724] <= 32'b11111111110000010000000100010011;
ROM[24725] <= 32'b00000000000000010010001110000011;
ROM[24726] <= 32'b11111111110000010000000100010011;
ROM[24727] <= 32'b00000000000000010010010000000011;
ROM[24728] <= 32'b01000000011101000000001110110011;
ROM[24729] <= 32'b00000000011100010010000000100011;
ROM[24730] <= 32'b00000000010000010000000100010011;
ROM[24731] <= 32'b11111111110000010000000100010011;
ROM[24732] <= 32'b00000000000000010010001110000011;
ROM[24733] <= 32'b00000000011100011010111000100011;
ROM[24734] <= 32'b00000111110001101010001110000011;
ROM[24735] <= 32'b00000000011100010010000000100011;
ROM[24736] <= 32'b00000000010000010000000100010011;
ROM[24737] <= 32'b00000001000000011010001110000011;
ROM[24738] <= 32'b00000000011100010010000000100011;
ROM[24739] <= 32'b00000000010000010000000100010011;
ROM[24740] <= 32'b11111111110000010000000100010011;
ROM[24741] <= 32'b00000000000000010010001110000011;
ROM[24742] <= 32'b11111111110000010000000100010011;
ROM[24743] <= 32'b00000000000000010010010000000011;
ROM[24744] <= 32'b00000000011101000000001110110011;
ROM[24745] <= 32'b00000000011100010010000000100011;
ROM[24746] <= 32'b00000000010000010000000100010011;
ROM[24747] <= 32'b11111111110000010000000100010011;
ROM[24748] <= 32'b00000000000000010010001110000011;
ROM[24749] <= 32'b00000000000000111000001100010011;
ROM[24750] <= 32'b00000000110100110000010000110011;
ROM[24751] <= 32'b00000000000001000010001110000011;
ROM[24752] <= 32'b00000000011100010010000000100011;
ROM[24753] <= 32'b00000000010000010000000100010011;
ROM[24754] <= 32'b00000001110000011010001110000011;
ROM[24755] <= 32'b00000000011100010010000000100011;
ROM[24756] <= 32'b00000000010000010000000100010011;
ROM[24757] <= 32'b11111111110000010000000100010011;
ROM[24758] <= 32'b00000000000000010010001110000011;
ROM[24759] <= 32'b11111111110000010000000100010011;
ROM[24760] <= 32'b00000000000000010010010000000011;
ROM[24761] <= 32'b00000000011101000111001110110011;
ROM[24762] <= 32'b00000000011100010010000000100011;
ROM[24763] <= 32'b00000000010000010000000100010011;
ROM[24764] <= 32'b11111111110000010000000100010011;
ROM[24765] <= 32'b00000000000000010010001110000011;
ROM[24766] <= 32'b00000010011100011010000000100011;
ROM[24767] <= 32'b00000010000000011010001110000011;
ROM[24768] <= 32'b00000000011100010010000000100011;
ROM[24769] <= 32'b00000000010000010000000100010011;
ROM[24770] <= 32'b00000111100001101010001110000011;
ROM[24771] <= 32'b00000000011100010010000000100011;
ROM[24772] <= 32'b00000000010000010000000100010011;
ROM[24773] <= 32'b00000001000000011010001110000011;
ROM[24774] <= 32'b00000000011100010010000000100011;
ROM[24775] <= 32'b00000000010000010000000100010011;
ROM[24776] <= 32'b11111111110000010000000100010011;
ROM[24777] <= 32'b00000000000000010010001110000011;
ROM[24778] <= 32'b11111111110000010000000100010011;
ROM[24779] <= 32'b00000000000000010010010000000011;
ROM[24780] <= 32'b00000000011101000000001110110011;
ROM[24781] <= 32'b00000000011100010010000000100011;
ROM[24782] <= 32'b00000000010000010000000100010011;
ROM[24783] <= 32'b11111111110000010000000100010011;
ROM[24784] <= 32'b00000000000000010010001110000011;
ROM[24785] <= 32'b00000000000000111000001100010011;
ROM[24786] <= 32'b11111111110000010000000100010011;
ROM[24787] <= 32'b00000000000000010010001110000011;
ROM[24788] <= 32'b00000000110100110000010000110011;
ROM[24789] <= 32'b00000000011101000010000000100011;
ROM[24790] <= 32'b00000010000000011010001110000011;
ROM[24791] <= 32'b00000000011100010010000000100011;
ROM[24792] <= 32'b00000000010000010000000100010011;
ROM[24793] <= 32'b00000111110001101010001110000011;
ROM[24794] <= 32'b00000000011100010010000000100011;
ROM[24795] <= 32'b00000000010000010000000100010011;
ROM[24796] <= 32'b00000001000000011010001110000011;
ROM[24797] <= 32'b00000000011100010010000000100011;
ROM[24798] <= 32'b00000000010000010000000100010011;
ROM[24799] <= 32'b11111111110000010000000100010011;
ROM[24800] <= 32'b00000000000000010010001110000011;
ROM[24801] <= 32'b11111111110000010000000100010011;
ROM[24802] <= 32'b00000000000000010010010000000011;
ROM[24803] <= 32'b00000000011101000000001110110011;
ROM[24804] <= 32'b00000000011100010010000000100011;
ROM[24805] <= 32'b00000000010000010000000100010011;
ROM[24806] <= 32'b11111111110000010000000100010011;
ROM[24807] <= 32'b00000000000000010010001110000011;
ROM[24808] <= 32'b00000000000000111000001100010011;
ROM[24809] <= 32'b11111111110000010000000100010011;
ROM[24810] <= 32'b00000000000000010010001110000011;
ROM[24811] <= 32'b00000000110100110000010000110011;
ROM[24812] <= 32'b00000000011101000010000000100011;
ROM[24813] <= 32'b00000000010000011010001110000011;
ROM[24814] <= 32'b00000000011100010010000000100011;
ROM[24815] <= 32'b00000000010000010000000100010011;
ROM[24816] <= 32'b00000000000100000000001110010011;
ROM[24817] <= 32'b00000000011100010010000000100011;
ROM[24818] <= 32'b00000000010000010000000100010011;
ROM[24819] <= 32'b11111111110000010000000100010011;
ROM[24820] <= 32'b00000000000000010010001110000011;
ROM[24821] <= 32'b11111111110000010000000100010011;
ROM[24822] <= 32'b00000000000000010010010000000011;
ROM[24823] <= 32'b00000000011101000000001110110011;
ROM[24824] <= 32'b00000000011100010010000000100011;
ROM[24825] <= 32'b00000000010000010000000100010011;
ROM[24826] <= 32'b11111111110000010000000100010011;
ROM[24827] <= 32'b00000000000000010010001110000011;
ROM[24828] <= 32'b00000000011100011010001000100011;
ROM[24829] <= 32'b11010000110011111111000011101111;
ROM[24830] <= 32'b00000000000000000000001110010011;
ROM[24831] <= 32'b00000000011100010010000000100011;
ROM[24832] <= 32'b00000000010000010000000100010011;
ROM[24833] <= 32'b00000001010000000000001110010011;
ROM[24834] <= 32'b01000000011100011000001110110011;
ROM[24835] <= 32'b00000000000000111010000010000011;
ROM[24836] <= 32'b11111111110000010000000100010011;
ROM[24837] <= 32'b00000000000000010010001110000011;
ROM[24838] <= 32'b00000000011100100010000000100011;
ROM[24839] <= 32'b00000000010000100000000100010011;
ROM[24840] <= 32'b00000001010000000000001110010011;
ROM[24841] <= 32'b01000000011100011000001110110011;
ROM[24842] <= 32'b00000000010000111010000110000011;
ROM[24843] <= 32'b00000000100000111010001000000011;
ROM[24844] <= 32'b00000000110000111010001010000011;
ROM[24845] <= 32'b00000001000000111010001100000011;
ROM[24846] <= 32'b00000000000000001000000011100111;
ROM[24847] <= 32'b00000000000000010010000000100011;
ROM[24848] <= 32'b00000000010000010000000100010011;
ROM[24849] <= 32'b00000000000000010010000000100011;
ROM[24850] <= 32'b00000000010000010000000100010011;
ROM[24851] <= 32'b00000000000000010010000000100011;
ROM[24852] <= 32'b00000000010000010000000100010011;
ROM[24853] <= 32'b00000001110100000000001110010011;
ROM[24854] <= 32'b00000000011100010010000000100011;
ROM[24855] <= 32'b00000000010000010000000100010011;
ROM[24856] <= 32'b00000000000000011000001110110111;
ROM[24857] <= 32'b01001010110000111000001110010011;
ROM[24858] <= 32'b00000000111000111000001110110011;
ROM[24859] <= 32'b00000000011100010010000000100011;
ROM[24860] <= 32'b00000000010000010000000100010011;
ROM[24861] <= 32'b00000000001100010010000000100011;
ROM[24862] <= 32'b00000000010000010000000100010011;
ROM[24863] <= 32'b00000000010000010010000000100011;
ROM[24864] <= 32'b00000000010000010000000100010011;
ROM[24865] <= 32'b00000000010100010010000000100011;
ROM[24866] <= 32'b00000000010000010000000100010011;
ROM[24867] <= 32'b00000000011000010010000000100011;
ROM[24868] <= 32'b00000000010000010000000100010011;
ROM[24869] <= 32'b00000001010000000000001110010011;
ROM[24870] <= 32'b00000000010000111000001110010011;
ROM[24871] <= 32'b01000000011100010000001110110011;
ROM[24872] <= 32'b00000000011100000000001000110011;
ROM[24873] <= 32'b00000000001000000000000110110011;
ROM[24874] <= 32'b00101001010000010001000011101111;
ROM[24875] <= 32'b00000100010100000000001110010011;
ROM[24876] <= 32'b00000000011100010010000000100011;
ROM[24877] <= 32'b00000000010000010000000100010011;
ROM[24878] <= 32'b00000000000000011000001110110111;
ROM[24879] <= 32'b01010000010000111000001110010011;
ROM[24880] <= 32'b00000000111000111000001110110011;
ROM[24881] <= 32'b00000000011100010010000000100011;
ROM[24882] <= 32'b00000000010000010000000100010011;
ROM[24883] <= 32'b00000000001100010010000000100011;
ROM[24884] <= 32'b00000000010000010000000100010011;
ROM[24885] <= 32'b00000000010000010010000000100011;
ROM[24886] <= 32'b00000000010000010000000100010011;
ROM[24887] <= 32'b00000000010100010010000000100011;
ROM[24888] <= 32'b00000000010000010000000100010011;
ROM[24889] <= 32'b00000000011000010010000000100011;
ROM[24890] <= 32'b00000000010000010000000100010011;
ROM[24891] <= 32'b00000001010000000000001110010011;
ROM[24892] <= 32'b00000000100000111000001110010011;
ROM[24893] <= 32'b01000000011100010000001110110011;
ROM[24894] <= 32'b00000000011100000000001000110011;
ROM[24895] <= 32'b00000000001000000000000110110011;
ROM[24896] <= 32'b01101010110000010001000011101111;
ROM[24897] <= 32'b00000110111000000000001110010011;
ROM[24898] <= 32'b00000000011100010010000000100011;
ROM[24899] <= 32'b00000000010000010000000100010011;
ROM[24900] <= 32'b00000000000000011000001110110111;
ROM[24901] <= 32'b01010101110000111000001110010011;
ROM[24902] <= 32'b00000000111000111000001110110011;
ROM[24903] <= 32'b00000000011100010010000000100011;
ROM[24904] <= 32'b00000000010000010000000100010011;
ROM[24905] <= 32'b00000000001100010010000000100011;
ROM[24906] <= 32'b00000000010000010000000100010011;
ROM[24907] <= 32'b00000000010000010010000000100011;
ROM[24908] <= 32'b00000000010000010000000100010011;
ROM[24909] <= 32'b00000000010100010010000000100011;
ROM[24910] <= 32'b00000000010000010000000100010011;
ROM[24911] <= 32'b00000000011000010010000000100011;
ROM[24912] <= 32'b00000000010000010000000100010011;
ROM[24913] <= 32'b00000001010000000000001110010011;
ROM[24914] <= 32'b00000000100000111000001110010011;
ROM[24915] <= 32'b01000000011100010000001110110011;
ROM[24916] <= 32'b00000000011100000000001000110011;
ROM[24917] <= 32'b00000000001000000000000110110011;
ROM[24918] <= 32'b01100101010000010001000011101111;
ROM[24919] <= 32'b00000111010000000000001110010011;
ROM[24920] <= 32'b00000000011100010010000000100011;
ROM[24921] <= 32'b00000000010000010000000100010011;
ROM[24922] <= 32'b00000000000000011000001110110111;
ROM[24923] <= 32'b01011011010000111000001110010011;
ROM[24924] <= 32'b00000000111000111000001110110011;
ROM[24925] <= 32'b00000000011100010010000000100011;
ROM[24926] <= 32'b00000000010000010000000100010011;
ROM[24927] <= 32'b00000000001100010010000000100011;
ROM[24928] <= 32'b00000000010000010000000100010011;
ROM[24929] <= 32'b00000000010000010010000000100011;
ROM[24930] <= 32'b00000000010000010000000100010011;
ROM[24931] <= 32'b00000000010100010010000000100011;
ROM[24932] <= 32'b00000000010000010000000100010011;
ROM[24933] <= 32'b00000000011000010010000000100011;
ROM[24934] <= 32'b00000000010000010000000100010011;
ROM[24935] <= 32'b00000001010000000000001110010011;
ROM[24936] <= 32'b00000000100000111000001110010011;
ROM[24937] <= 32'b01000000011100010000001110110011;
ROM[24938] <= 32'b00000000011100000000001000110011;
ROM[24939] <= 32'b00000000001000000000000110110011;
ROM[24940] <= 32'b01011111110000010001000011101111;
ROM[24941] <= 32'b00000110010100000000001110010011;
ROM[24942] <= 32'b00000000011100010010000000100011;
ROM[24943] <= 32'b00000000010000010000000100010011;
ROM[24944] <= 32'b00000000000000011000001110110111;
ROM[24945] <= 32'b01100000110000111000001110010011;
ROM[24946] <= 32'b00000000111000111000001110110011;
ROM[24947] <= 32'b00000000011100010010000000100011;
ROM[24948] <= 32'b00000000010000010000000100010011;
ROM[24949] <= 32'b00000000001100010010000000100011;
ROM[24950] <= 32'b00000000010000010000000100010011;
ROM[24951] <= 32'b00000000010000010010000000100011;
ROM[24952] <= 32'b00000000010000010000000100010011;
ROM[24953] <= 32'b00000000010100010010000000100011;
ROM[24954] <= 32'b00000000010000010000000100010011;
ROM[24955] <= 32'b00000000011000010010000000100011;
ROM[24956] <= 32'b00000000010000010000000100010011;
ROM[24957] <= 32'b00000001010000000000001110010011;
ROM[24958] <= 32'b00000000100000111000001110010011;
ROM[24959] <= 32'b01000000011100010000001110110011;
ROM[24960] <= 32'b00000000011100000000001000110011;
ROM[24961] <= 32'b00000000001000000000000110110011;
ROM[24962] <= 32'b01011010010000010001000011101111;
ROM[24963] <= 32'b00000111001000000000001110010011;
ROM[24964] <= 32'b00000000011100010010000000100011;
ROM[24965] <= 32'b00000000010000010000000100010011;
ROM[24966] <= 32'b00000000000000011000001110110111;
ROM[24967] <= 32'b01100110010000111000001110010011;
ROM[24968] <= 32'b00000000111000111000001110110011;
ROM[24969] <= 32'b00000000011100010010000000100011;
ROM[24970] <= 32'b00000000010000010000000100010011;
ROM[24971] <= 32'b00000000001100010010000000100011;
ROM[24972] <= 32'b00000000010000010000000100010011;
ROM[24973] <= 32'b00000000010000010010000000100011;
ROM[24974] <= 32'b00000000010000010000000100010011;
ROM[24975] <= 32'b00000000010100010010000000100011;
ROM[24976] <= 32'b00000000010000010000000100010011;
ROM[24977] <= 32'b00000000011000010010000000100011;
ROM[24978] <= 32'b00000000010000010000000100010011;
ROM[24979] <= 32'b00000001010000000000001110010011;
ROM[24980] <= 32'b00000000100000111000001110010011;
ROM[24981] <= 32'b01000000011100010000001110110011;
ROM[24982] <= 32'b00000000011100000000001000110011;
ROM[24983] <= 32'b00000000001000000000000110110011;
ROM[24984] <= 32'b01010100110000010001000011101111;
ROM[24985] <= 32'b00000010000000000000001110010011;
ROM[24986] <= 32'b00000000011100010010000000100011;
ROM[24987] <= 32'b00000000010000010000000100010011;
ROM[24988] <= 32'b00000000000000011000001110110111;
ROM[24989] <= 32'b01101011110000111000001110010011;
ROM[24990] <= 32'b00000000111000111000001110110011;
ROM[24991] <= 32'b00000000011100010010000000100011;
ROM[24992] <= 32'b00000000010000010000000100010011;
ROM[24993] <= 32'b00000000001100010010000000100011;
ROM[24994] <= 32'b00000000010000010000000100010011;
ROM[24995] <= 32'b00000000010000010010000000100011;
ROM[24996] <= 32'b00000000010000010000000100010011;
ROM[24997] <= 32'b00000000010100010010000000100011;
ROM[24998] <= 32'b00000000010000010000000100010011;
ROM[24999] <= 32'b00000000011000010010000000100011;
ROM[25000] <= 32'b00000000010000010000000100010011;
ROM[25001] <= 32'b00000001010000000000001110010011;
ROM[25002] <= 32'b00000000100000111000001110010011;
ROM[25003] <= 32'b01000000011100010000001110110011;
ROM[25004] <= 32'b00000000011100000000001000110011;
ROM[25005] <= 32'b00000000001000000000000110110011;
ROM[25006] <= 32'b01001111010000010001000011101111;
ROM[25007] <= 32'b00000111010000000000001110010011;
ROM[25008] <= 32'b00000000011100010010000000100011;
ROM[25009] <= 32'b00000000010000010000000100010011;
ROM[25010] <= 32'b00000000000000011000001110110111;
ROM[25011] <= 32'b01110001010000111000001110010011;
ROM[25012] <= 32'b00000000111000111000001110110011;
ROM[25013] <= 32'b00000000011100010010000000100011;
ROM[25014] <= 32'b00000000010000010000000100010011;
ROM[25015] <= 32'b00000000001100010010000000100011;
ROM[25016] <= 32'b00000000010000010000000100010011;
ROM[25017] <= 32'b00000000010000010010000000100011;
ROM[25018] <= 32'b00000000010000010000000100010011;
ROM[25019] <= 32'b00000000010100010010000000100011;
ROM[25020] <= 32'b00000000010000010000000100010011;
ROM[25021] <= 32'b00000000011000010010000000100011;
ROM[25022] <= 32'b00000000010000010000000100010011;
ROM[25023] <= 32'b00000001010000000000001110010011;
ROM[25024] <= 32'b00000000100000111000001110010011;
ROM[25025] <= 32'b01000000011100010000001110110011;
ROM[25026] <= 32'b00000000011100000000001000110011;
ROM[25027] <= 32'b00000000001000000000000110110011;
ROM[25028] <= 32'b01001001110000010001000011101111;
ROM[25029] <= 32'b00000110100000000000001110010011;
ROM[25030] <= 32'b00000000011100010010000000100011;
ROM[25031] <= 32'b00000000010000010000000100010011;
ROM[25032] <= 32'b00000000000000011000001110110111;
ROM[25033] <= 32'b01110110110000111000001110010011;
ROM[25034] <= 32'b00000000111000111000001110110011;
ROM[25035] <= 32'b00000000011100010010000000100011;
ROM[25036] <= 32'b00000000010000010000000100010011;
ROM[25037] <= 32'b00000000001100010010000000100011;
ROM[25038] <= 32'b00000000010000010000000100010011;
ROM[25039] <= 32'b00000000010000010010000000100011;
ROM[25040] <= 32'b00000000010000010000000100010011;
ROM[25041] <= 32'b00000000010100010010000000100011;
ROM[25042] <= 32'b00000000010000010000000100010011;
ROM[25043] <= 32'b00000000011000010010000000100011;
ROM[25044] <= 32'b00000000010000010000000100010011;
ROM[25045] <= 32'b00000001010000000000001110010011;
ROM[25046] <= 32'b00000000100000111000001110010011;
ROM[25047] <= 32'b01000000011100010000001110110011;
ROM[25048] <= 32'b00000000011100000000001000110011;
ROM[25049] <= 32'b00000000001000000000000110110011;
ROM[25050] <= 32'b01000100010000010001000011101111;
ROM[25051] <= 32'b00000110010100000000001110010011;
ROM[25052] <= 32'b00000000011100010010000000100011;
ROM[25053] <= 32'b00000000010000010000000100010011;
ROM[25054] <= 32'b00000000000000011000001110110111;
ROM[25055] <= 32'b01111100010000111000001110010011;
ROM[25056] <= 32'b00000000111000111000001110110011;
ROM[25057] <= 32'b00000000011100010010000000100011;
ROM[25058] <= 32'b00000000010000010000000100010011;
ROM[25059] <= 32'b00000000001100010010000000100011;
ROM[25060] <= 32'b00000000010000010000000100010011;
ROM[25061] <= 32'b00000000010000010010000000100011;
ROM[25062] <= 32'b00000000010000010000000100010011;
ROM[25063] <= 32'b00000000010100010010000000100011;
ROM[25064] <= 32'b00000000010000010000000100010011;
ROM[25065] <= 32'b00000000011000010010000000100011;
ROM[25066] <= 32'b00000000010000010000000100010011;
ROM[25067] <= 32'b00000001010000000000001110010011;
ROM[25068] <= 32'b00000000100000111000001110010011;
ROM[25069] <= 32'b01000000011100010000001110110011;
ROM[25070] <= 32'b00000000011100000000001000110011;
ROM[25071] <= 32'b00000000001000000000000110110011;
ROM[25072] <= 32'b00111110110000010001000011101111;
ROM[25073] <= 32'b00000010000000000000001110010011;
ROM[25074] <= 32'b00000000011100010010000000100011;
ROM[25075] <= 32'b00000000010000010000000100010011;
ROM[25076] <= 32'b00000000000000011001001110110111;
ROM[25077] <= 32'b10000001110000111000001110010011;
ROM[25078] <= 32'b00000000111000111000001110110011;
ROM[25079] <= 32'b00000000011100010010000000100011;
ROM[25080] <= 32'b00000000010000010000000100010011;
ROM[25081] <= 32'b00000000001100010010000000100011;
ROM[25082] <= 32'b00000000010000010000000100010011;
ROM[25083] <= 32'b00000000010000010010000000100011;
ROM[25084] <= 32'b00000000010000010000000100010011;
ROM[25085] <= 32'b00000000010100010010000000100011;
ROM[25086] <= 32'b00000000010000010000000100010011;
ROM[25087] <= 32'b00000000011000010010000000100011;
ROM[25088] <= 32'b00000000010000010000000100010011;
ROM[25089] <= 32'b00000001010000000000001110010011;
ROM[25090] <= 32'b00000000100000111000001110010011;
ROM[25091] <= 32'b01000000011100010000001110110011;
ROM[25092] <= 32'b00000000011100000000001000110011;
ROM[25093] <= 32'b00000000001000000000000110110011;
ROM[25094] <= 32'b00111001010000010001000011101111;
ROM[25095] <= 32'b00000111001100000000001110010011;
ROM[25096] <= 32'b00000000011100010010000000100011;
ROM[25097] <= 32'b00000000010000010000000100010011;
ROM[25098] <= 32'b00000000000000011001001110110111;
ROM[25099] <= 32'b10000111010000111000001110010011;
ROM[25100] <= 32'b00000000111000111000001110110011;
ROM[25101] <= 32'b00000000011100010010000000100011;
ROM[25102] <= 32'b00000000010000010000000100010011;
ROM[25103] <= 32'b00000000001100010010000000100011;
ROM[25104] <= 32'b00000000010000010000000100010011;
ROM[25105] <= 32'b00000000010000010010000000100011;
ROM[25106] <= 32'b00000000010000010000000100010011;
ROM[25107] <= 32'b00000000010100010010000000100011;
ROM[25108] <= 32'b00000000010000010000000100010011;
ROM[25109] <= 32'b00000000011000010010000000100011;
ROM[25110] <= 32'b00000000010000010000000100010011;
ROM[25111] <= 32'b00000001010000000000001110010011;
ROM[25112] <= 32'b00000000100000111000001110010011;
ROM[25113] <= 32'b01000000011100010000001110110011;
ROM[25114] <= 32'b00000000011100000000001000110011;
ROM[25115] <= 32'b00000000001000000000000110110011;
ROM[25116] <= 32'b00110011110000010001000011101111;
ROM[25117] <= 32'b00000110100100000000001110010011;
ROM[25118] <= 32'b00000000011100010010000000100011;
ROM[25119] <= 32'b00000000010000010000000100010011;
ROM[25120] <= 32'b00000000000000011001001110110111;
ROM[25121] <= 32'b10001100110000111000001110010011;
ROM[25122] <= 32'b00000000111000111000001110110011;
ROM[25123] <= 32'b00000000011100010010000000100011;
ROM[25124] <= 32'b00000000010000010000000100010011;
ROM[25125] <= 32'b00000000001100010010000000100011;
ROM[25126] <= 32'b00000000010000010000000100010011;
ROM[25127] <= 32'b00000000010000010010000000100011;
ROM[25128] <= 32'b00000000010000010000000100010011;
ROM[25129] <= 32'b00000000010100010010000000100011;
ROM[25130] <= 32'b00000000010000010000000100010011;
ROM[25131] <= 32'b00000000011000010010000000100011;
ROM[25132] <= 32'b00000000010000010000000100010011;
ROM[25133] <= 32'b00000001010000000000001110010011;
ROM[25134] <= 32'b00000000100000111000001110010011;
ROM[25135] <= 32'b01000000011100010000001110110011;
ROM[25136] <= 32'b00000000011100000000001000110011;
ROM[25137] <= 32'b00000000001000000000000110110011;
ROM[25138] <= 32'b00101110010000010001000011101111;
ROM[25139] <= 32'b00000111101000000000001110010011;
ROM[25140] <= 32'b00000000011100010010000000100011;
ROM[25141] <= 32'b00000000010000010000000100010011;
ROM[25142] <= 32'b00000000000000011001001110110111;
ROM[25143] <= 32'b10010010010000111000001110010011;
ROM[25144] <= 32'b00000000111000111000001110110011;
ROM[25145] <= 32'b00000000011100010010000000100011;
ROM[25146] <= 32'b00000000010000010000000100010011;
ROM[25147] <= 32'b00000000001100010010000000100011;
ROM[25148] <= 32'b00000000010000010000000100010011;
ROM[25149] <= 32'b00000000010000010010000000100011;
ROM[25150] <= 32'b00000000010000010000000100010011;
ROM[25151] <= 32'b00000000010100010010000000100011;
ROM[25152] <= 32'b00000000010000010000000100010011;
ROM[25153] <= 32'b00000000011000010010000000100011;
ROM[25154] <= 32'b00000000010000010000000100010011;
ROM[25155] <= 32'b00000001010000000000001110010011;
ROM[25156] <= 32'b00000000100000111000001110010011;
ROM[25157] <= 32'b01000000011100010000001110110011;
ROM[25158] <= 32'b00000000011100000000001000110011;
ROM[25159] <= 32'b00000000001000000000000110110011;
ROM[25160] <= 32'b00101000110000010001000011101111;
ROM[25161] <= 32'b00000110010100000000001110010011;
ROM[25162] <= 32'b00000000011100010010000000100011;
ROM[25163] <= 32'b00000000010000010000000100010011;
ROM[25164] <= 32'b00000000000000011001001110110111;
ROM[25165] <= 32'b10010111110000111000001110010011;
ROM[25166] <= 32'b00000000111000111000001110110011;
ROM[25167] <= 32'b00000000011100010010000000100011;
ROM[25168] <= 32'b00000000010000010000000100010011;
ROM[25169] <= 32'b00000000001100010010000000100011;
ROM[25170] <= 32'b00000000010000010000000100010011;
ROM[25171] <= 32'b00000000010000010010000000100011;
ROM[25172] <= 32'b00000000010000010000000100010011;
ROM[25173] <= 32'b00000000010100010010000000100011;
ROM[25174] <= 32'b00000000010000010000000100010011;
ROM[25175] <= 32'b00000000011000010010000000100011;
ROM[25176] <= 32'b00000000010000010000000100010011;
ROM[25177] <= 32'b00000001010000000000001110010011;
ROM[25178] <= 32'b00000000100000111000001110010011;
ROM[25179] <= 32'b01000000011100010000001110110011;
ROM[25180] <= 32'b00000000011100000000001000110011;
ROM[25181] <= 32'b00000000001000000000000110110011;
ROM[25182] <= 32'b00100011010000010001000011101111;
ROM[25183] <= 32'b00000010000000000000001110010011;
ROM[25184] <= 32'b00000000011100010010000000100011;
ROM[25185] <= 32'b00000000010000010000000100010011;
ROM[25186] <= 32'b00000000000000011001001110110111;
ROM[25187] <= 32'b10011101010000111000001110010011;
ROM[25188] <= 32'b00000000111000111000001110110011;
ROM[25189] <= 32'b00000000011100010010000000100011;
ROM[25190] <= 32'b00000000010000010000000100010011;
ROM[25191] <= 32'b00000000001100010010000000100011;
ROM[25192] <= 32'b00000000010000010000000100010011;
ROM[25193] <= 32'b00000000010000010010000000100011;
ROM[25194] <= 32'b00000000010000010000000100010011;
ROM[25195] <= 32'b00000000010100010010000000100011;
ROM[25196] <= 32'b00000000010000010000000100010011;
ROM[25197] <= 32'b00000000011000010010000000100011;
ROM[25198] <= 32'b00000000010000010000000100010011;
ROM[25199] <= 32'b00000001010000000000001110010011;
ROM[25200] <= 32'b00000000100000111000001110010011;
ROM[25201] <= 32'b01000000011100010000001110110011;
ROM[25202] <= 32'b00000000011100000000001000110011;
ROM[25203] <= 32'b00000000001000000000000110110011;
ROM[25204] <= 32'b00011101110000010001000011101111;
ROM[25205] <= 32'b00000110111100000000001110010011;
ROM[25206] <= 32'b00000000011100010010000000100011;
ROM[25207] <= 32'b00000000010000010000000100010011;
ROM[25208] <= 32'b00000000000000011001001110110111;
ROM[25209] <= 32'b10100010110000111000001110010011;
ROM[25210] <= 32'b00000000111000111000001110110011;
ROM[25211] <= 32'b00000000011100010010000000100011;
ROM[25212] <= 32'b00000000010000010000000100010011;
ROM[25213] <= 32'b00000000001100010010000000100011;
ROM[25214] <= 32'b00000000010000010000000100010011;
ROM[25215] <= 32'b00000000010000010010000000100011;
ROM[25216] <= 32'b00000000010000010000000100010011;
ROM[25217] <= 32'b00000000010100010010000000100011;
ROM[25218] <= 32'b00000000010000010000000100010011;
ROM[25219] <= 32'b00000000011000010010000000100011;
ROM[25220] <= 32'b00000000010000010000000100010011;
ROM[25221] <= 32'b00000001010000000000001110010011;
ROM[25222] <= 32'b00000000100000111000001110010011;
ROM[25223] <= 32'b01000000011100010000001110110011;
ROM[25224] <= 32'b00000000011100000000001000110011;
ROM[25225] <= 32'b00000000001000000000000110110011;
ROM[25226] <= 32'b00011000010000010001000011101111;
ROM[25227] <= 32'b00000110011000000000001110010011;
ROM[25228] <= 32'b00000000011100010010000000100011;
ROM[25229] <= 32'b00000000010000010000000100010011;
ROM[25230] <= 32'b00000000000000011001001110110111;
ROM[25231] <= 32'b10101000010000111000001110010011;
ROM[25232] <= 32'b00000000111000111000001110110011;
ROM[25233] <= 32'b00000000011100010010000000100011;
ROM[25234] <= 32'b00000000010000010000000100010011;
ROM[25235] <= 32'b00000000001100010010000000100011;
ROM[25236] <= 32'b00000000010000010000000100010011;
ROM[25237] <= 32'b00000000010000010010000000100011;
ROM[25238] <= 32'b00000000010000010000000100010011;
ROM[25239] <= 32'b00000000010100010010000000100011;
ROM[25240] <= 32'b00000000010000010000000100010011;
ROM[25241] <= 32'b00000000011000010010000000100011;
ROM[25242] <= 32'b00000000010000010000000100010011;
ROM[25243] <= 32'b00000001010000000000001110010011;
ROM[25244] <= 32'b00000000100000111000001110010011;
ROM[25245] <= 32'b01000000011100010000001110110011;
ROM[25246] <= 32'b00000000011100000000001000110011;
ROM[25247] <= 32'b00000000001000000000000110110011;
ROM[25248] <= 32'b00010010110000010001000011101111;
ROM[25249] <= 32'b00000010000000000000001110010011;
ROM[25250] <= 32'b00000000011100010010000000100011;
ROM[25251] <= 32'b00000000010000010000000100010011;
ROM[25252] <= 32'b00000000000000011001001110110111;
ROM[25253] <= 32'b10101101110000111000001110010011;
ROM[25254] <= 32'b00000000111000111000001110110011;
ROM[25255] <= 32'b00000000011100010010000000100011;
ROM[25256] <= 32'b00000000010000010000000100010011;
ROM[25257] <= 32'b00000000001100010010000000100011;
ROM[25258] <= 32'b00000000010000010000000100010011;
ROM[25259] <= 32'b00000000010000010010000000100011;
ROM[25260] <= 32'b00000000010000010000000100010011;
ROM[25261] <= 32'b00000000010100010010000000100011;
ROM[25262] <= 32'b00000000010000010000000100010011;
ROM[25263] <= 32'b00000000011000010010000000100011;
ROM[25264] <= 32'b00000000010000010000000100010011;
ROM[25265] <= 32'b00000001010000000000001110010011;
ROM[25266] <= 32'b00000000100000111000001110010011;
ROM[25267] <= 32'b01000000011100010000001110110011;
ROM[25268] <= 32'b00000000011100000000001000110011;
ROM[25269] <= 32'b00000000001000000000000110110011;
ROM[25270] <= 32'b00001101010000010001000011101111;
ROM[25271] <= 32'b00000111010000000000001110010011;
ROM[25272] <= 32'b00000000011100010010000000100011;
ROM[25273] <= 32'b00000000010000010000000100010011;
ROM[25274] <= 32'b00000000000000011001001110110111;
ROM[25275] <= 32'b10110011010000111000001110010011;
ROM[25276] <= 32'b00000000111000111000001110110011;
ROM[25277] <= 32'b00000000011100010010000000100011;
ROM[25278] <= 32'b00000000010000010000000100010011;
ROM[25279] <= 32'b00000000001100010010000000100011;
ROM[25280] <= 32'b00000000010000010000000100010011;
ROM[25281] <= 32'b00000000010000010010000000100011;
ROM[25282] <= 32'b00000000010000010000000100010011;
ROM[25283] <= 32'b00000000010100010010000000100011;
ROM[25284] <= 32'b00000000010000010000000100010011;
ROM[25285] <= 32'b00000000011000010010000000100011;
ROM[25286] <= 32'b00000000010000010000000100010011;
ROM[25287] <= 32'b00000001010000000000001110010011;
ROM[25288] <= 32'b00000000100000111000001110010011;
ROM[25289] <= 32'b01000000011100010000001110110011;
ROM[25290] <= 32'b00000000011100000000001000110011;
ROM[25291] <= 32'b00000000001000000000000110110011;
ROM[25292] <= 32'b00000111110000010001000011101111;
ROM[25293] <= 32'b00000110100000000000001110010011;
ROM[25294] <= 32'b00000000011100010010000000100011;
ROM[25295] <= 32'b00000000010000010000000100010011;
ROM[25296] <= 32'b00000000000000011001001110110111;
ROM[25297] <= 32'b10111000110000111000001110010011;
ROM[25298] <= 32'b00000000111000111000001110110011;
ROM[25299] <= 32'b00000000011100010010000000100011;
ROM[25300] <= 32'b00000000010000010000000100010011;
ROM[25301] <= 32'b00000000001100010010000000100011;
ROM[25302] <= 32'b00000000010000010000000100010011;
ROM[25303] <= 32'b00000000010000010010000000100011;
ROM[25304] <= 32'b00000000010000010000000100010011;
ROM[25305] <= 32'b00000000010100010010000000100011;
ROM[25306] <= 32'b00000000010000010000000100010011;
ROM[25307] <= 32'b00000000011000010010000000100011;
ROM[25308] <= 32'b00000000010000010000000100010011;
ROM[25309] <= 32'b00000001010000000000001110010011;
ROM[25310] <= 32'b00000000100000111000001110010011;
ROM[25311] <= 32'b01000000011100010000001110110011;
ROM[25312] <= 32'b00000000011100000000001000110011;
ROM[25313] <= 32'b00000000001000000000000110110011;
ROM[25314] <= 32'b00000010010000010001000011101111;
ROM[25315] <= 32'b00000110010100000000001110010011;
ROM[25316] <= 32'b00000000011100010010000000100011;
ROM[25317] <= 32'b00000000010000010000000100010011;
ROM[25318] <= 32'b00000000000000011001001110110111;
ROM[25319] <= 32'b10111110010000111000001110010011;
ROM[25320] <= 32'b00000000111000111000001110110011;
ROM[25321] <= 32'b00000000011100010010000000100011;
ROM[25322] <= 32'b00000000010000010000000100010011;
ROM[25323] <= 32'b00000000001100010010000000100011;
ROM[25324] <= 32'b00000000010000010000000100010011;
ROM[25325] <= 32'b00000000010000010010000000100011;
ROM[25326] <= 32'b00000000010000010000000100010011;
ROM[25327] <= 32'b00000000010100010010000000100011;
ROM[25328] <= 32'b00000000010000010000000100010011;
ROM[25329] <= 32'b00000000011000010010000000100011;
ROM[25330] <= 32'b00000000010000010000000100010011;
ROM[25331] <= 32'b00000001010000000000001110010011;
ROM[25332] <= 32'b00000000100000111000001110010011;
ROM[25333] <= 32'b01000000011100010000001110110011;
ROM[25334] <= 32'b00000000011100000000001000110011;
ROM[25335] <= 32'b00000000001000000000000110110011;
ROM[25336] <= 32'b01111100110100010000000011101111;
ROM[25337] <= 32'b00000010000000000000001110010011;
ROM[25338] <= 32'b00000000011100010010000000100011;
ROM[25339] <= 32'b00000000010000010000000100010011;
ROM[25340] <= 32'b00000000000000011001001110110111;
ROM[25341] <= 32'b11000011110000111000001110010011;
ROM[25342] <= 32'b00000000111000111000001110110011;
ROM[25343] <= 32'b00000000011100010010000000100011;
ROM[25344] <= 32'b00000000010000010000000100010011;
ROM[25345] <= 32'b00000000001100010010000000100011;
ROM[25346] <= 32'b00000000010000010000000100010011;
ROM[25347] <= 32'b00000000010000010010000000100011;
ROM[25348] <= 32'b00000000010000010000000100010011;
ROM[25349] <= 32'b00000000010100010010000000100011;
ROM[25350] <= 32'b00000000010000010000000100010011;
ROM[25351] <= 32'b00000000011000010010000000100011;
ROM[25352] <= 32'b00000000010000010000000100010011;
ROM[25353] <= 32'b00000001010000000000001110010011;
ROM[25354] <= 32'b00000000100000111000001110010011;
ROM[25355] <= 32'b01000000011100010000001110110011;
ROM[25356] <= 32'b00000000011100000000001000110011;
ROM[25357] <= 32'b00000000001000000000000110110011;
ROM[25358] <= 32'b01110111010100010000000011101111;
ROM[25359] <= 32'b00000110000100000000001110010011;
ROM[25360] <= 32'b00000000011100010010000000100011;
ROM[25361] <= 32'b00000000010000010000000100010011;
ROM[25362] <= 32'b00000000000000011001001110110111;
ROM[25363] <= 32'b11001001010000111000001110010011;
ROM[25364] <= 32'b00000000111000111000001110110011;
ROM[25365] <= 32'b00000000011100010010000000100011;
ROM[25366] <= 32'b00000000010000010000000100010011;
ROM[25367] <= 32'b00000000001100010010000000100011;
ROM[25368] <= 32'b00000000010000010000000100010011;
ROM[25369] <= 32'b00000000010000010010000000100011;
ROM[25370] <= 32'b00000000010000010000000100010011;
ROM[25371] <= 32'b00000000010100010010000000100011;
ROM[25372] <= 32'b00000000010000010000000100010011;
ROM[25373] <= 32'b00000000011000010010000000100011;
ROM[25374] <= 32'b00000000010000010000000100010011;
ROM[25375] <= 32'b00000001010000000000001110010011;
ROM[25376] <= 32'b00000000100000111000001110010011;
ROM[25377] <= 32'b01000000011100010000001110110011;
ROM[25378] <= 32'b00000000011100000000001000110011;
ROM[25379] <= 32'b00000000001000000000000110110011;
ROM[25380] <= 32'b01110001110100010000000011101111;
ROM[25381] <= 32'b00000111001000000000001110010011;
ROM[25382] <= 32'b00000000011100010010000000100011;
ROM[25383] <= 32'b00000000010000010000000100010011;
ROM[25384] <= 32'b00000000000000011001001110110111;
ROM[25385] <= 32'b11001110110000111000001110010011;
ROM[25386] <= 32'b00000000111000111000001110110011;
ROM[25387] <= 32'b00000000011100010010000000100011;
ROM[25388] <= 32'b00000000010000010000000100010011;
ROM[25389] <= 32'b00000000001100010010000000100011;
ROM[25390] <= 32'b00000000010000010000000100010011;
ROM[25391] <= 32'b00000000010000010010000000100011;
ROM[25392] <= 32'b00000000010000010000000100010011;
ROM[25393] <= 32'b00000000010100010010000000100011;
ROM[25394] <= 32'b00000000010000010000000100010011;
ROM[25395] <= 32'b00000000011000010010000000100011;
ROM[25396] <= 32'b00000000010000010000000100010011;
ROM[25397] <= 32'b00000001010000000000001110010011;
ROM[25398] <= 32'b00000000100000111000001110010011;
ROM[25399] <= 32'b01000000011100010000001110110011;
ROM[25400] <= 32'b00000000011100000000001000110011;
ROM[25401] <= 32'b00000000001000000000000110110011;
ROM[25402] <= 32'b01101100010100010000000011101111;
ROM[25403] <= 32'b00000111001000000000001110010011;
ROM[25404] <= 32'b00000000011100010010000000100011;
ROM[25405] <= 32'b00000000010000010000000100010011;
ROM[25406] <= 32'b00000000000000011001001110110111;
ROM[25407] <= 32'b11010100010000111000001110010011;
ROM[25408] <= 32'b00000000111000111000001110110011;
ROM[25409] <= 32'b00000000011100010010000000100011;
ROM[25410] <= 32'b00000000010000010000000100010011;
ROM[25411] <= 32'b00000000001100010010000000100011;
ROM[25412] <= 32'b00000000010000010000000100010011;
ROM[25413] <= 32'b00000000010000010010000000100011;
ROM[25414] <= 32'b00000000010000010000000100010011;
ROM[25415] <= 32'b00000000010100010010000000100011;
ROM[25416] <= 32'b00000000010000010000000100010011;
ROM[25417] <= 32'b00000000011000010010000000100011;
ROM[25418] <= 32'b00000000010000010000000100010011;
ROM[25419] <= 32'b00000001010000000000001110010011;
ROM[25420] <= 32'b00000000100000111000001110010011;
ROM[25421] <= 32'b01000000011100010000001110110011;
ROM[25422] <= 32'b00000000011100000000001000110011;
ROM[25423] <= 32'b00000000001000000000000110110011;
ROM[25424] <= 32'b01100110110100010000000011101111;
ROM[25425] <= 32'b00000110000100000000001110010011;
ROM[25426] <= 32'b00000000011100010010000000100011;
ROM[25427] <= 32'b00000000010000010000000100010011;
ROM[25428] <= 32'b00000000000000011001001110110111;
ROM[25429] <= 32'b11011001110000111000001110010011;
ROM[25430] <= 32'b00000000111000111000001110110011;
ROM[25431] <= 32'b00000000011100010010000000100011;
ROM[25432] <= 32'b00000000010000010000000100010011;
ROM[25433] <= 32'b00000000001100010010000000100011;
ROM[25434] <= 32'b00000000010000010000000100010011;
ROM[25435] <= 32'b00000000010000010010000000100011;
ROM[25436] <= 32'b00000000010000010000000100010011;
ROM[25437] <= 32'b00000000010100010010000000100011;
ROM[25438] <= 32'b00000000010000010000000100010011;
ROM[25439] <= 32'b00000000011000010010000000100011;
ROM[25440] <= 32'b00000000010000010000000100010011;
ROM[25441] <= 32'b00000001010000000000001110010011;
ROM[25442] <= 32'b00000000100000111000001110010011;
ROM[25443] <= 32'b01000000011100010000001110110011;
ROM[25444] <= 32'b00000000011100000000001000110011;
ROM[25445] <= 32'b00000000001000000000000110110011;
ROM[25446] <= 32'b01100001010100010000000011101111;
ROM[25447] <= 32'b00000111100100000000001110010011;
ROM[25448] <= 32'b00000000011100010010000000100011;
ROM[25449] <= 32'b00000000010000010000000100010011;
ROM[25450] <= 32'b00000000000000011001001110110111;
ROM[25451] <= 32'b11011111010000111000001110010011;
ROM[25452] <= 32'b00000000111000111000001110110011;
ROM[25453] <= 32'b00000000011100010010000000100011;
ROM[25454] <= 32'b00000000010000010000000100010011;
ROM[25455] <= 32'b00000000001100010010000000100011;
ROM[25456] <= 32'b00000000010000010000000100010011;
ROM[25457] <= 32'b00000000010000010010000000100011;
ROM[25458] <= 32'b00000000010000010000000100010011;
ROM[25459] <= 32'b00000000010100010010000000100011;
ROM[25460] <= 32'b00000000010000010000000100010011;
ROM[25461] <= 32'b00000000011000010010000000100011;
ROM[25462] <= 32'b00000000010000010000000100010011;
ROM[25463] <= 32'b00000001010000000000001110010011;
ROM[25464] <= 32'b00000000100000111000001110010011;
ROM[25465] <= 32'b01000000011100010000001110110011;
ROM[25466] <= 32'b00000000011100000000001000110011;
ROM[25467] <= 32'b00000000001000000000000110110011;
ROM[25468] <= 32'b01011011110100010000000011101111;
ROM[25469] <= 32'b00000011101000000000001110010011;
ROM[25470] <= 32'b00000000011100010010000000100011;
ROM[25471] <= 32'b00000000010000010000000100010011;
ROM[25472] <= 32'b00000000000000011001001110110111;
ROM[25473] <= 32'b11100100110000111000001110010011;
ROM[25474] <= 32'b00000000111000111000001110110011;
ROM[25475] <= 32'b00000000011100010010000000100011;
ROM[25476] <= 32'b00000000010000010000000100010011;
ROM[25477] <= 32'b00000000001100010010000000100011;
ROM[25478] <= 32'b00000000010000010000000100010011;
ROM[25479] <= 32'b00000000010000010010000000100011;
ROM[25480] <= 32'b00000000010000010000000100010011;
ROM[25481] <= 32'b00000000010100010010000000100011;
ROM[25482] <= 32'b00000000010000010000000100010011;
ROM[25483] <= 32'b00000000011000010010000000100011;
ROM[25484] <= 32'b00000000010000010000000100010011;
ROM[25485] <= 32'b00000001010000000000001110010011;
ROM[25486] <= 32'b00000000100000111000001110010011;
ROM[25487] <= 32'b01000000011100010000001110110011;
ROM[25488] <= 32'b00000000011100000000001000110011;
ROM[25489] <= 32'b00000000001000000000000110110011;
ROM[25490] <= 32'b01010110010100010000000011101111;
ROM[25491] <= 32'b00000010000000000000001110010011;
ROM[25492] <= 32'b00000000011100010010000000100011;
ROM[25493] <= 32'b00000000010000010000000100010011;
ROM[25494] <= 32'b00000000000000011001001110110111;
ROM[25495] <= 32'b11101010010000111000001110010011;
ROM[25496] <= 32'b00000000111000111000001110110011;
ROM[25497] <= 32'b00000000011100010010000000100011;
ROM[25498] <= 32'b00000000010000010000000100010011;
ROM[25499] <= 32'b00000000001100010010000000100011;
ROM[25500] <= 32'b00000000010000010000000100010011;
ROM[25501] <= 32'b00000000010000010010000000100011;
ROM[25502] <= 32'b00000000010000010000000100010011;
ROM[25503] <= 32'b00000000010100010010000000100011;
ROM[25504] <= 32'b00000000010000010000000100010011;
ROM[25505] <= 32'b00000000011000010010000000100011;
ROM[25506] <= 32'b00000000010000010000000100010011;
ROM[25507] <= 32'b00000001010000000000001110010011;
ROM[25508] <= 32'b00000000100000111000001110010011;
ROM[25509] <= 32'b01000000011100010000001110110011;
ROM[25510] <= 32'b00000000011100000000001000110011;
ROM[25511] <= 32'b00000000001000000000000110110011;
ROM[25512] <= 32'b01010000110100010000000011101111;
ROM[25513] <= 32'b00000000000000011001001110110111;
ROM[25514] <= 32'b11101111000000111000001110010011;
ROM[25515] <= 32'b00000000111000111000001110110011;
ROM[25516] <= 32'b00000000011100010010000000100011;
ROM[25517] <= 32'b00000000010000010000000100010011;
ROM[25518] <= 32'b00000000001100010010000000100011;
ROM[25519] <= 32'b00000000010000010000000100010011;
ROM[25520] <= 32'b00000000010000010010000000100011;
ROM[25521] <= 32'b00000000010000010000000100010011;
ROM[25522] <= 32'b00000000010100010010000000100011;
ROM[25523] <= 32'b00000000010000010000000100010011;
ROM[25524] <= 32'b00000000011000010010000000100011;
ROM[25525] <= 32'b00000000010000010000000100010011;
ROM[25526] <= 32'b00000001010000000000001110010011;
ROM[25527] <= 32'b00000000010000111000001110010011;
ROM[25528] <= 32'b01000000011100010000001110110011;
ROM[25529] <= 32'b00000000011100000000001000110011;
ROM[25530] <= 32'b00000000001000000000000110110011;
ROM[25531] <= 32'b10011101110011110101000011101111;
ROM[25532] <= 32'b11111111110000010000000100010011;
ROM[25533] <= 32'b00000000000000010010001110000011;
ROM[25534] <= 32'b00000000011100011010001000100011;
ROM[25535] <= 32'b00000000010000011010001110000011;
ROM[25536] <= 32'b00000000011100010010000000100011;
ROM[25537] <= 32'b00000000010000010000000100010011;
ROM[25538] <= 32'b00000000000000011001001110110111;
ROM[25539] <= 32'b11110101010000111000001110010011;
ROM[25540] <= 32'b00000000111000111000001110110011;
ROM[25541] <= 32'b00000000011100010010000000100011;
ROM[25542] <= 32'b00000000010000010000000100010011;
ROM[25543] <= 32'b00000000001100010010000000100011;
ROM[25544] <= 32'b00000000010000010000000100010011;
ROM[25545] <= 32'b00000000010000010010000000100011;
ROM[25546] <= 32'b00000000010000010000000100010011;
ROM[25547] <= 32'b00000000010100010010000000100011;
ROM[25548] <= 32'b00000000010000010000000100010011;
ROM[25549] <= 32'b00000000011000010010000000100011;
ROM[25550] <= 32'b00000000010000010000000100010011;
ROM[25551] <= 32'b00000001010000000000001110010011;
ROM[25552] <= 32'b00000000010000111000001110010011;
ROM[25553] <= 32'b01000000011100010000001110110011;
ROM[25554] <= 32'b00000000011100000000001000110011;
ROM[25555] <= 32'b00000000001000000000000110110011;
ROM[25556] <= 32'b10010011000011100111000011101111;
ROM[25557] <= 32'b11111111110000010000000100010011;
ROM[25558] <= 32'b00000000000000010010001110000011;
ROM[25559] <= 32'b00000000011100011010000000100011;
ROM[25560] <= 32'b00000010000100000000001110010011;
ROM[25561] <= 32'b00000000011100010010000000100011;
ROM[25562] <= 32'b00000000010000010000000100010011;
ROM[25563] <= 32'b00000000000000011001001110110111;
ROM[25564] <= 32'b11111011100000111000001110010011;
ROM[25565] <= 32'b00000000111000111000001110110011;
ROM[25566] <= 32'b00000000011100010010000000100011;
ROM[25567] <= 32'b00000000010000010000000100010011;
ROM[25568] <= 32'b00000000001100010010000000100011;
ROM[25569] <= 32'b00000000010000010000000100010011;
ROM[25570] <= 32'b00000000010000010010000000100011;
ROM[25571] <= 32'b00000000010000010000000100010011;
ROM[25572] <= 32'b00000000010100010010000000100011;
ROM[25573] <= 32'b00000000010000010000000100010011;
ROM[25574] <= 32'b00000000011000010010000000100011;
ROM[25575] <= 32'b00000000010000010000000100010011;
ROM[25576] <= 32'b00000001010000000000001110010011;
ROM[25577] <= 32'b00000000010000111000001110010011;
ROM[25578] <= 32'b01000000011100010000001110110011;
ROM[25579] <= 32'b00000000011100000000001000110011;
ROM[25580] <= 32'b00000000001000000000000110110011;
ROM[25581] <= 32'b01111000100000010000000011101111;
ROM[25582] <= 32'b00000100010100000000001110010011;
ROM[25583] <= 32'b00000000011100010010000000100011;
ROM[25584] <= 32'b00000000010000010000000100010011;
ROM[25585] <= 32'b00000000000000011001001110110111;
ROM[25586] <= 32'b00000001000000111000001110010011;
ROM[25587] <= 32'b00000000111000111000001110110011;
ROM[25588] <= 32'b00000000011100010010000000100011;
ROM[25589] <= 32'b00000000010000010000000100010011;
ROM[25590] <= 32'b00000000001100010010000000100011;
ROM[25591] <= 32'b00000000010000010000000100010011;
ROM[25592] <= 32'b00000000010000010010000000100011;
ROM[25593] <= 32'b00000000010000010000000100010011;
ROM[25594] <= 32'b00000000010100010010000000100011;
ROM[25595] <= 32'b00000000010000010000000100010011;
ROM[25596] <= 32'b00000000011000010010000000100011;
ROM[25597] <= 32'b00000000010000010000000100010011;
ROM[25598] <= 32'b00000001010000000000001110010011;
ROM[25599] <= 32'b00000000100000111000001110010011;
ROM[25600] <= 32'b01000000011100010000001110110011;
ROM[25601] <= 32'b00000000011100000000001000110011;
ROM[25602] <= 32'b00000000001000000000000110110011;
ROM[25603] <= 32'b00111010000100010000000011101111;
ROM[25604] <= 32'b00000110111000000000001110010011;
ROM[25605] <= 32'b00000000011100010010000000100011;
ROM[25606] <= 32'b00000000010000010000000100010011;
ROM[25607] <= 32'b00000000000000011001001110110111;
ROM[25608] <= 32'b00000110100000111000001110010011;
ROM[25609] <= 32'b00000000111000111000001110110011;
ROM[25610] <= 32'b00000000011100010010000000100011;
ROM[25611] <= 32'b00000000010000010000000100010011;
ROM[25612] <= 32'b00000000001100010010000000100011;
ROM[25613] <= 32'b00000000010000010000000100010011;
ROM[25614] <= 32'b00000000010000010010000000100011;
ROM[25615] <= 32'b00000000010000010000000100010011;
ROM[25616] <= 32'b00000000010100010010000000100011;
ROM[25617] <= 32'b00000000010000010000000100010011;
ROM[25618] <= 32'b00000000011000010010000000100011;
ROM[25619] <= 32'b00000000010000010000000100010011;
ROM[25620] <= 32'b00000001010000000000001110010011;
ROM[25621] <= 32'b00000000100000111000001110010011;
ROM[25622] <= 32'b01000000011100010000001110110011;
ROM[25623] <= 32'b00000000011100000000001000110011;
ROM[25624] <= 32'b00000000001000000000000110110011;
ROM[25625] <= 32'b00110100100100010000000011101111;
ROM[25626] <= 32'b00000111010000000000001110010011;
ROM[25627] <= 32'b00000000011100010010000000100011;
ROM[25628] <= 32'b00000000010000010000000100010011;
ROM[25629] <= 32'b00000000000000011001001110110111;
ROM[25630] <= 32'b00001100000000111000001110010011;
ROM[25631] <= 32'b00000000111000111000001110110011;
ROM[25632] <= 32'b00000000011100010010000000100011;
ROM[25633] <= 32'b00000000010000010000000100010011;
ROM[25634] <= 32'b00000000001100010010000000100011;
ROM[25635] <= 32'b00000000010000010000000100010011;
ROM[25636] <= 32'b00000000010000010010000000100011;
ROM[25637] <= 32'b00000000010000010000000100010011;
ROM[25638] <= 32'b00000000010100010010000000100011;
ROM[25639] <= 32'b00000000010000010000000100010011;
ROM[25640] <= 32'b00000000011000010010000000100011;
ROM[25641] <= 32'b00000000010000010000000100010011;
ROM[25642] <= 32'b00000001010000000000001110010011;
ROM[25643] <= 32'b00000000100000111000001110010011;
ROM[25644] <= 32'b01000000011100010000001110110011;
ROM[25645] <= 32'b00000000011100000000001000110011;
ROM[25646] <= 32'b00000000001000000000000110110011;
ROM[25647] <= 32'b00101111000100010000000011101111;
ROM[25648] <= 32'b00000110010100000000001110010011;
ROM[25649] <= 32'b00000000011100010010000000100011;
ROM[25650] <= 32'b00000000010000010000000100010011;
ROM[25651] <= 32'b00000000000000011001001110110111;
ROM[25652] <= 32'b00010001100000111000001110010011;
ROM[25653] <= 32'b00000000111000111000001110110011;
ROM[25654] <= 32'b00000000011100010010000000100011;
ROM[25655] <= 32'b00000000010000010000000100010011;
ROM[25656] <= 32'b00000000001100010010000000100011;
ROM[25657] <= 32'b00000000010000010000000100010011;
ROM[25658] <= 32'b00000000010000010010000000100011;
ROM[25659] <= 32'b00000000010000010000000100010011;
ROM[25660] <= 32'b00000000010100010010000000100011;
ROM[25661] <= 32'b00000000010000010000000100010011;
ROM[25662] <= 32'b00000000011000010010000000100011;
ROM[25663] <= 32'b00000000010000010000000100010011;
ROM[25664] <= 32'b00000001010000000000001110010011;
ROM[25665] <= 32'b00000000100000111000001110010011;
ROM[25666] <= 32'b01000000011100010000001110110011;
ROM[25667] <= 32'b00000000011100000000001000110011;
ROM[25668] <= 32'b00000000001000000000000110110011;
ROM[25669] <= 32'b00101001100100010000000011101111;
ROM[25670] <= 32'b00000111001000000000001110010011;
ROM[25671] <= 32'b00000000011100010010000000100011;
ROM[25672] <= 32'b00000000010000010000000100010011;
ROM[25673] <= 32'b00000000000000011001001110110111;
ROM[25674] <= 32'b00010111000000111000001110010011;
ROM[25675] <= 32'b00000000111000111000001110110011;
ROM[25676] <= 32'b00000000011100010010000000100011;
ROM[25677] <= 32'b00000000010000010000000100010011;
ROM[25678] <= 32'b00000000001100010010000000100011;
ROM[25679] <= 32'b00000000010000010000000100010011;
ROM[25680] <= 32'b00000000010000010010000000100011;
ROM[25681] <= 32'b00000000010000010000000100010011;
ROM[25682] <= 32'b00000000010100010010000000100011;
ROM[25683] <= 32'b00000000010000010000000100010011;
ROM[25684] <= 32'b00000000011000010010000000100011;
ROM[25685] <= 32'b00000000010000010000000100010011;
ROM[25686] <= 32'b00000001010000000000001110010011;
ROM[25687] <= 32'b00000000100000111000001110010011;
ROM[25688] <= 32'b01000000011100010000001110110011;
ROM[25689] <= 32'b00000000011100000000001000110011;
ROM[25690] <= 32'b00000000001000000000000110110011;
ROM[25691] <= 32'b00100100000100010000000011101111;
ROM[25692] <= 32'b00000010000000000000001110010011;
ROM[25693] <= 32'b00000000011100010010000000100011;
ROM[25694] <= 32'b00000000010000010000000100010011;
ROM[25695] <= 32'b00000000000000011001001110110111;
ROM[25696] <= 32'b00011100100000111000001110010011;
ROM[25697] <= 32'b00000000111000111000001110110011;
ROM[25698] <= 32'b00000000011100010010000000100011;
ROM[25699] <= 32'b00000000010000010000000100010011;
ROM[25700] <= 32'b00000000001100010010000000100011;
ROM[25701] <= 32'b00000000010000010000000100010011;
ROM[25702] <= 32'b00000000010000010010000000100011;
ROM[25703] <= 32'b00000000010000010000000100010011;
ROM[25704] <= 32'b00000000010100010010000000100011;
ROM[25705] <= 32'b00000000010000010000000100010011;
ROM[25706] <= 32'b00000000011000010010000000100011;
ROM[25707] <= 32'b00000000010000010000000100010011;
ROM[25708] <= 32'b00000001010000000000001110010011;
ROM[25709] <= 32'b00000000100000111000001110010011;
ROM[25710] <= 32'b01000000011100010000001110110011;
ROM[25711] <= 32'b00000000011100000000001000110011;
ROM[25712] <= 32'b00000000001000000000000110110011;
ROM[25713] <= 32'b00011110100100010000000011101111;
ROM[25714] <= 32'b00000111010000000000001110010011;
ROM[25715] <= 32'b00000000011100010010000000100011;
ROM[25716] <= 32'b00000000010000010000000100010011;
ROM[25717] <= 32'b00000000000000011001001110110111;
ROM[25718] <= 32'b00100010000000111000001110010011;
ROM[25719] <= 32'b00000000111000111000001110110011;
ROM[25720] <= 32'b00000000011100010010000000100011;
ROM[25721] <= 32'b00000000010000010000000100010011;
ROM[25722] <= 32'b00000000001100010010000000100011;
ROM[25723] <= 32'b00000000010000010000000100010011;
ROM[25724] <= 32'b00000000010000010010000000100011;
ROM[25725] <= 32'b00000000010000010000000100010011;
ROM[25726] <= 32'b00000000010100010010000000100011;
ROM[25727] <= 32'b00000000010000010000000100010011;
ROM[25728] <= 32'b00000000011000010010000000100011;
ROM[25729] <= 32'b00000000010000010000000100010011;
ROM[25730] <= 32'b00000001010000000000001110010011;
ROM[25731] <= 32'b00000000100000111000001110010011;
ROM[25732] <= 32'b01000000011100010000001110110011;
ROM[25733] <= 32'b00000000011100000000001000110011;
ROM[25734] <= 32'b00000000001000000000000110110011;
ROM[25735] <= 32'b00011001000100010000000011101111;
ROM[25736] <= 32'b00000110100000000000001110010011;
ROM[25737] <= 32'b00000000011100010010000000100011;
ROM[25738] <= 32'b00000000010000010000000100010011;
ROM[25739] <= 32'b00000000000000011001001110110111;
ROM[25740] <= 32'b00100111100000111000001110010011;
ROM[25741] <= 32'b00000000111000111000001110110011;
ROM[25742] <= 32'b00000000011100010010000000100011;
ROM[25743] <= 32'b00000000010000010000000100010011;
ROM[25744] <= 32'b00000000001100010010000000100011;
ROM[25745] <= 32'b00000000010000010000000100010011;
ROM[25746] <= 32'b00000000010000010010000000100011;
ROM[25747] <= 32'b00000000010000010000000100010011;
ROM[25748] <= 32'b00000000010100010010000000100011;
ROM[25749] <= 32'b00000000010000010000000100010011;
ROM[25750] <= 32'b00000000011000010010000000100011;
ROM[25751] <= 32'b00000000010000010000000100010011;
ROM[25752] <= 32'b00000001010000000000001110010011;
ROM[25753] <= 32'b00000000100000111000001110010011;
ROM[25754] <= 32'b01000000011100010000001110110011;
ROM[25755] <= 32'b00000000011100000000001000110011;
ROM[25756] <= 32'b00000000001000000000000110110011;
ROM[25757] <= 32'b00010011100100010000000011101111;
ROM[25758] <= 32'b00000110010100000000001110010011;
ROM[25759] <= 32'b00000000011100010010000000100011;
ROM[25760] <= 32'b00000000010000010000000100010011;
ROM[25761] <= 32'b00000000000000011001001110110111;
ROM[25762] <= 32'b00101101000000111000001110010011;
ROM[25763] <= 32'b00000000111000111000001110110011;
ROM[25764] <= 32'b00000000011100010010000000100011;
ROM[25765] <= 32'b00000000010000010000000100010011;
ROM[25766] <= 32'b00000000001100010010000000100011;
ROM[25767] <= 32'b00000000010000010000000100010011;
ROM[25768] <= 32'b00000000010000010010000000100011;
ROM[25769] <= 32'b00000000010000010000000100010011;
ROM[25770] <= 32'b00000000010100010010000000100011;
ROM[25771] <= 32'b00000000010000010000000100010011;
ROM[25772] <= 32'b00000000011000010010000000100011;
ROM[25773] <= 32'b00000000010000010000000100010011;
ROM[25774] <= 32'b00000001010000000000001110010011;
ROM[25775] <= 32'b00000000100000111000001110010011;
ROM[25776] <= 32'b01000000011100010000001110110011;
ROM[25777] <= 32'b00000000011100000000001000110011;
ROM[25778] <= 32'b00000000001000000000000110110011;
ROM[25779] <= 32'b00001110000100010000000011101111;
ROM[25780] <= 32'b00000010000000000000001110010011;
ROM[25781] <= 32'b00000000011100010010000000100011;
ROM[25782] <= 32'b00000000010000010000000100010011;
ROM[25783] <= 32'b00000000000000011001001110110111;
ROM[25784] <= 32'b00110010100000111000001110010011;
ROM[25785] <= 32'b00000000111000111000001110110011;
ROM[25786] <= 32'b00000000011100010010000000100011;
ROM[25787] <= 32'b00000000010000010000000100010011;
ROM[25788] <= 32'b00000000001100010010000000100011;
ROM[25789] <= 32'b00000000010000010000000100010011;
ROM[25790] <= 32'b00000000010000010010000000100011;
ROM[25791] <= 32'b00000000010000010000000100010011;
ROM[25792] <= 32'b00000000010100010010000000100011;
ROM[25793] <= 32'b00000000010000010000000100010011;
ROM[25794] <= 32'b00000000011000010010000000100011;
ROM[25795] <= 32'b00000000010000010000000100010011;
ROM[25796] <= 32'b00000001010000000000001110010011;
ROM[25797] <= 32'b00000000100000111000001110010011;
ROM[25798] <= 32'b01000000011100010000001110110011;
ROM[25799] <= 32'b00000000011100000000001000110011;
ROM[25800] <= 32'b00000000001000000000000110110011;
ROM[25801] <= 32'b00001000100100010000000011101111;
ROM[25802] <= 32'b00000110010100000000001110010011;
ROM[25803] <= 32'b00000000011100010010000000100011;
ROM[25804] <= 32'b00000000010000010000000100010011;
ROM[25805] <= 32'b00000000000000011001001110110111;
ROM[25806] <= 32'b00111000000000111000001110010011;
ROM[25807] <= 32'b00000000111000111000001110110011;
ROM[25808] <= 32'b00000000011100010010000000100011;
ROM[25809] <= 32'b00000000010000010000000100010011;
ROM[25810] <= 32'b00000000001100010010000000100011;
ROM[25811] <= 32'b00000000010000010000000100010011;
ROM[25812] <= 32'b00000000010000010010000000100011;
ROM[25813] <= 32'b00000000010000010000000100010011;
ROM[25814] <= 32'b00000000010100010010000000100011;
ROM[25815] <= 32'b00000000010000010000000100010011;
ROM[25816] <= 32'b00000000011000010010000000100011;
ROM[25817] <= 32'b00000000010000010000000100010011;
ROM[25818] <= 32'b00000001010000000000001110010011;
ROM[25819] <= 32'b00000000100000111000001110010011;
ROM[25820] <= 32'b01000000011100010000001110110011;
ROM[25821] <= 32'b00000000011100000000001000110011;
ROM[25822] <= 32'b00000000001000000000000110110011;
ROM[25823] <= 32'b00000011000100010000000011101111;
ROM[25824] <= 32'b00000110110000000000001110010011;
ROM[25825] <= 32'b00000000011100010010000000100011;
ROM[25826] <= 32'b00000000010000010000000100010011;
ROM[25827] <= 32'b00000000000000011001001110110111;
ROM[25828] <= 32'b00111101100000111000001110010011;
ROM[25829] <= 32'b00000000111000111000001110110011;
ROM[25830] <= 32'b00000000011100010010000000100011;
ROM[25831] <= 32'b00000000010000010000000100010011;
ROM[25832] <= 32'b00000000001100010010000000100011;
ROM[25833] <= 32'b00000000010000010000000100010011;
ROM[25834] <= 32'b00000000010000010010000000100011;
ROM[25835] <= 32'b00000000010000010000000100010011;
ROM[25836] <= 32'b00000000010100010010000000100011;
ROM[25837] <= 32'b00000000010000010000000100010011;
ROM[25838] <= 32'b00000000011000010010000000100011;
ROM[25839] <= 32'b00000000010000010000000100010011;
ROM[25840] <= 32'b00000001010000000000001110010011;
ROM[25841] <= 32'b00000000100000111000001110010011;
ROM[25842] <= 32'b01000000011100010000001110110011;
ROM[25843] <= 32'b00000000011100000000001000110011;
ROM[25844] <= 32'b00000000001000000000000110110011;
ROM[25845] <= 32'b01111101100000010000000011101111;
ROM[25846] <= 32'b00000110010100000000001110010011;
ROM[25847] <= 32'b00000000011100010010000000100011;
ROM[25848] <= 32'b00000000010000010000000100010011;
ROM[25849] <= 32'b00000000000000011001001110110111;
ROM[25850] <= 32'b01000011000000111000001110010011;
ROM[25851] <= 32'b00000000111000111000001110110011;
ROM[25852] <= 32'b00000000011100010010000000100011;
ROM[25853] <= 32'b00000000010000010000000100010011;
ROM[25854] <= 32'b00000000001100010010000000100011;
ROM[25855] <= 32'b00000000010000010000000100010011;
ROM[25856] <= 32'b00000000010000010010000000100011;
ROM[25857] <= 32'b00000000010000010000000100010011;
ROM[25858] <= 32'b00000000010100010010000000100011;
ROM[25859] <= 32'b00000000010000010000000100010011;
ROM[25860] <= 32'b00000000011000010010000000100011;
ROM[25861] <= 32'b00000000010000010000000100010011;
ROM[25862] <= 32'b00000001010000000000001110010011;
ROM[25863] <= 32'b00000000100000111000001110010011;
ROM[25864] <= 32'b01000000011100010000001110110011;
ROM[25865] <= 32'b00000000011100000000001000110011;
ROM[25866] <= 32'b00000000001000000000000110110011;
ROM[25867] <= 32'b01111000000000010000000011101111;
ROM[25868] <= 32'b00000110110100000000001110010011;
ROM[25869] <= 32'b00000000011100010010000000100011;
ROM[25870] <= 32'b00000000010000010000000100010011;
ROM[25871] <= 32'b00000000000000011001001110110111;
ROM[25872] <= 32'b01001000100000111000001110010011;
ROM[25873] <= 32'b00000000111000111000001110110011;
ROM[25874] <= 32'b00000000011100010010000000100011;
ROM[25875] <= 32'b00000000010000010000000100010011;
ROM[25876] <= 32'b00000000001100010010000000100011;
ROM[25877] <= 32'b00000000010000010000000100010011;
ROM[25878] <= 32'b00000000010000010010000000100011;
ROM[25879] <= 32'b00000000010000010000000100010011;
ROM[25880] <= 32'b00000000010100010010000000100011;
ROM[25881] <= 32'b00000000010000010000000100010011;
ROM[25882] <= 32'b00000000011000010010000000100011;
ROM[25883] <= 32'b00000000010000010000000100010011;
ROM[25884] <= 32'b00000001010000000000001110010011;
ROM[25885] <= 32'b00000000100000111000001110010011;
ROM[25886] <= 32'b01000000011100010000001110110011;
ROM[25887] <= 32'b00000000011100000000001000110011;
ROM[25888] <= 32'b00000000001000000000000110110011;
ROM[25889] <= 32'b01110010100000010000000011101111;
ROM[25890] <= 32'b00000110010100000000001110010011;
ROM[25891] <= 32'b00000000011100010010000000100011;
ROM[25892] <= 32'b00000000010000010000000100010011;
ROM[25893] <= 32'b00000000000000011001001110110111;
ROM[25894] <= 32'b01001110000000111000001110010011;
ROM[25895] <= 32'b00000000111000111000001110110011;
ROM[25896] <= 32'b00000000011100010010000000100011;
ROM[25897] <= 32'b00000000010000010000000100010011;
ROM[25898] <= 32'b00000000001100010010000000100011;
ROM[25899] <= 32'b00000000010000010000000100010011;
ROM[25900] <= 32'b00000000010000010010000000100011;
ROM[25901] <= 32'b00000000010000010000000100010011;
ROM[25902] <= 32'b00000000010100010010000000100011;
ROM[25903] <= 32'b00000000010000010000000100010011;
ROM[25904] <= 32'b00000000011000010010000000100011;
ROM[25905] <= 32'b00000000010000010000000100010011;
ROM[25906] <= 32'b00000001010000000000001110010011;
ROM[25907] <= 32'b00000000100000111000001110010011;
ROM[25908] <= 32'b01000000011100010000001110110011;
ROM[25909] <= 32'b00000000011100000000001000110011;
ROM[25910] <= 32'b00000000001000000000000110110011;
ROM[25911] <= 32'b01101101000000010000000011101111;
ROM[25912] <= 32'b00000110111000000000001110010011;
ROM[25913] <= 32'b00000000011100010010000000100011;
ROM[25914] <= 32'b00000000010000010000000100010011;
ROM[25915] <= 32'b00000000000000011001001110110111;
ROM[25916] <= 32'b01010011100000111000001110010011;
ROM[25917] <= 32'b00000000111000111000001110110011;
ROM[25918] <= 32'b00000000011100010010000000100011;
ROM[25919] <= 32'b00000000010000010000000100010011;
ROM[25920] <= 32'b00000000001100010010000000100011;
ROM[25921] <= 32'b00000000010000010000000100010011;
ROM[25922] <= 32'b00000000010000010010000000100011;
ROM[25923] <= 32'b00000000010000010000000100010011;
ROM[25924] <= 32'b00000000010100010010000000100011;
ROM[25925] <= 32'b00000000010000010000000100010011;
ROM[25926] <= 32'b00000000011000010010000000100011;
ROM[25927] <= 32'b00000000010000010000000100010011;
ROM[25928] <= 32'b00000001010000000000001110010011;
ROM[25929] <= 32'b00000000100000111000001110010011;
ROM[25930] <= 32'b01000000011100010000001110110011;
ROM[25931] <= 32'b00000000011100000000001000110011;
ROM[25932] <= 32'b00000000001000000000000110110011;
ROM[25933] <= 32'b01100111100000010000000011101111;
ROM[25934] <= 32'b00000111010000000000001110010011;
ROM[25935] <= 32'b00000000011100010010000000100011;
ROM[25936] <= 32'b00000000010000010000000100010011;
ROM[25937] <= 32'b00000000000000011001001110110111;
ROM[25938] <= 32'b01011001000000111000001110010011;
ROM[25939] <= 32'b00000000111000111000001110110011;
ROM[25940] <= 32'b00000000011100010010000000100011;
ROM[25941] <= 32'b00000000010000010000000100010011;
ROM[25942] <= 32'b00000000001100010010000000100011;
ROM[25943] <= 32'b00000000010000010000000100010011;
ROM[25944] <= 32'b00000000010000010010000000100011;
ROM[25945] <= 32'b00000000010000010000000100010011;
ROM[25946] <= 32'b00000000010100010010000000100011;
ROM[25947] <= 32'b00000000010000010000000100010011;
ROM[25948] <= 32'b00000000011000010010000000100011;
ROM[25949] <= 32'b00000000010000010000000100010011;
ROM[25950] <= 32'b00000001010000000000001110010011;
ROM[25951] <= 32'b00000000100000111000001110010011;
ROM[25952] <= 32'b01000000011100010000001110110011;
ROM[25953] <= 32'b00000000011100000000001000110011;
ROM[25954] <= 32'b00000000001000000000000110110011;
ROM[25955] <= 32'b01100010000000010000000011101111;
ROM[25956] <= 32'b00000111001100000000001110010011;
ROM[25957] <= 32'b00000000011100010010000000100011;
ROM[25958] <= 32'b00000000010000010000000100010011;
ROM[25959] <= 32'b00000000000000011001001110110111;
ROM[25960] <= 32'b01011110100000111000001110010011;
ROM[25961] <= 32'b00000000111000111000001110110011;
ROM[25962] <= 32'b00000000011100010010000000100011;
ROM[25963] <= 32'b00000000010000010000000100010011;
ROM[25964] <= 32'b00000000001100010010000000100011;
ROM[25965] <= 32'b00000000010000010000000100010011;
ROM[25966] <= 32'b00000000010000010010000000100011;
ROM[25967] <= 32'b00000000010000010000000100010011;
ROM[25968] <= 32'b00000000010100010010000000100011;
ROM[25969] <= 32'b00000000010000010000000100010011;
ROM[25970] <= 32'b00000000011000010010000000100011;
ROM[25971] <= 32'b00000000010000010000000100010011;
ROM[25972] <= 32'b00000001010000000000001110010011;
ROM[25973] <= 32'b00000000100000111000001110010011;
ROM[25974] <= 32'b01000000011100010000001110110011;
ROM[25975] <= 32'b00000000011100000000001000110011;
ROM[25976] <= 32'b00000000001000000000000110110011;
ROM[25977] <= 32'b01011100100000010000000011101111;
ROM[25978] <= 32'b00000010000000000000001110010011;
ROM[25979] <= 32'b00000000011100010010000000100011;
ROM[25980] <= 32'b00000000010000010000000100010011;
ROM[25981] <= 32'b00000000000000011001001110110111;
ROM[25982] <= 32'b01100100000000111000001110010011;
ROM[25983] <= 32'b00000000111000111000001110110011;
ROM[25984] <= 32'b00000000011100010010000000100011;
ROM[25985] <= 32'b00000000010000010000000100010011;
ROM[25986] <= 32'b00000000001100010010000000100011;
ROM[25987] <= 32'b00000000010000010000000100010011;
ROM[25988] <= 32'b00000000010000010010000000100011;
ROM[25989] <= 32'b00000000010000010000000100010011;
ROM[25990] <= 32'b00000000010100010010000000100011;
ROM[25991] <= 32'b00000000010000010000000100010011;
ROM[25992] <= 32'b00000000011000010010000000100011;
ROM[25993] <= 32'b00000000010000010000000100010011;
ROM[25994] <= 32'b00000001010000000000001110010011;
ROM[25995] <= 32'b00000000100000111000001110010011;
ROM[25996] <= 32'b01000000011100010000001110110011;
ROM[25997] <= 32'b00000000011100000000001000110011;
ROM[25998] <= 32'b00000000001000000000000110110011;
ROM[25999] <= 32'b01010111000000010000000011101111;
ROM[26000] <= 32'b00000110111100000000001110010011;
ROM[26001] <= 32'b00000000011100010010000000100011;
ROM[26002] <= 32'b00000000010000010000000100010011;
ROM[26003] <= 32'b00000000000000011001001110110111;
ROM[26004] <= 32'b01101001100000111000001110010011;
ROM[26005] <= 32'b00000000111000111000001110110011;
ROM[26006] <= 32'b00000000011100010010000000100011;
ROM[26007] <= 32'b00000000010000010000000100010011;
ROM[26008] <= 32'b00000000001100010010000000100011;
ROM[26009] <= 32'b00000000010000010000000100010011;
ROM[26010] <= 32'b00000000010000010010000000100011;
ROM[26011] <= 32'b00000000010000010000000100010011;
ROM[26012] <= 32'b00000000010100010010000000100011;
ROM[26013] <= 32'b00000000010000010000000100010011;
ROM[26014] <= 32'b00000000011000010010000000100011;
ROM[26015] <= 32'b00000000010000010000000100010011;
ROM[26016] <= 32'b00000001010000000000001110010011;
ROM[26017] <= 32'b00000000100000111000001110010011;
ROM[26018] <= 32'b01000000011100010000001110110011;
ROM[26019] <= 32'b00000000011100000000001000110011;
ROM[26020] <= 32'b00000000001000000000000110110011;
ROM[26021] <= 32'b01010001100000010000000011101111;
ROM[26022] <= 32'b00000110011000000000001110010011;
ROM[26023] <= 32'b00000000011100010010000000100011;
ROM[26024] <= 32'b00000000010000010000000100010011;
ROM[26025] <= 32'b00000000000000011001001110110111;
ROM[26026] <= 32'b01101111000000111000001110010011;
ROM[26027] <= 32'b00000000111000111000001110110011;
ROM[26028] <= 32'b00000000011100010010000000100011;
ROM[26029] <= 32'b00000000010000010000000100010011;
ROM[26030] <= 32'b00000000001100010010000000100011;
ROM[26031] <= 32'b00000000010000010000000100010011;
ROM[26032] <= 32'b00000000010000010010000000100011;
ROM[26033] <= 32'b00000000010000010000000100010011;
ROM[26034] <= 32'b00000000010100010010000000100011;
ROM[26035] <= 32'b00000000010000010000000100010011;
ROM[26036] <= 32'b00000000011000010010000000100011;
ROM[26037] <= 32'b00000000010000010000000100010011;
ROM[26038] <= 32'b00000001010000000000001110010011;
ROM[26039] <= 32'b00000000100000111000001110010011;
ROM[26040] <= 32'b01000000011100010000001110110011;
ROM[26041] <= 32'b00000000011100000000001000110011;
ROM[26042] <= 32'b00000000001000000000000110110011;
ROM[26043] <= 32'b01001100000000010000000011101111;
ROM[26044] <= 32'b00000010000000000000001110010011;
ROM[26045] <= 32'b00000000011100010010000000100011;
ROM[26046] <= 32'b00000000010000010000000100010011;
ROM[26047] <= 32'b00000000000000011001001110110111;
ROM[26048] <= 32'b01110100100000111000001110010011;
ROM[26049] <= 32'b00000000111000111000001110110011;
ROM[26050] <= 32'b00000000011100010010000000100011;
ROM[26051] <= 32'b00000000010000010000000100010011;
ROM[26052] <= 32'b00000000001100010010000000100011;
ROM[26053] <= 32'b00000000010000010000000100010011;
ROM[26054] <= 32'b00000000010000010010000000100011;
ROM[26055] <= 32'b00000000010000010000000100010011;
ROM[26056] <= 32'b00000000010100010010000000100011;
ROM[26057] <= 32'b00000000010000010000000100010011;
ROM[26058] <= 32'b00000000011000010010000000100011;
ROM[26059] <= 32'b00000000010000010000000100010011;
ROM[26060] <= 32'b00000001010000000000001110010011;
ROM[26061] <= 32'b00000000100000111000001110010011;
ROM[26062] <= 32'b01000000011100010000001110110011;
ROM[26063] <= 32'b00000000011100000000001000110011;
ROM[26064] <= 32'b00000000001000000000000110110011;
ROM[26065] <= 32'b01000110100000010000000011101111;
ROM[26066] <= 32'b00000111010000000000001110010011;
ROM[26067] <= 32'b00000000011100010010000000100011;
ROM[26068] <= 32'b00000000010000010000000100010011;
ROM[26069] <= 32'b00000000000000011001001110110111;
ROM[26070] <= 32'b01111010000000111000001110010011;
ROM[26071] <= 32'b00000000111000111000001110110011;
ROM[26072] <= 32'b00000000011100010010000000100011;
ROM[26073] <= 32'b00000000010000010000000100010011;
ROM[26074] <= 32'b00000000001100010010000000100011;
ROM[26075] <= 32'b00000000010000010000000100010011;
ROM[26076] <= 32'b00000000010000010010000000100011;
ROM[26077] <= 32'b00000000010000010000000100010011;
ROM[26078] <= 32'b00000000010100010010000000100011;
ROM[26079] <= 32'b00000000010000010000000100010011;
ROM[26080] <= 32'b00000000011000010010000000100011;
ROM[26081] <= 32'b00000000010000010000000100010011;
ROM[26082] <= 32'b00000001010000000000001110010011;
ROM[26083] <= 32'b00000000100000111000001110010011;
ROM[26084] <= 32'b01000000011100010000001110110011;
ROM[26085] <= 32'b00000000011100000000001000110011;
ROM[26086] <= 32'b00000000001000000000000110110011;
ROM[26087] <= 32'b01000001000000010000000011101111;
ROM[26088] <= 32'b00000110100000000000001110010011;
ROM[26089] <= 32'b00000000011100010010000000100011;
ROM[26090] <= 32'b00000000010000010000000100010011;
ROM[26091] <= 32'b00000000000000011001001110110111;
ROM[26092] <= 32'b01111111100000111000001110010011;
ROM[26093] <= 32'b00000000111000111000001110110011;
ROM[26094] <= 32'b00000000011100010010000000100011;
ROM[26095] <= 32'b00000000010000010000000100010011;
ROM[26096] <= 32'b00000000001100010010000000100011;
ROM[26097] <= 32'b00000000010000010000000100010011;
ROM[26098] <= 32'b00000000010000010010000000100011;
ROM[26099] <= 32'b00000000010000010000000100010011;
ROM[26100] <= 32'b00000000010100010010000000100011;
ROM[26101] <= 32'b00000000010000010000000100010011;
ROM[26102] <= 32'b00000000011000010010000000100011;
ROM[26103] <= 32'b00000000010000010000000100010011;
ROM[26104] <= 32'b00000001010000000000001110010011;
ROM[26105] <= 32'b00000000100000111000001110010011;
ROM[26106] <= 32'b01000000011100010000001110110011;
ROM[26107] <= 32'b00000000011100000000001000110011;
ROM[26108] <= 32'b00000000001000000000000110110011;
ROM[26109] <= 32'b00111011100000010000000011101111;
ROM[26110] <= 32'b00000110010100000000001110010011;
ROM[26111] <= 32'b00000000011100010010000000100011;
ROM[26112] <= 32'b00000000010000010000000100010011;
ROM[26113] <= 32'b00000000000000011010001110110111;
ROM[26114] <= 32'b10000101000000111000001110010011;
ROM[26115] <= 32'b00000000111000111000001110110011;
ROM[26116] <= 32'b00000000011100010010000000100011;
ROM[26117] <= 32'b00000000010000010000000100010011;
ROM[26118] <= 32'b00000000001100010010000000100011;
ROM[26119] <= 32'b00000000010000010000000100010011;
ROM[26120] <= 32'b00000000010000010010000000100011;
ROM[26121] <= 32'b00000000010000010000000100010011;
ROM[26122] <= 32'b00000000010100010010000000100011;
ROM[26123] <= 32'b00000000010000010000000100010011;
ROM[26124] <= 32'b00000000011000010010000000100011;
ROM[26125] <= 32'b00000000010000010000000100010011;
ROM[26126] <= 32'b00000001010000000000001110010011;
ROM[26127] <= 32'b00000000100000111000001110010011;
ROM[26128] <= 32'b01000000011100010000001110110011;
ROM[26129] <= 32'b00000000011100000000001000110011;
ROM[26130] <= 32'b00000000001000000000000110110011;
ROM[26131] <= 32'b00110110000000010000000011101111;
ROM[26132] <= 32'b00000010000000000000001110010011;
ROM[26133] <= 32'b00000000011100010010000000100011;
ROM[26134] <= 32'b00000000010000010000000100010011;
ROM[26135] <= 32'b00000000000000011010001110110111;
ROM[26136] <= 32'b10001010100000111000001110010011;
ROM[26137] <= 32'b00000000111000111000001110110011;
ROM[26138] <= 32'b00000000011100010010000000100011;
ROM[26139] <= 32'b00000000010000010000000100010011;
ROM[26140] <= 32'b00000000001100010010000000100011;
ROM[26141] <= 32'b00000000010000010000000100010011;
ROM[26142] <= 32'b00000000010000010010000000100011;
ROM[26143] <= 32'b00000000010000010000000100010011;
ROM[26144] <= 32'b00000000010100010010000000100011;
ROM[26145] <= 32'b00000000010000010000000100010011;
ROM[26146] <= 32'b00000000011000010010000000100011;
ROM[26147] <= 32'b00000000010000010000000100010011;
ROM[26148] <= 32'b00000001010000000000001110010011;
ROM[26149] <= 32'b00000000100000111000001110010011;
ROM[26150] <= 32'b01000000011100010000001110110011;
ROM[26151] <= 32'b00000000011100000000001000110011;
ROM[26152] <= 32'b00000000001000000000000110110011;
ROM[26153] <= 32'b00110000100000010000000011101111;
ROM[26154] <= 32'b00000110000100000000001110010011;
ROM[26155] <= 32'b00000000011100010010000000100011;
ROM[26156] <= 32'b00000000010000010000000100010011;
ROM[26157] <= 32'b00000000000000011010001110110111;
ROM[26158] <= 32'b10010000000000111000001110010011;
ROM[26159] <= 32'b00000000111000111000001110110011;
ROM[26160] <= 32'b00000000011100010010000000100011;
ROM[26161] <= 32'b00000000010000010000000100010011;
ROM[26162] <= 32'b00000000001100010010000000100011;
ROM[26163] <= 32'b00000000010000010000000100010011;
ROM[26164] <= 32'b00000000010000010010000000100011;
ROM[26165] <= 32'b00000000010000010000000100010011;
ROM[26166] <= 32'b00000000010100010010000000100011;
ROM[26167] <= 32'b00000000010000010000000100010011;
ROM[26168] <= 32'b00000000011000010010000000100011;
ROM[26169] <= 32'b00000000010000010000000100010011;
ROM[26170] <= 32'b00000001010000000000001110010011;
ROM[26171] <= 32'b00000000100000111000001110010011;
ROM[26172] <= 32'b01000000011100010000001110110011;
ROM[26173] <= 32'b00000000011100000000001000110011;
ROM[26174] <= 32'b00000000001000000000000110110011;
ROM[26175] <= 32'b00101011000000010000000011101111;
ROM[26176] <= 32'b00000111001000000000001110010011;
ROM[26177] <= 32'b00000000011100010010000000100011;
ROM[26178] <= 32'b00000000010000010000000100010011;
ROM[26179] <= 32'b00000000000000011010001110110111;
ROM[26180] <= 32'b10010101100000111000001110010011;
ROM[26181] <= 32'b00000000111000111000001110110011;
ROM[26182] <= 32'b00000000011100010010000000100011;
ROM[26183] <= 32'b00000000010000010000000100010011;
ROM[26184] <= 32'b00000000001100010010000000100011;
ROM[26185] <= 32'b00000000010000010000000100010011;
ROM[26186] <= 32'b00000000010000010010000000100011;
ROM[26187] <= 32'b00000000010000010000000100010011;
ROM[26188] <= 32'b00000000010100010010000000100011;
ROM[26189] <= 32'b00000000010000010000000100010011;
ROM[26190] <= 32'b00000000011000010010000000100011;
ROM[26191] <= 32'b00000000010000010000000100010011;
ROM[26192] <= 32'b00000001010000000000001110010011;
ROM[26193] <= 32'b00000000100000111000001110010011;
ROM[26194] <= 32'b01000000011100010000001110110011;
ROM[26195] <= 32'b00000000011100000000001000110011;
ROM[26196] <= 32'b00000000001000000000000110110011;
ROM[26197] <= 32'b00100101100000010000000011101111;
ROM[26198] <= 32'b00000111001000000000001110010011;
ROM[26199] <= 32'b00000000011100010010000000100011;
ROM[26200] <= 32'b00000000010000010000000100010011;
ROM[26201] <= 32'b00000000000000011010001110110111;
ROM[26202] <= 32'b10011011000000111000001110010011;
ROM[26203] <= 32'b00000000111000111000001110110011;
ROM[26204] <= 32'b00000000011100010010000000100011;
ROM[26205] <= 32'b00000000010000010000000100010011;
ROM[26206] <= 32'b00000000001100010010000000100011;
ROM[26207] <= 32'b00000000010000010000000100010011;
ROM[26208] <= 32'b00000000010000010010000000100011;
ROM[26209] <= 32'b00000000010000010000000100010011;
ROM[26210] <= 32'b00000000010100010010000000100011;
ROM[26211] <= 32'b00000000010000010000000100010011;
ROM[26212] <= 32'b00000000011000010010000000100011;
ROM[26213] <= 32'b00000000010000010000000100010011;
ROM[26214] <= 32'b00000001010000000000001110010011;
ROM[26215] <= 32'b00000000100000111000001110010011;
ROM[26216] <= 32'b01000000011100010000001110110011;
ROM[26217] <= 32'b00000000011100000000001000110011;
ROM[26218] <= 32'b00000000001000000000000110110011;
ROM[26219] <= 32'b00100000000000010000000011101111;
ROM[26220] <= 32'b00000110000100000000001110010011;
ROM[26221] <= 32'b00000000011100010010000000100011;
ROM[26222] <= 32'b00000000010000010000000100010011;
ROM[26223] <= 32'b00000000000000011010001110110111;
ROM[26224] <= 32'b10100000100000111000001110010011;
ROM[26225] <= 32'b00000000111000111000001110110011;
ROM[26226] <= 32'b00000000011100010010000000100011;
ROM[26227] <= 32'b00000000010000010000000100010011;
ROM[26228] <= 32'b00000000001100010010000000100011;
ROM[26229] <= 32'b00000000010000010000000100010011;
ROM[26230] <= 32'b00000000010000010010000000100011;
ROM[26231] <= 32'b00000000010000010000000100010011;
ROM[26232] <= 32'b00000000010100010010000000100011;
ROM[26233] <= 32'b00000000010000010000000100010011;
ROM[26234] <= 32'b00000000011000010010000000100011;
ROM[26235] <= 32'b00000000010000010000000100010011;
ROM[26236] <= 32'b00000001010000000000001110010011;
ROM[26237] <= 32'b00000000100000111000001110010011;
ROM[26238] <= 32'b01000000011100010000001110110011;
ROM[26239] <= 32'b00000000011100000000001000110011;
ROM[26240] <= 32'b00000000001000000000000110110011;
ROM[26241] <= 32'b00011010100000010000000011101111;
ROM[26242] <= 32'b00000111100100000000001110010011;
ROM[26243] <= 32'b00000000011100010010000000100011;
ROM[26244] <= 32'b00000000010000010000000100010011;
ROM[26245] <= 32'b00000000000000011010001110110111;
ROM[26246] <= 32'b10100110000000111000001110010011;
ROM[26247] <= 32'b00000000111000111000001110110011;
ROM[26248] <= 32'b00000000011100010010000000100011;
ROM[26249] <= 32'b00000000010000010000000100010011;
ROM[26250] <= 32'b00000000001100010010000000100011;
ROM[26251] <= 32'b00000000010000010000000100010011;
ROM[26252] <= 32'b00000000010000010010000000100011;
ROM[26253] <= 32'b00000000010000010000000100010011;
ROM[26254] <= 32'b00000000010100010010000000100011;
ROM[26255] <= 32'b00000000010000010000000100010011;
ROM[26256] <= 32'b00000000011000010010000000100011;
ROM[26257] <= 32'b00000000010000010000000100010011;
ROM[26258] <= 32'b00000001010000000000001110010011;
ROM[26259] <= 32'b00000000100000111000001110010011;
ROM[26260] <= 32'b01000000011100010000001110110011;
ROM[26261] <= 32'b00000000011100000000001000110011;
ROM[26262] <= 32'b00000000001000000000000110110011;
ROM[26263] <= 32'b00010101000000010000000011101111;
ROM[26264] <= 32'b00000011101000000000001110010011;
ROM[26265] <= 32'b00000000011100010010000000100011;
ROM[26266] <= 32'b00000000010000010000000100010011;
ROM[26267] <= 32'b00000000000000011010001110110111;
ROM[26268] <= 32'b10101011100000111000001110010011;
ROM[26269] <= 32'b00000000111000111000001110110011;
ROM[26270] <= 32'b00000000011100010010000000100011;
ROM[26271] <= 32'b00000000010000010000000100010011;
ROM[26272] <= 32'b00000000001100010010000000100011;
ROM[26273] <= 32'b00000000010000010000000100010011;
ROM[26274] <= 32'b00000000010000010010000000100011;
ROM[26275] <= 32'b00000000010000010000000100010011;
ROM[26276] <= 32'b00000000010100010010000000100011;
ROM[26277] <= 32'b00000000010000010000000100010011;
ROM[26278] <= 32'b00000000011000010010000000100011;
ROM[26279] <= 32'b00000000010000010000000100010011;
ROM[26280] <= 32'b00000001010000000000001110010011;
ROM[26281] <= 32'b00000000100000111000001110010011;
ROM[26282] <= 32'b01000000011100010000001110110011;
ROM[26283] <= 32'b00000000011100000000001000110011;
ROM[26284] <= 32'b00000000001000000000000110110011;
ROM[26285] <= 32'b00001111100000010000000011101111;
ROM[26286] <= 32'b00000010000000000000001110010011;
ROM[26287] <= 32'b00000000011100010010000000100011;
ROM[26288] <= 32'b00000000010000010000000100010011;
ROM[26289] <= 32'b00000000000000011010001110110111;
ROM[26290] <= 32'b10110001000000111000001110010011;
ROM[26291] <= 32'b00000000111000111000001110110011;
ROM[26292] <= 32'b00000000011100010010000000100011;
ROM[26293] <= 32'b00000000010000010000000100010011;
ROM[26294] <= 32'b00000000001100010010000000100011;
ROM[26295] <= 32'b00000000010000010000000100010011;
ROM[26296] <= 32'b00000000010000010010000000100011;
ROM[26297] <= 32'b00000000010000010000000100010011;
ROM[26298] <= 32'b00000000010100010010000000100011;
ROM[26299] <= 32'b00000000010000010000000100010011;
ROM[26300] <= 32'b00000000011000010010000000100011;
ROM[26301] <= 32'b00000000010000010000000100010011;
ROM[26302] <= 32'b00000001010000000000001110010011;
ROM[26303] <= 32'b00000000100000111000001110010011;
ROM[26304] <= 32'b01000000011100010000001110110011;
ROM[26305] <= 32'b00000000011100000000001000110011;
ROM[26306] <= 32'b00000000001000000000000110110011;
ROM[26307] <= 32'b00001010000000010000000011101111;
ROM[26308] <= 32'b00000000000000011010001110110111;
ROM[26309] <= 32'b10110101110000111000001110010011;
ROM[26310] <= 32'b00000000111000111000001110110011;
ROM[26311] <= 32'b00000000011100010010000000100011;
ROM[26312] <= 32'b00000000010000010000000100010011;
ROM[26313] <= 32'b00000000001100010010000000100011;
ROM[26314] <= 32'b00000000010000010000000100010011;
ROM[26315] <= 32'b00000000010000010010000000100011;
ROM[26316] <= 32'b00000000010000010000000100010011;
ROM[26317] <= 32'b00000000010100010010000000100011;
ROM[26318] <= 32'b00000000010000010000000100010011;
ROM[26319] <= 32'b00000000011000010010000000100011;
ROM[26320] <= 32'b00000000010000010000000100010011;
ROM[26321] <= 32'b00000001010000000000001110010011;
ROM[26322] <= 32'b00000000010000111000001110010011;
ROM[26323] <= 32'b01000000011100010000001110110011;
ROM[26324] <= 32'b00000000011100000000001000110011;
ROM[26325] <= 32'b00000000001000000000000110110011;
ROM[26326] <= 32'b11000001000011111101000011101111;
ROM[26327] <= 32'b11111111110000010000000100010011;
ROM[26328] <= 32'b00000000000000010010001110000011;
ROM[26329] <= 32'b00000000011101100010000000100011;
ROM[26330] <= 32'b00000000000000011010001110110111;
ROM[26331] <= 32'b10111011010000111000001110010011;
ROM[26332] <= 32'b00000000111000111000001110110011;
ROM[26333] <= 32'b00000000011100010010000000100011;
ROM[26334] <= 32'b00000000010000010000000100010011;
ROM[26335] <= 32'b00000000001100010010000000100011;
ROM[26336] <= 32'b00000000010000010000000100010011;
ROM[26337] <= 32'b00000000010000010010000000100011;
ROM[26338] <= 32'b00000000010000010000000100010011;
ROM[26339] <= 32'b00000000010100010010000000100011;
ROM[26340] <= 32'b00000000010000010000000100010011;
ROM[26341] <= 32'b00000000011000010010000000100011;
ROM[26342] <= 32'b00000000010000010000000100010011;
ROM[26343] <= 32'b00000001010000000000001110010011;
ROM[26344] <= 32'b00000000000000111000001110010011;
ROM[26345] <= 32'b01000000011100010000001110110011;
ROM[26346] <= 32'b00000000011100000000001000110011;
ROM[26347] <= 32'b00000000001000000000000110110011;
ROM[26348] <= 32'b11111011100011111101000011101111;
ROM[26349] <= 32'b11111111110000010000000100010011;
ROM[26350] <= 32'b00000000000000010010001110000011;
ROM[26351] <= 32'b00000000011101100010000000100011;
ROM[26352] <= 32'b00000000000000000000001110010011;
ROM[26353] <= 32'b00000000011100010010000000100011;
ROM[26354] <= 32'b00000000010000010000000100010011;
ROM[26355] <= 32'b11111111110000010000000100010011;
ROM[26356] <= 32'b00000000000000010010001110000011;
ROM[26357] <= 32'b00000000011100011010010000100011;
ROM[26358] <= 32'b00000000100000011010001110000011;
ROM[26359] <= 32'b00000000011100010010000000100011;
ROM[26360] <= 32'b00000000010000010000000100010011;
ROM[26361] <= 32'b00000000010000011010001110000011;
ROM[26362] <= 32'b00000000011100010010000000100011;
ROM[26363] <= 32'b00000000010000010000000100010011;
ROM[26364] <= 32'b11111111110000010000000100010011;
ROM[26365] <= 32'b00000000000000010010001110000011;
ROM[26366] <= 32'b11111111110000010000000100010011;
ROM[26367] <= 32'b00000000000000010010010000000011;
ROM[26368] <= 32'b00000000011101000010001110110011;
ROM[26369] <= 32'b00000000011100010010000000100011;
ROM[26370] <= 32'b00000000010000010000000100010011;
ROM[26371] <= 32'b11111111110000010000000100010011;
ROM[26372] <= 32'b00000000000000010010001110000011;
ROM[26373] <= 32'b01000000011100000000001110110011;
ROM[26374] <= 32'b00000000000100111000001110010011;
ROM[26375] <= 32'b00000000011100010010000000100011;
ROM[26376] <= 32'b00000000010000010000000100010011;
ROM[26377] <= 32'b11111111110000010000000100010011;
ROM[26378] <= 32'b00000000000000010010001110000011;
ROM[26379] <= 32'b00000000000000111000101001100011;
ROM[26380] <= 32'b00000000000000011010001110110111;
ROM[26381] <= 32'b11011101000000111000001110010011;
ROM[26382] <= 32'b00000000111000111000001110110011;
ROM[26383] <= 32'b00000000000000111000000011100111;
ROM[26384] <= 32'b00000000000000000000001110010011;
ROM[26385] <= 32'b00000000011100010010000000100011;
ROM[26386] <= 32'b00000000010000010000000100010011;
ROM[26387] <= 32'b00000000000000011010001110110111;
ROM[26388] <= 32'b11001001100000111000001110010011;
ROM[26389] <= 32'b00000000111000111000001110110011;
ROM[26390] <= 32'b00000000011100010010000000100011;
ROM[26391] <= 32'b00000000010000010000000100010011;
ROM[26392] <= 32'b00000000001100010010000000100011;
ROM[26393] <= 32'b00000000010000010000000100010011;
ROM[26394] <= 32'b00000000010000010010000000100011;
ROM[26395] <= 32'b00000000010000010000000100010011;
ROM[26396] <= 32'b00000000010100010010000000100011;
ROM[26397] <= 32'b00000000010000010000000100010011;
ROM[26398] <= 32'b00000000011000010010000000100011;
ROM[26399] <= 32'b00000000010000010000000100010011;
ROM[26400] <= 32'b00000001010000000000001110010011;
ROM[26401] <= 32'b00000000010000111000001110010011;
ROM[26402] <= 32'b01000000011100010000001110110011;
ROM[26403] <= 32'b00000000011100000000001000110011;
ROM[26404] <= 32'b00000000001000000000000110110011;
ROM[26405] <= 32'b00101010100100001111000011101111;
ROM[26406] <= 32'b00000000000000011010001110110111;
ROM[26407] <= 32'b11001110010000111000001110010011;
ROM[26408] <= 32'b00000000111000111000001110110011;
ROM[26409] <= 32'b00000000011100010010000000100011;
ROM[26410] <= 32'b00000000010000010000000100010011;
ROM[26411] <= 32'b00000000001100010010000000100011;
ROM[26412] <= 32'b00000000010000010000000100010011;
ROM[26413] <= 32'b00000000010000010010000000100011;
ROM[26414] <= 32'b00000000010000010000000100010011;
ROM[26415] <= 32'b00000000010100010010000000100011;
ROM[26416] <= 32'b00000000010000010000000100010011;
ROM[26417] <= 32'b00000000011000010010000000100011;
ROM[26418] <= 32'b00000000010000010000000100010011;
ROM[26419] <= 32'b00000001010000000000001110010011;
ROM[26420] <= 32'b00000000010000111000001110010011;
ROM[26421] <= 32'b01000000011100010000001110110011;
ROM[26422] <= 32'b00000000011100000000001000110011;
ROM[26423] <= 32'b00000000001000000000000110110011;
ROM[26424] <= 32'b10111110100011110100000011101111;
ROM[26425] <= 32'b00000000000000011010001110000011;
ROM[26426] <= 32'b00000000011100010010000000100011;
ROM[26427] <= 32'b00000000010000010000000100010011;
ROM[26428] <= 32'b00000000100000011010001110000011;
ROM[26429] <= 32'b00000000011100010010000000100011;
ROM[26430] <= 32'b00000000010000010000000100010011;
ROM[26431] <= 32'b00000000010000000000001110010011;
ROM[26432] <= 32'b00000000011100010010000000100011;
ROM[26433] <= 32'b00000000010000010000000100010011;
ROM[26434] <= 32'b00000000000000011010001110110111;
ROM[26435] <= 32'b11010101010000111000001110010011;
ROM[26436] <= 32'b00000000111000111000001110110011;
ROM[26437] <= 32'b00000000011100010010000000100011;
ROM[26438] <= 32'b00000000010000010000000100010011;
ROM[26439] <= 32'b00000000001100010010000000100011;
ROM[26440] <= 32'b00000000010000010000000100010011;
ROM[26441] <= 32'b00000000010000010010000000100011;
ROM[26442] <= 32'b00000000010000010000000100010011;
ROM[26443] <= 32'b00000000010100010010000000100011;
ROM[26444] <= 32'b00000000010000010000000100010011;
ROM[26445] <= 32'b00000000011000010010000000100011;
ROM[26446] <= 32'b00000000010000010000000100010011;
ROM[26447] <= 32'b00000001010000000000001110010011;
ROM[26448] <= 32'b00000000100000111000001110010011;
ROM[26449] <= 32'b01000000011100010000001110110011;
ROM[26450] <= 32'b00000000011100000000001000110011;
ROM[26451] <= 32'b00000000001000000000000110110011;
ROM[26452] <= 32'b10101101110111110111000011101111;
ROM[26453] <= 32'b11111111110000010000000100010011;
ROM[26454] <= 32'b00000000000000010010001110000011;
ROM[26455] <= 32'b11111111110000010000000100010011;
ROM[26456] <= 32'b00000000000000010010010000000011;
ROM[26457] <= 32'b00000000011101000000001110110011;
ROM[26458] <= 32'b00000000011100010010000000100011;
ROM[26459] <= 32'b00000000010000010000000100010011;
ROM[26460] <= 32'b11111111110000010000000100010011;
ROM[26461] <= 32'b00000000000000010010001110000011;
ROM[26462] <= 32'b00000000000000111000001100010011;
ROM[26463] <= 32'b11111111110000010000000100010011;
ROM[26464] <= 32'b00000000000000010010001110000011;
ROM[26465] <= 32'b00000000110100110000010000110011;
ROM[26466] <= 32'b00000000011101000010000000100011;
ROM[26467] <= 32'b00000000100000011010001110000011;
ROM[26468] <= 32'b00000000011100010010000000100011;
ROM[26469] <= 32'b00000000010000010000000100010011;
ROM[26470] <= 32'b00000000000100000000001110010011;
ROM[26471] <= 32'b00000000011100010010000000100011;
ROM[26472] <= 32'b00000000010000010000000100010011;
ROM[26473] <= 32'b11111111110000010000000100010011;
ROM[26474] <= 32'b00000000000000010010001110000011;
ROM[26475] <= 32'b11111111110000010000000100010011;
ROM[26476] <= 32'b00000000000000010010010000000011;
ROM[26477] <= 32'b00000000011101000000001110110011;
ROM[26478] <= 32'b00000000011100010010000000100011;
ROM[26479] <= 32'b00000000010000010000000100010011;
ROM[26480] <= 32'b11111111110000010000000100010011;
ROM[26481] <= 32'b00000000000000010010001110000011;
ROM[26482] <= 32'b00000000011100011010010000100011;
ROM[26483] <= 32'b11100000110111111111000011101111;
ROM[26484] <= 32'b00000000000000011010001110000011;
ROM[26485] <= 32'b00000000011100010010000000100011;
ROM[26486] <= 32'b00000000010000010000000100010011;
ROM[26487] <= 32'b00000000000000000000001110010011;
ROM[26488] <= 32'b00000000011100010010000000100011;
ROM[26489] <= 32'b00000000010000010000000100010011;
ROM[26490] <= 32'b00000000010000011010001110000011;
ROM[26491] <= 32'b00000000011100010010000000100011;
ROM[26492] <= 32'b00000000010000010000000100010011;
ROM[26493] <= 32'b00000000000100000000001110010011;
ROM[26494] <= 32'b00000000011100010010000000100011;
ROM[26495] <= 32'b00000000010000010000000100010011;
ROM[26496] <= 32'b11111111110000010000000100010011;
ROM[26497] <= 32'b00000000000000010010001110000011;
ROM[26498] <= 32'b11111111110000010000000100010011;
ROM[26499] <= 32'b00000000000000010010010000000011;
ROM[26500] <= 32'b01000000011101000000001110110011;
ROM[26501] <= 32'b00000000011100010010000000100011;
ROM[26502] <= 32'b00000000010000010000000100010011;
ROM[26503] <= 32'b00000000000000011010001110110111;
ROM[26504] <= 32'b11100110100000111000001110010011;
ROM[26505] <= 32'b00000000111000111000001110110011;
ROM[26506] <= 32'b00000000011100010010000000100011;
ROM[26507] <= 32'b00000000010000010000000100010011;
ROM[26508] <= 32'b00000000001100010010000000100011;
ROM[26509] <= 32'b00000000010000010000000100010011;
ROM[26510] <= 32'b00000000010000010010000000100011;
ROM[26511] <= 32'b00000000010000010000000100010011;
ROM[26512] <= 32'b00000000010100010010000000100011;
ROM[26513] <= 32'b00000000010000010000000100010011;
ROM[26514] <= 32'b00000000011000010010000000100011;
ROM[26515] <= 32'b00000000010000010000000100010011;
ROM[26516] <= 32'b00000001010000000000001110010011;
ROM[26517] <= 32'b00000000110000111000001110010011;
ROM[26518] <= 32'b01000000011100010000001110110011;
ROM[26519] <= 32'b00000000011100000000001000110011;
ROM[26520] <= 32'b00000000001000000000000110110011;
ROM[26521] <= 32'b01010001010100000000000011101111;
ROM[26522] <= 32'b11111111110000010000000100010011;
ROM[26523] <= 32'b00000000000000010010001110000011;
ROM[26524] <= 32'b00000000011101100010000000100011;
ROM[26525] <= 32'b00000001010100000000001110010011;
ROM[26526] <= 32'b00000000011100010010000000100011;
ROM[26527] <= 32'b00000000010000010000000100010011;
ROM[26528] <= 32'b00000000000000011010001110110111;
ROM[26529] <= 32'b11101100110000111000001110010011;
ROM[26530] <= 32'b00000000111000111000001110110011;
ROM[26531] <= 32'b00000000011100010010000000100011;
ROM[26532] <= 32'b00000000010000010000000100010011;
ROM[26533] <= 32'b00000000001100010010000000100011;
ROM[26534] <= 32'b00000000010000010000000100010011;
ROM[26535] <= 32'b00000000010000010010000000100011;
ROM[26536] <= 32'b00000000010000010000000100010011;
ROM[26537] <= 32'b00000000010100010010000000100011;
ROM[26538] <= 32'b00000000010000010000000100010011;
ROM[26539] <= 32'b00000000011000010010000000100011;
ROM[26540] <= 32'b00000000010000010000000100010011;
ROM[26541] <= 32'b00000001010000000000001110010011;
ROM[26542] <= 32'b00000000010000111000001110010011;
ROM[26543] <= 32'b01000000011100010000001110110011;
ROM[26544] <= 32'b00000000011100000000001000110011;
ROM[26545] <= 32'b00000000001000000000000110110011;
ROM[26546] <= 32'b00000111010100001111000011101111;
ROM[26547] <= 32'b00000101010000000000001110010011;
ROM[26548] <= 32'b00000000011100010010000000100011;
ROM[26549] <= 32'b00000000010000010000000100010011;
ROM[26550] <= 32'b00000000000000011010001110110111;
ROM[26551] <= 32'b11110010010000111000001110010011;
ROM[26552] <= 32'b00000000111000111000001110110011;
ROM[26553] <= 32'b00000000011100010010000000100011;
ROM[26554] <= 32'b00000000010000010000000100010011;
ROM[26555] <= 32'b00000000001100010010000000100011;
ROM[26556] <= 32'b00000000010000010000000100010011;
ROM[26557] <= 32'b00000000010000010010000000100011;
ROM[26558] <= 32'b00000000010000010000000100010011;
ROM[26559] <= 32'b00000000010100010010000000100011;
ROM[26560] <= 32'b00000000010000010000000100010011;
ROM[26561] <= 32'b00000000011000010010000000100011;
ROM[26562] <= 32'b00000000010000010000000100010011;
ROM[26563] <= 32'b00000001010000000000001110010011;
ROM[26564] <= 32'b00000000100000111000001110010011;
ROM[26565] <= 32'b01000000011100010000001110110011;
ROM[26566] <= 32'b00000000011100000000001000110011;
ROM[26567] <= 32'b00000000001000000000000110110011;
ROM[26568] <= 32'b01001000110100001111000011101111;
ROM[26569] <= 32'b00000110100000000000001110010011;
ROM[26570] <= 32'b00000000011100010010000000100011;
ROM[26571] <= 32'b00000000010000010000000100010011;
ROM[26572] <= 32'b00000000000000011010001110110111;
ROM[26573] <= 32'b11110111110000111000001110010011;
ROM[26574] <= 32'b00000000111000111000001110110011;
ROM[26575] <= 32'b00000000011100010010000000100011;
ROM[26576] <= 32'b00000000010000010000000100010011;
ROM[26577] <= 32'b00000000001100010010000000100011;
ROM[26578] <= 32'b00000000010000010000000100010011;
ROM[26579] <= 32'b00000000010000010010000000100011;
ROM[26580] <= 32'b00000000010000010000000100010011;
ROM[26581] <= 32'b00000000010100010010000000100011;
ROM[26582] <= 32'b00000000010000010000000100010011;
ROM[26583] <= 32'b00000000011000010010000000100011;
ROM[26584] <= 32'b00000000010000010000000100010011;
ROM[26585] <= 32'b00000001010000000000001110010011;
ROM[26586] <= 32'b00000000100000111000001110010011;
ROM[26587] <= 32'b01000000011100010000001110110011;
ROM[26588] <= 32'b00000000011100000000001000110011;
ROM[26589] <= 32'b00000000001000000000000110110011;
ROM[26590] <= 32'b01000011010100001111000011101111;
ROM[26591] <= 32'b00000110010100000000001110010011;
ROM[26592] <= 32'b00000000011100010010000000100011;
ROM[26593] <= 32'b00000000010000010000000100010011;
ROM[26594] <= 32'b00000000000000011010001110110111;
ROM[26595] <= 32'b11111101010000111000001110010011;
ROM[26596] <= 32'b00000000111000111000001110110011;
ROM[26597] <= 32'b00000000011100010010000000100011;
ROM[26598] <= 32'b00000000010000010000000100010011;
ROM[26599] <= 32'b00000000001100010010000000100011;
ROM[26600] <= 32'b00000000010000010000000100010011;
ROM[26601] <= 32'b00000000010000010010000000100011;
ROM[26602] <= 32'b00000000010000010000000100010011;
ROM[26603] <= 32'b00000000010100010010000000100011;
ROM[26604] <= 32'b00000000010000010000000100010011;
ROM[26605] <= 32'b00000000011000010010000000100011;
ROM[26606] <= 32'b00000000010000010000000100010011;
ROM[26607] <= 32'b00000001010000000000001110010011;
ROM[26608] <= 32'b00000000100000111000001110010011;
ROM[26609] <= 32'b01000000011100010000001110110011;
ROM[26610] <= 32'b00000000011100000000001000110011;
ROM[26611] <= 32'b00000000001000000000000110110011;
ROM[26612] <= 32'b00111101110100001111000011101111;
ROM[26613] <= 32'b00000010000000000000001110010011;
ROM[26614] <= 32'b00000000011100010010000000100011;
ROM[26615] <= 32'b00000000010000010000000100010011;
ROM[26616] <= 32'b00000000000000011010001110110111;
ROM[26617] <= 32'b00000010110000111000001110010011;
ROM[26618] <= 32'b00000000111000111000001110110011;
ROM[26619] <= 32'b00000000011100010010000000100011;
ROM[26620] <= 32'b00000000010000010000000100010011;
ROM[26621] <= 32'b00000000001100010010000000100011;
ROM[26622] <= 32'b00000000010000010000000100010011;
ROM[26623] <= 32'b00000000010000010010000000100011;
ROM[26624] <= 32'b00000000010000010000000100010011;
ROM[26625] <= 32'b00000000010100010010000000100011;
ROM[26626] <= 32'b00000000010000010000000100010011;
ROM[26627] <= 32'b00000000011000010010000000100011;
ROM[26628] <= 32'b00000000010000010000000100010011;
ROM[26629] <= 32'b00000001010000000000001110010011;
ROM[26630] <= 32'b00000000100000111000001110010011;
ROM[26631] <= 32'b01000000011100010000001110110011;
ROM[26632] <= 32'b00000000011100000000001000110011;
ROM[26633] <= 32'b00000000001000000000000110110011;
ROM[26634] <= 32'b00111000010100001111000011101111;
ROM[26635] <= 32'b00000111001100000000001110010011;
ROM[26636] <= 32'b00000000011100010010000000100011;
ROM[26637] <= 32'b00000000010000010000000100010011;
ROM[26638] <= 32'b00000000000000011010001110110111;
ROM[26639] <= 32'b00001000010000111000001110010011;
ROM[26640] <= 32'b00000000111000111000001110110011;
ROM[26641] <= 32'b00000000011100010010000000100011;
ROM[26642] <= 32'b00000000010000010000000100010011;
ROM[26643] <= 32'b00000000001100010010000000100011;
ROM[26644] <= 32'b00000000010000010000000100010011;
ROM[26645] <= 32'b00000000010000010010000000100011;
ROM[26646] <= 32'b00000000010000010000000100010011;
ROM[26647] <= 32'b00000000010100010010000000100011;
ROM[26648] <= 32'b00000000010000010000000100010011;
ROM[26649] <= 32'b00000000011000010010000000100011;
ROM[26650] <= 32'b00000000010000010000000100010011;
ROM[26651] <= 32'b00000001010000000000001110010011;
ROM[26652] <= 32'b00000000100000111000001110010011;
ROM[26653] <= 32'b01000000011100010000001110110011;
ROM[26654] <= 32'b00000000011100000000001000110011;
ROM[26655] <= 32'b00000000001000000000000110110011;
ROM[26656] <= 32'b00110010110100001111000011101111;
ROM[26657] <= 32'b00000110111100000000001110010011;
ROM[26658] <= 32'b00000000011100010010000000100011;
ROM[26659] <= 32'b00000000010000010000000100010011;
ROM[26660] <= 32'b00000000000000011010001110110111;
ROM[26661] <= 32'b00001101110000111000001110010011;
ROM[26662] <= 32'b00000000111000111000001110110011;
ROM[26663] <= 32'b00000000011100010010000000100011;
ROM[26664] <= 32'b00000000010000010000000100010011;
ROM[26665] <= 32'b00000000001100010010000000100011;
ROM[26666] <= 32'b00000000010000010000000100010011;
ROM[26667] <= 32'b00000000010000010010000000100011;
ROM[26668] <= 32'b00000000010000010000000100010011;
ROM[26669] <= 32'b00000000010100010010000000100011;
ROM[26670] <= 32'b00000000010000010000000100010011;
ROM[26671] <= 32'b00000000011000010010000000100011;
ROM[26672] <= 32'b00000000010000010000000100010011;
ROM[26673] <= 32'b00000001010000000000001110010011;
ROM[26674] <= 32'b00000000100000111000001110010011;
ROM[26675] <= 32'b01000000011100010000001110110011;
ROM[26676] <= 32'b00000000011100000000001000110011;
ROM[26677] <= 32'b00000000001000000000000110110011;
ROM[26678] <= 32'b00101101010100001111000011101111;
ROM[26679] <= 32'b00000111001000000000001110010011;
ROM[26680] <= 32'b00000000011100010010000000100011;
ROM[26681] <= 32'b00000000010000010000000100010011;
ROM[26682] <= 32'b00000000000000011010001110110111;
ROM[26683] <= 32'b00010011010000111000001110010011;
ROM[26684] <= 32'b00000000111000111000001110110011;
ROM[26685] <= 32'b00000000011100010010000000100011;
ROM[26686] <= 32'b00000000010000010000000100010011;
ROM[26687] <= 32'b00000000001100010010000000100011;
ROM[26688] <= 32'b00000000010000010000000100010011;
ROM[26689] <= 32'b00000000010000010010000000100011;
ROM[26690] <= 32'b00000000010000010000000100010011;
ROM[26691] <= 32'b00000000010100010010000000100011;
ROM[26692] <= 32'b00000000010000010000000100010011;
ROM[26693] <= 32'b00000000011000010010000000100011;
ROM[26694] <= 32'b00000000010000010000000100010011;
ROM[26695] <= 32'b00000001010000000000001110010011;
ROM[26696] <= 32'b00000000100000111000001110010011;
ROM[26697] <= 32'b01000000011100010000001110110011;
ROM[26698] <= 32'b00000000011100000000001000110011;
ROM[26699] <= 32'b00000000001000000000000110110011;
ROM[26700] <= 32'b00100111110100001111000011101111;
ROM[26701] <= 32'b00000111010000000000001110010011;
ROM[26702] <= 32'b00000000011100010010000000100011;
ROM[26703] <= 32'b00000000010000010000000100010011;
ROM[26704] <= 32'b00000000000000011010001110110111;
ROM[26705] <= 32'b00011000110000111000001110010011;
ROM[26706] <= 32'b00000000111000111000001110110011;
ROM[26707] <= 32'b00000000011100010010000000100011;
ROM[26708] <= 32'b00000000010000010000000100010011;
ROM[26709] <= 32'b00000000001100010010000000100011;
ROM[26710] <= 32'b00000000010000010000000100010011;
ROM[26711] <= 32'b00000000010000010010000000100011;
ROM[26712] <= 32'b00000000010000010000000100010011;
ROM[26713] <= 32'b00000000010100010010000000100011;
ROM[26714] <= 32'b00000000010000010000000100010011;
ROM[26715] <= 32'b00000000011000010010000000100011;
ROM[26716] <= 32'b00000000010000010000000100010011;
ROM[26717] <= 32'b00000001010000000000001110010011;
ROM[26718] <= 32'b00000000100000111000001110010011;
ROM[26719] <= 32'b01000000011100010000001110110011;
ROM[26720] <= 32'b00000000011100000000001000110011;
ROM[26721] <= 32'b00000000001000000000000110110011;
ROM[26722] <= 32'b00100010010100001111000011101111;
ROM[26723] <= 32'b00000110010100000000001110010011;
ROM[26724] <= 32'b00000000011100010010000000100011;
ROM[26725] <= 32'b00000000010000010000000100010011;
ROM[26726] <= 32'b00000000000000011010001110110111;
ROM[26727] <= 32'b00011110010000111000001110010011;
ROM[26728] <= 32'b00000000111000111000001110110011;
ROM[26729] <= 32'b00000000011100010010000000100011;
ROM[26730] <= 32'b00000000010000010000000100010011;
ROM[26731] <= 32'b00000000001100010010000000100011;
ROM[26732] <= 32'b00000000010000010000000100010011;
ROM[26733] <= 32'b00000000010000010010000000100011;
ROM[26734] <= 32'b00000000010000010000000100010011;
ROM[26735] <= 32'b00000000010100010010000000100011;
ROM[26736] <= 32'b00000000010000010000000100010011;
ROM[26737] <= 32'b00000000011000010010000000100011;
ROM[26738] <= 32'b00000000010000010000000100010011;
ROM[26739] <= 32'b00000001010000000000001110010011;
ROM[26740] <= 32'b00000000100000111000001110010011;
ROM[26741] <= 32'b01000000011100010000001110110011;
ROM[26742] <= 32'b00000000011100000000001000110011;
ROM[26743] <= 32'b00000000001000000000000110110011;
ROM[26744] <= 32'b00011100110100001111000011101111;
ROM[26745] <= 32'b00000110010000000000001110010011;
ROM[26746] <= 32'b00000000011100010010000000100011;
ROM[26747] <= 32'b00000000010000010000000100010011;
ROM[26748] <= 32'b00000000000000011010001110110111;
ROM[26749] <= 32'b00100011110000111000001110010011;
ROM[26750] <= 32'b00000000111000111000001110110011;
ROM[26751] <= 32'b00000000011100010010000000100011;
ROM[26752] <= 32'b00000000010000010000000100010011;
ROM[26753] <= 32'b00000000001100010010000000100011;
ROM[26754] <= 32'b00000000010000010000000100010011;
ROM[26755] <= 32'b00000000010000010010000000100011;
ROM[26756] <= 32'b00000000010000010000000100010011;
ROM[26757] <= 32'b00000000010100010010000000100011;
ROM[26758] <= 32'b00000000010000010000000100010011;
ROM[26759] <= 32'b00000000011000010010000000100011;
ROM[26760] <= 32'b00000000010000010000000100010011;
ROM[26761] <= 32'b00000001010000000000001110010011;
ROM[26762] <= 32'b00000000100000111000001110010011;
ROM[26763] <= 32'b01000000011100010000001110110011;
ROM[26764] <= 32'b00000000011100000000001000110011;
ROM[26765] <= 32'b00000000001000000000000110110011;
ROM[26766] <= 32'b00010111010100001111000011101111;
ROM[26767] <= 32'b00000010000000000000001110010011;
ROM[26768] <= 32'b00000000011100010010000000100011;
ROM[26769] <= 32'b00000000010000010000000100010011;
ROM[26770] <= 32'b00000000000000011010001110110111;
ROM[26771] <= 32'b00101001010000111000001110010011;
ROM[26772] <= 32'b00000000111000111000001110110011;
ROM[26773] <= 32'b00000000011100010010000000100011;
ROM[26774] <= 32'b00000000010000010000000100010011;
ROM[26775] <= 32'b00000000001100010010000000100011;
ROM[26776] <= 32'b00000000010000010000000100010011;
ROM[26777] <= 32'b00000000010000010010000000100011;
ROM[26778] <= 32'b00000000010000010000000100010011;
ROM[26779] <= 32'b00000000010100010010000000100011;
ROM[26780] <= 32'b00000000010000010000000100010011;
ROM[26781] <= 32'b00000000011000010010000000100011;
ROM[26782] <= 32'b00000000010000010000000100010011;
ROM[26783] <= 32'b00000001010000000000001110010011;
ROM[26784] <= 32'b00000000100000111000001110010011;
ROM[26785] <= 32'b01000000011100010000001110110011;
ROM[26786] <= 32'b00000000011100000000001000110011;
ROM[26787] <= 32'b00000000001000000000000110110011;
ROM[26788] <= 32'b00010001110100001111000011101111;
ROM[26789] <= 32'b00000110000100000000001110010011;
ROM[26790] <= 32'b00000000011100010010000000100011;
ROM[26791] <= 32'b00000000010000010000000100010011;
ROM[26792] <= 32'b00000000000000011010001110110111;
ROM[26793] <= 32'b00101110110000111000001110010011;
ROM[26794] <= 32'b00000000111000111000001110110011;
ROM[26795] <= 32'b00000000011100010010000000100011;
ROM[26796] <= 32'b00000000010000010000000100010011;
ROM[26797] <= 32'b00000000001100010010000000100011;
ROM[26798] <= 32'b00000000010000010000000100010011;
ROM[26799] <= 32'b00000000010000010010000000100011;
ROM[26800] <= 32'b00000000010000010000000100010011;
ROM[26801] <= 32'b00000000010100010010000000100011;
ROM[26802] <= 32'b00000000010000010000000100010011;
ROM[26803] <= 32'b00000000011000010010000000100011;
ROM[26804] <= 32'b00000000010000010000000100010011;
ROM[26805] <= 32'b00000001010000000000001110010011;
ROM[26806] <= 32'b00000000100000111000001110010011;
ROM[26807] <= 32'b01000000011100010000001110110011;
ROM[26808] <= 32'b00000000011100000000001000110011;
ROM[26809] <= 32'b00000000001000000000000110110011;
ROM[26810] <= 32'b00001100010100001111000011101111;
ROM[26811] <= 32'b00000111001000000000001110010011;
ROM[26812] <= 32'b00000000011100010010000000100011;
ROM[26813] <= 32'b00000000010000010000000100010011;
ROM[26814] <= 32'b00000000000000011010001110110111;
ROM[26815] <= 32'b00110100010000111000001110010011;
ROM[26816] <= 32'b00000000111000111000001110110011;
ROM[26817] <= 32'b00000000011100010010000000100011;
ROM[26818] <= 32'b00000000010000010000000100010011;
ROM[26819] <= 32'b00000000001100010010000000100011;
ROM[26820] <= 32'b00000000010000010000000100010011;
ROM[26821] <= 32'b00000000010000010010000000100011;
ROM[26822] <= 32'b00000000010000010000000100010011;
ROM[26823] <= 32'b00000000010100010010000000100011;
ROM[26824] <= 32'b00000000010000010000000100010011;
ROM[26825] <= 32'b00000000011000010010000000100011;
ROM[26826] <= 32'b00000000010000010000000100010011;
ROM[26827] <= 32'b00000001010000000000001110010011;
ROM[26828] <= 32'b00000000100000111000001110010011;
ROM[26829] <= 32'b01000000011100010000001110110011;
ROM[26830] <= 32'b00000000011100000000001000110011;
ROM[26831] <= 32'b00000000001000000000000110110011;
ROM[26832] <= 32'b00000110110100001111000011101111;
ROM[26833] <= 32'b00000111001000000000001110010011;
ROM[26834] <= 32'b00000000011100010010000000100011;
ROM[26835] <= 32'b00000000010000010000000100010011;
ROM[26836] <= 32'b00000000000000011010001110110111;
ROM[26837] <= 32'b00111001110000111000001110010011;
ROM[26838] <= 32'b00000000111000111000001110110011;
ROM[26839] <= 32'b00000000011100010010000000100011;
ROM[26840] <= 32'b00000000010000010000000100010011;
ROM[26841] <= 32'b00000000001100010010000000100011;
ROM[26842] <= 32'b00000000010000010000000100010011;
ROM[26843] <= 32'b00000000010000010010000000100011;
ROM[26844] <= 32'b00000000010000010000000100010011;
ROM[26845] <= 32'b00000000010100010010000000100011;
ROM[26846] <= 32'b00000000010000010000000100010011;
ROM[26847] <= 32'b00000000011000010010000000100011;
ROM[26848] <= 32'b00000000010000010000000100010011;
ROM[26849] <= 32'b00000001010000000000001110010011;
ROM[26850] <= 32'b00000000100000111000001110010011;
ROM[26851] <= 32'b01000000011100010000001110110011;
ROM[26852] <= 32'b00000000011100000000001000110011;
ROM[26853] <= 32'b00000000001000000000000110110011;
ROM[26854] <= 32'b00000001010100001111000011101111;
ROM[26855] <= 32'b00000110000100000000001110010011;
ROM[26856] <= 32'b00000000011100010010000000100011;
ROM[26857] <= 32'b00000000010000010000000100010011;
ROM[26858] <= 32'b00000000000000011010001110110111;
ROM[26859] <= 32'b00111111010000111000001110010011;
ROM[26860] <= 32'b00000000111000111000001110110011;
ROM[26861] <= 32'b00000000011100010010000000100011;
ROM[26862] <= 32'b00000000010000010000000100010011;
ROM[26863] <= 32'b00000000001100010010000000100011;
ROM[26864] <= 32'b00000000010000010000000100010011;
ROM[26865] <= 32'b00000000010000010010000000100011;
ROM[26866] <= 32'b00000000010000010000000100010011;
ROM[26867] <= 32'b00000000010100010010000000100011;
ROM[26868] <= 32'b00000000010000010000000100010011;
ROM[26869] <= 32'b00000000011000010010000000100011;
ROM[26870] <= 32'b00000000010000010000000100010011;
ROM[26871] <= 32'b00000001010000000000001110010011;
ROM[26872] <= 32'b00000000100000111000001110010011;
ROM[26873] <= 32'b01000000011100010000001110110011;
ROM[26874] <= 32'b00000000011100000000001000110011;
ROM[26875] <= 32'b00000000001000000000000110110011;
ROM[26876] <= 32'b01111011110000001111000011101111;
ROM[26877] <= 32'b00000111100100000000001110010011;
ROM[26878] <= 32'b00000000011100010010000000100011;
ROM[26879] <= 32'b00000000010000010000000100010011;
ROM[26880] <= 32'b00000000000000011010001110110111;
ROM[26881] <= 32'b01000100110000111000001110010011;
ROM[26882] <= 32'b00000000111000111000001110110011;
ROM[26883] <= 32'b00000000011100010010000000100011;
ROM[26884] <= 32'b00000000010000010000000100010011;
ROM[26885] <= 32'b00000000001100010010000000100011;
ROM[26886] <= 32'b00000000010000010000000100010011;
ROM[26887] <= 32'b00000000010000010010000000100011;
ROM[26888] <= 32'b00000000010000010000000100010011;
ROM[26889] <= 32'b00000000010100010010000000100011;
ROM[26890] <= 32'b00000000010000010000000100010011;
ROM[26891] <= 32'b00000000011000010010000000100011;
ROM[26892] <= 32'b00000000010000010000000100010011;
ROM[26893] <= 32'b00000001010000000000001110010011;
ROM[26894] <= 32'b00000000100000111000001110010011;
ROM[26895] <= 32'b01000000011100010000001110110011;
ROM[26896] <= 32'b00000000011100000000001000110011;
ROM[26897] <= 32'b00000000001000000000000110110011;
ROM[26898] <= 32'b01110110010000001111000011101111;
ROM[26899] <= 32'b00000010000000000000001110010011;
ROM[26900] <= 32'b00000000011100010010000000100011;
ROM[26901] <= 32'b00000000010000010000000100010011;
ROM[26902] <= 32'b00000000000000011010001110110111;
ROM[26903] <= 32'b01001010010000111000001110010011;
ROM[26904] <= 32'b00000000111000111000001110110011;
ROM[26905] <= 32'b00000000011100010010000000100011;
ROM[26906] <= 32'b00000000010000010000000100010011;
ROM[26907] <= 32'b00000000001100010010000000100011;
ROM[26908] <= 32'b00000000010000010000000100010011;
ROM[26909] <= 32'b00000000010000010010000000100011;
ROM[26910] <= 32'b00000000010000010000000100010011;
ROM[26911] <= 32'b00000000010100010010000000100011;
ROM[26912] <= 32'b00000000010000010000000100010011;
ROM[26913] <= 32'b00000000011000010010000000100011;
ROM[26914] <= 32'b00000000010000010000000100010011;
ROM[26915] <= 32'b00000001010000000000001110010011;
ROM[26916] <= 32'b00000000100000111000001110010011;
ROM[26917] <= 32'b01000000011100010000001110110011;
ROM[26918] <= 32'b00000000011100000000001000110011;
ROM[26919] <= 32'b00000000001000000000000110110011;
ROM[26920] <= 32'b01110000110000001111000011101111;
ROM[26921] <= 32'b00000110100100000000001110010011;
ROM[26922] <= 32'b00000000011100010010000000100011;
ROM[26923] <= 32'b00000000010000010000000100010011;
ROM[26924] <= 32'b00000000000000011010001110110111;
ROM[26925] <= 32'b01001111110000111000001110010011;
ROM[26926] <= 32'b00000000111000111000001110110011;
ROM[26927] <= 32'b00000000011100010010000000100011;
ROM[26928] <= 32'b00000000010000010000000100010011;
ROM[26929] <= 32'b00000000001100010010000000100011;
ROM[26930] <= 32'b00000000010000010000000100010011;
ROM[26931] <= 32'b00000000010000010010000000100011;
ROM[26932] <= 32'b00000000010000010000000100010011;
ROM[26933] <= 32'b00000000010100010010000000100011;
ROM[26934] <= 32'b00000000010000010000000100010011;
ROM[26935] <= 32'b00000000011000010010000000100011;
ROM[26936] <= 32'b00000000010000010000000100010011;
ROM[26937] <= 32'b00000001010000000000001110010011;
ROM[26938] <= 32'b00000000100000111000001110010011;
ROM[26939] <= 32'b01000000011100010000001110110011;
ROM[26940] <= 32'b00000000011100000000001000110011;
ROM[26941] <= 32'b00000000001000000000000110110011;
ROM[26942] <= 32'b01101011010000001111000011101111;
ROM[26943] <= 32'b00000111001100000000001110010011;
ROM[26944] <= 32'b00000000011100010010000000100011;
ROM[26945] <= 32'b00000000010000010000000100010011;
ROM[26946] <= 32'b00000000000000011010001110110111;
ROM[26947] <= 32'b01010101010000111000001110010011;
ROM[26948] <= 32'b00000000111000111000001110110011;
ROM[26949] <= 32'b00000000011100010010000000100011;
ROM[26950] <= 32'b00000000010000010000000100010011;
ROM[26951] <= 32'b00000000001100010010000000100011;
ROM[26952] <= 32'b00000000010000010000000100010011;
ROM[26953] <= 32'b00000000010000010010000000100011;
ROM[26954] <= 32'b00000000010000010000000100010011;
ROM[26955] <= 32'b00000000010100010010000000100011;
ROM[26956] <= 32'b00000000010000010000000100010011;
ROM[26957] <= 32'b00000000011000010010000000100011;
ROM[26958] <= 32'b00000000010000010000000100010011;
ROM[26959] <= 32'b00000001010000000000001110010011;
ROM[26960] <= 32'b00000000100000111000001110010011;
ROM[26961] <= 32'b01000000011100010000001110110011;
ROM[26962] <= 32'b00000000011100000000001000110011;
ROM[26963] <= 32'b00000000001000000000000110110011;
ROM[26964] <= 32'b01100101110000001111000011101111;
ROM[26965] <= 32'b00000011101000000000001110010011;
ROM[26966] <= 32'b00000000011100010010000000100011;
ROM[26967] <= 32'b00000000010000010000000100010011;
ROM[26968] <= 32'b00000000000000011010001110110111;
ROM[26969] <= 32'b01011010110000111000001110010011;
ROM[26970] <= 32'b00000000111000111000001110110011;
ROM[26971] <= 32'b00000000011100010010000000100011;
ROM[26972] <= 32'b00000000010000010000000100010011;
ROM[26973] <= 32'b00000000001100010010000000100011;
ROM[26974] <= 32'b00000000010000010000000100010011;
ROM[26975] <= 32'b00000000010000010010000000100011;
ROM[26976] <= 32'b00000000010000010000000100010011;
ROM[26977] <= 32'b00000000010100010010000000100011;
ROM[26978] <= 32'b00000000010000010000000100010011;
ROM[26979] <= 32'b00000000011000010010000000100011;
ROM[26980] <= 32'b00000000010000010000000100010011;
ROM[26981] <= 32'b00000001010000000000001110010011;
ROM[26982] <= 32'b00000000100000111000001110010011;
ROM[26983] <= 32'b01000000011100010000001110110011;
ROM[26984] <= 32'b00000000011100000000001000110011;
ROM[26985] <= 32'b00000000001000000000000110110011;
ROM[26986] <= 32'b01100000010000001111000011101111;
ROM[26987] <= 32'b00000010000000000000001110010011;
ROM[26988] <= 32'b00000000011100010010000000100011;
ROM[26989] <= 32'b00000000010000010000000100010011;
ROM[26990] <= 32'b00000000000000011010001110110111;
ROM[26991] <= 32'b01100000010000111000001110010011;
ROM[26992] <= 32'b00000000111000111000001110110011;
ROM[26993] <= 32'b00000000011100010010000000100011;
ROM[26994] <= 32'b00000000010000010000000100010011;
ROM[26995] <= 32'b00000000001100010010000000100011;
ROM[26996] <= 32'b00000000010000010000000100010011;
ROM[26997] <= 32'b00000000010000010010000000100011;
ROM[26998] <= 32'b00000000010000010000000100010011;
ROM[26999] <= 32'b00000000010100010010000000100011;
ROM[27000] <= 32'b00000000010000010000000100010011;
ROM[27001] <= 32'b00000000011000010010000000100011;
ROM[27002] <= 32'b00000000010000010000000100010011;
ROM[27003] <= 32'b00000001010000000000001110010011;
ROM[27004] <= 32'b00000000100000111000001110010011;
ROM[27005] <= 32'b01000000011100010000001110110011;
ROM[27006] <= 32'b00000000011100000000001000110011;
ROM[27007] <= 32'b00000000001000000000000110110011;
ROM[27008] <= 32'b01011010110000001111000011101111;
ROM[27009] <= 32'b00000000000000011010001110110111;
ROM[27010] <= 32'b01100101000000111000001110010011;
ROM[27011] <= 32'b00000000111000111000001110110011;
ROM[27012] <= 32'b00000000011100010010000000100011;
ROM[27013] <= 32'b00000000010000010000000100010011;
ROM[27014] <= 32'b00000000001100010010000000100011;
ROM[27015] <= 32'b00000000010000010000000100010011;
ROM[27016] <= 32'b00000000010000010010000000100011;
ROM[27017] <= 32'b00000000010000010000000100010011;
ROM[27018] <= 32'b00000000010100010010000000100011;
ROM[27019] <= 32'b00000000010000010000000100010011;
ROM[27020] <= 32'b00000000011000010010000000100011;
ROM[27021] <= 32'b00000000010000010000000100010011;
ROM[27022] <= 32'b00000001010000000000001110010011;
ROM[27023] <= 32'b00000000010000111000001110010011;
ROM[27024] <= 32'b01000000011100010000001110110011;
ROM[27025] <= 32'b00000000011100000000001000110011;
ROM[27026] <= 32'b00000000001000000000000110110011;
ROM[27027] <= 32'b10010001110111111100000011101111;
ROM[27028] <= 32'b11111111110000010000000100010011;
ROM[27029] <= 32'b00000000000000010010001110000011;
ROM[27030] <= 32'b00000000011101100010000000100011;
ROM[27031] <= 32'b00000000000000000000001110010011;
ROM[27032] <= 32'b00000000011100010010000000100011;
ROM[27033] <= 32'b00000000010000010000000100010011;
ROM[27034] <= 32'b11111111110000010000000100010011;
ROM[27035] <= 32'b00000000000000010010001110000011;
ROM[27036] <= 32'b00000000011100011010010000100011;
ROM[27037] <= 32'b00000000100000011010001110000011;
ROM[27038] <= 32'b00000000011100010010000000100011;
ROM[27039] <= 32'b00000000010000010000000100010011;
ROM[27040] <= 32'b00000000010000011010001110000011;
ROM[27041] <= 32'b00000000011100010010000000100011;
ROM[27042] <= 32'b00000000010000010000000100010011;
ROM[27043] <= 32'b11111111110000010000000100010011;
ROM[27044] <= 32'b00000000000000010010001110000011;
ROM[27045] <= 32'b11111111110000010000000100010011;
ROM[27046] <= 32'b00000000000000010010010000000011;
ROM[27047] <= 32'b00000000011101000010001110110011;
ROM[27048] <= 32'b00000000011100010010000000100011;
ROM[27049] <= 32'b00000000010000010000000100010011;
ROM[27050] <= 32'b11111111110000010000000100010011;
ROM[27051] <= 32'b00000000000000010010001110000011;
ROM[27052] <= 32'b01000000011100000000001110110011;
ROM[27053] <= 32'b00000000000100111000001110010011;
ROM[27054] <= 32'b00000000011100010010000000100011;
ROM[27055] <= 32'b00000000010000010000000100010011;
ROM[27056] <= 32'b11111111110000010000000100010011;
ROM[27057] <= 32'b00000000000000010010001110000011;
ROM[27058] <= 32'b00000000000000111000101001100011;
ROM[27059] <= 32'b00000000000000011011001110110111;
ROM[27060] <= 32'b10110011010000111000001110010011;
ROM[27061] <= 32'b00000000111000111000001110110011;
ROM[27062] <= 32'b00000000000000111000000011100111;
ROM[27063] <= 32'b00000000000000011010001110000011;
ROM[27064] <= 32'b00000000011100010010000000100011;
ROM[27065] <= 32'b00000000010000010000000100010011;
ROM[27066] <= 32'b00000000100000011010001110000011;
ROM[27067] <= 32'b00000000011100010010000000100011;
ROM[27068] <= 32'b00000000010000010000000100010011;
ROM[27069] <= 32'b00000000010000000000001110010011;
ROM[27070] <= 32'b00000000011100010010000000100011;
ROM[27071] <= 32'b00000000010000010000000100010011;
ROM[27072] <= 32'b00000000000000011010001110110111;
ROM[27073] <= 32'b01110100110000111000001110010011;
ROM[27074] <= 32'b00000000111000111000001110110011;
ROM[27075] <= 32'b00000000011100010010000000100011;
ROM[27076] <= 32'b00000000010000010000000100010011;
ROM[27077] <= 32'b00000000001100010010000000100011;
ROM[27078] <= 32'b00000000010000010000000100010011;
ROM[27079] <= 32'b00000000010000010010000000100011;
ROM[27080] <= 32'b00000000010000010000000100010011;
ROM[27081] <= 32'b00000000010100010010000000100011;
ROM[27082] <= 32'b00000000010000010000000100010011;
ROM[27083] <= 32'b00000000011000010010000000100011;
ROM[27084] <= 32'b00000000010000010000000100010011;
ROM[27085] <= 32'b00000001010000000000001110010011;
ROM[27086] <= 32'b00000000100000111000001110010011;
ROM[27087] <= 32'b01000000011100010000001110110011;
ROM[27088] <= 32'b00000000011100000000001000110011;
ROM[27089] <= 32'b00000000001000000000000110110011;
ROM[27090] <= 32'b10001110010011110111000011101111;
ROM[27091] <= 32'b11111111110000010000000100010011;
ROM[27092] <= 32'b00000000000000010010001110000011;
ROM[27093] <= 32'b11111111110000010000000100010011;
ROM[27094] <= 32'b00000000000000010010010000000011;
ROM[27095] <= 32'b00000000011101000000001110110011;
ROM[27096] <= 32'b00000000011100010010000000100011;
ROM[27097] <= 32'b00000000010000010000000100010011;
ROM[27098] <= 32'b11111111110000010000000100010011;
ROM[27099] <= 32'b00000000000000010010001110000011;
ROM[27100] <= 32'b00000000000000111000001100010011;
ROM[27101] <= 32'b00000000110100110000010000110011;
ROM[27102] <= 32'b00000000000001000010001110000011;
ROM[27103] <= 32'b00000000011100010010000000100011;
ROM[27104] <= 32'b00000000010000010000000100010011;
ROM[27105] <= 32'b00000000000000011010001110110111;
ROM[27106] <= 32'b01111101000000111000001110010011;
ROM[27107] <= 32'b00000000111000111000001110110011;
ROM[27108] <= 32'b00000000011100010010000000100011;
ROM[27109] <= 32'b00000000010000010000000100010011;
ROM[27110] <= 32'b00000000001100010010000000100011;
ROM[27111] <= 32'b00000000010000010000000100010011;
ROM[27112] <= 32'b00000000010000010010000000100011;
ROM[27113] <= 32'b00000000010000010000000100010011;
ROM[27114] <= 32'b00000000010100010010000000100011;
ROM[27115] <= 32'b00000000010000010000000100010011;
ROM[27116] <= 32'b00000000011000010010000000100011;
ROM[27117] <= 32'b00000000010000010000000100010011;
ROM[27118] <= 32'b00000001010000000000001110010011;
ROM[27119] <= 32'b00000000010000111000001110010011;
ROM[27120] <= 32'b01000000011100010000001110110011;
ROM[27121] <= 32'b00000000011100000000001000110011;
ROM[27122] <= 32'b00000000001000000000000110110011;
ROM[27123] <= 32'b10011011010111111100000011101111;
ROM[27124] <= 32'b11111111110000010000000100010011;
ROM[27125] <= 32'b00000000000000010010001110000011;
ROM[27126] <= 32'b00000000011101100010000000100011;
ROM[27127] <= 32'b00000000100000011010001110000011;
ROM[27128] <= 32'b00000000011100010010000000100011;
ROM[27129] <= 32'b00000000010000010000000100010011;
ROM[27130] <= 32'b00000000000100000000001110010011;
ROM[27131] <= 32'b00000000011100010010000000100011;
ROM[27132] <= 32'b00000000010000010000000100010011;
ROM[27133] <= 32'b11111111110000010000000100010011;
ROM[27134] <= 32'b00000000000000010010001110000011;
ROM[27135] <= 32'b11111111110000010000000100010011;
ROM[27136] <= 32'b00000000000000010010010000000011;
ROM[27137] <= 32'b00000000011101000000001110110011;
ROM[27138] <= 32'b00000000011100010010000000100011;
ROM[27139] <= 32'b00000000010000010000000100010011;
ROM[27140] <= 32'b11111111110000010000000100010011;
ROM[27141] <= 32'b00000000000000010010001110000011;
ROM[27142] <= 32'b00000000011100011010010000100011;
ROM[27143] <= 32'b00000000100000011010001110000011;
ROM[27144] <= 32'b00000000011100010010000000100011;
ROM[27145] <= 32'b00000000010000010000000100010011;
ROM[27146] <= 32'b00000000010000011010001110000011;
ROM[27147] <= 32'b00000000011100010010000000100011;
ROM[27148] <= 32'b00000000010000010000000100010011;
ROM[27149] <= 32'b11111111110000010000000100010011;
ROM[27150] <= 32'b00000000000000010010001110000011;
ROM[27151] <= 32'b11111111110000010000000100010011;
ROM[27152] <= 32'b00000000000000010010010000000011;
ROM[27153] <= 32'b00000000011101000010001110110011;
ROM[27154] <= 32'b00000000011100010010000000100011;
ROM[27155] <= 32'b00000000010000010000000100010011;
ROM[27156] <= 32'b11111111110000010000000100010011;
ROM[27157] <= 32'b00000000000000010010001110000011;
ROM[27158] <= 32'b00000000000000111000101001100011;
ROM[27159] <= 32'b00000000000000011011001110110111;
ROM[27160] <= 32'b10011101000000111000001110010011;
ROM[27161] <= 32'b00000000111000111000001110110011;
ROM[27162] <= 32'b00000000000000111000000011100111;
ROM[27163] <= 32'b00000000001000000000001110010011;
ROM[27164] <= 32'b00000000011100010010000000100011;
ROM[27165] <= 32'b00000000010000010000000100010011;
ROM[27166] <= 32'b00000000000000011011001110110111;
ROM[27167] <= 32'b10001100010000111000001110010011;
ROM[27168] <= 32'b00000000111000111000001110110011;
ROM[27169] <= 32'b00000000011100010010000000100011;
ROM[27170] <= 32'b00000000010000010000000100010011;
ROM[27171] <= 32'b00000000001100010010000000100011;
ROM[27172] <= 32'b00000000010000010000000100010011;
ROM[27173] <= 32'b00000000010000010010000000100011;
ROM[27174] <= 32'b00000000010000010000000100010011;
ROM[27175] <= 32'b00000000010100010010000000100011;
ROM[27176] <= 32'b00000000010000010000000100010011;
ROM[27177] <= 32'b00000000011000010010000000100011;
ROM[27178] <= 32'b00000000010000010000000100010011;
ROM[27179] <= 32'b00000001010000000000001110010011;
ROM[27180] <= 32'b00000000010000111000001110010011;
ROM[27181] <= 32'b01000000011100010000001110110011;
ROM[27182] <= 32'b00000000011100000000001000110011;
ROM[27183] <= 32'b00000000001000000000000110110011;
ROM[27184] <= 32'b01100111110100001110000011101111;
ROM[27185] <= 32'b00000101110000000000001110010011;
ROM[27186] <= 32'b00000000011100010010000000100011;
ROM[27187] <= 32'b00000000010000010000000100010011;
ROM[27188] <= 32'b00000000000000011011001110110111;
ROM[27189] <= 32'b10010001110000111000001110010011;
ROM[27190] <= 32'b00000000111000111000001110110011;
ROM[27191] <= 32'b00000000011100010010000000100011;
ROM[27192] <= 32'b00000000010000010000000100010011;
ROM[27193] <= 32'b00000000001100010010000000100011;
ROM[27194] <= 32'b00000000010000010000000100010011;
ROM[27195] <= 32'b00000000010000010010000000100011;
ROM[27196] <= 32'b00000000010000010000000100010011;
ROM[27197] <= 32'b00000000010100010010000000100011;
ROM[27198] <= 32'b00000000010000010000000100010011;
ROM[27199] <= 32'b00000000011000010010000000100011;
ROM[27200] <= 32'b00000000010000010000000100010011;
ROM[27201] <= 32'b00000001010000000000001110010011;
ROM[27202] <= 32'b00000000100000111000001110010011;
ROM[27203] <= 32'b01000000011100010000001110110011;
ROM[27204] <= 32'b00000000011100000000001000110011;
ROM[27205] <= 32'b00000000001000000000000110110011;
ROM[27206] <= 32'b00101001010000001111000011101111;
ROM[27207] <= 32'b00000110111000000000001110010011;
ROM[27208] <= 32'b00000000011100010010000000100011;
ROM[27209] <= 32'b00000000010000010000000100010011;
ROM[27210] <= 32'b00000000000000011011001110110111;
ROM[27211] <= 32'b10010111010000111000001110010011;
ROM[27212] <= 32'b00000000111000111000001110110011;
ROM[27213] <= 32'b00000000011100010010000000100011;
ROM[27214] <= 32'b00000000010000010000000100010011;
ROM[27215] <= 32'b00000000001100010010000000100011;
ROM[27216] <= 32'b00000000010000010000000100010011;
ROM[27217] <= 32'b00000000010000010010000000100011;
ROM[27218] <= 32'b00000000010000010000000100010011;
ROM[27219] <= 32'b00000000010100010010000000100011;
ROM[27220] <= 32'b00000000010000010000000100010011;
ROM[27221] <= 32'b00000000011000010010000000100011;
ROM[27222] <= 32'b00000000010000010000000100010011;
ROM[27223] <= 32'b00000001010000000000001110010011;
ROM[27224] <= 32'b00000000100000111000001110010011;
ROM[27225] <= 32'b01000000011100010000001110110011;
ROM[27226] <= 32'b00000000011100000000001000110011;
ROM[27227] <= 32'b00000000001000000000000110110011;
ROM[27228] <= 32'b00100011110000001111000011101111;
ROM[27229] <= 32'b00000000000000011011001110110111;
ROM[27230] <= 32'b10011100000000111000001110010011;
ROM[27231] <= 32'b00000000111000111000001110110011;
ROM[27232] <= 32'b00000000011100010010000000100011;
ROM[27233] <= 32'b00000000010000010000000100010011;
ROM[27234] <= 32'b00000000001100010010000000100011;
ROM[27235] <= 32'b00000000010000010000000100010011;
ROM[27236] <= 32'b00000000010000010010000000100011;
ROM[27237] <= 32'b00000000010000010000000100010011;
ROM[27238] <= 32'b00000000010100010010000000100011;
ROM[27239] <= 32'b00000000010000010000000100010011;
ROM[27240] <= 32'b00000000011000010010000000100011;
ROM[27241] <= 32'b00000000010000010000000100010011;
ROM[27242] <= 32'b00000001010000000000001110010011;
ROM[27243] <= 32'b00000000010000111000001110010011;
ROM[27244] <= 32'b01000000011100010000001110110011;
ROM[27245] <= 32'b00000000011100000000001000110011;
ROM[27246] <= 32'b00000000001000000000000110110011;
ROM[27247] <= 32'b11011010110011111100000011101111;
ROM[27248] <= 32'b11111111110000010000000100010011;
ROM[27249] <= 32'b00000000000000010010001110000011;
ROM[27250] <= 32'b00000000011101100010000000100011;
ROM[27251] <= 32'b00010110010000000000000011101111;
ROM[27252] <= 32'b00000000001000000000001110010011;
ROM[27253] <= 32'b00000000011100010010000000100011;
ROM[27254] <= 32'b00000000010000010000000100010011;
ROM[27255] <= 32'b00000000000000011011001110110111;
ROM[27256] <= 32'b10100010100000111000001110010011;
ROM[27257] <= 32'b00000000111000111000001110110011;
ROM[27258] <= 32'b00000000011100010010000000100011;
ROM[27259] <= 32'b00000000010000010000000100010011;
ROM[27260] <= 32'b00000000001100010010000000100011;
ROM[27261] <= 32'b00000000010000010000000100010011;
ROM[27262] <= 32'b00000000010000010010000000100011;
ROM[27263] <= 32'b00000000010000010000000100010011;
ROM[27264] <= 32'b00000000010100010010000000100011;
ROM[27265] <= 32'b00000000010000010000000100010011;
ROM[27266] <= 32'b00000000011000010010000000100011;
ROM[27267] <= 32'b00000000010000010000000100010011;
ROM[27268] <= 32'b00000001010000000000001110010011;
ROM[27269] <= 32'b00000000010000111000001110010011;
ROM[27270] <= 32'b01000000011100010000001110110011;
ROM[27271] <= 32'b00000000011100000000001000110011;
ROM[27272] <= 32'b00000000001000000000000110110011;
ROM[27273] <= 32'b01010001100100001110000011101111;
ROM[27274] <= 32'b00000010110000000000001110010011;
ROM[27275] <= 32'b00000000011100010010000000100011;
ROM[27276] <= 32'b00000000010000010000000100010011;
ROM[27277] <= 32'b00000000000000011011001110110111;
ROM[27278] <= 32'b10101000000000111000001110010011;
ROM[27279] <= 32'b00000000111000111000001110110011;
ROM[27280] <= 32'b00000000011100010010000000100011;
ROM[27281] <= 32'b00000000010000010000000100010011;
ROM[27282] <= 32'b00000000001100010010000000100011;
ROM[27283] <= 32'b00000000010000010000000100010011;
ROM[27284] <= 32'b00000000010000010010000000100011;
ROM[27285] <= 32'b00000000010000010000000100010011;
ROM[27286] <= 32'b00000000010100010010000000100011;
ROM[27287] <= 32'b00000000010000010000000100010011;
ROM[27288] <= 32'b00000000011000010010000000100011;
ROM[27289] <= 32'b00000000010000010000000100010011;
ROM[27290] <= 32'b00000001010000000000001110010011;
ROM[27291] <= 32'b00000000100000111000001110010011;
ROM[27292] <= 32'b01000000011100010000001110110011;
ROM[27293] <= 32'b00000000011100000000001000110011;
ROM[27294] <= 32'b00000000001000000000000110110011;
ROM[27295] <= 32'b00010011000000001111000011101111;
ROM[27296] <= 32'b00000010000000000000001110010011;
ROM[27297] <= 32'b00000000011100010010000000100011;
ROM[27298] <= 32'b00000000010000010000000100010011;
ROM[27299] <= 32'b00000000000000011011001110110111;
ROM[27300] <= 32'b10101101100000111000001110010011;
ROM[27301] <= 32'b00000000111000111000001110110011;
ROM[27302] <= 32'b00000000011100010010000000100011;
ROM[27303] <= 32'b00000000010000010000000100010011;
ROM[27304] <= 32'b00000000001100010010000000100011;
ROM[27305] <= 32'b00000000010000010000000100010011;
ROM[27306] <= 32'b00000000010000010010000000100011;
ROM[27307] <= 32'b00000000010000010000000100010011;
ROM[27308] <= 32'b00000000010100010010000000100011;
ROM[27309] <= 32'b00000000010000010000000100010011;
ROM[27310] <= 32'b00000000011000010010000000100011;
ROM[27311] <= 32'b00000000010000010000000100010011;
ROM[27312] <= 32'b00000001010000000000001110010011;
ROM[27313] <= 32'b00000000100000111000001110010011;
ROM[27314] <= 32'b01000000011100010000001110110011;
ROM[27315] <= 32'b00000000011100000000001000110011;
ROM[27316] <= 32'b00000000001000000000000110110011;
ROM[27317] <= 32'b00001101100000001111000011101111;
ROM[27318] <= 32'b00000000000000011011001110110111;
ROM[27319] <= 32'b10110010010000111000001110010011;
ROM[27320] <= 32'b00000000111000111000001110110011;
ROM[27321] <= 32'b00000000011100010010000000100011;
ROM[27322] <= 32'b00000000010000010000000100010011;
ROM[27323] <= 32'b00000000001100010010000000100011;
ROM[27324] <= 32'b00000000010000010000000100010011;
ROM[27325] <= 32'b00000000010000010010000000100011;
ROM[27326] <= 32'b00000000010000010000000100010011;
ROM[27327] <= 32'b00000000010100010010000000100011;
ROM[27328] <= 32'b00000000010000010000000100010011;
ROM[27329] <= 32'b00000000011000010010000000100011;
ROM[27330] <= 32'b00000000010000010000000100010011;
ROM[27331] <= 32'b00000001010000000000001110010011;
ROM[27332] <= 32'b00000000010000111000001110010011;
ROM[27333] <= 32'b01000000011100010000001110110011;
ROM[27334] <= 32'b00000000011100000000001000110011;
ROM[27335] <= 32'b00000000001000000000000110110011;
ROM[27336] <= 32'b11000100100011111100000011101111;
ROM[27337] <= 32'b11111111110000010000000100010011;
ROM[27338] <= 32'b00000000000000010010001110000011;
ROM[27339] <= 32'b00000000011101100010000000100011;
ROM[27340] <= 32'b10110100010111111111000011101111;
ROM[27341] <= 32'b00000000000000000000001110010011;
ROM[27342] <= 32'b00000000011100010010000000100011;
ROM[27343] <= 32'b00000000010000010000000100010011;
ROM[27344] <= 32'b00000001010000000000001110010011;
ROM[27345] <= 32'b01000000011100011000001110110011;
ROM[27346] <= 32'b00000000000000111010000010000011;
ROM[27347] <= 32'b11111111110000010000000100010011;
ROM[27348] <= 32'b00000000000000010010001110000011;
ROM[27349] <= 32'b00000000011100100010000000100011;
ROM[27350] <= 32'b00000000010000100000000100010011;
ROM[27351] <= 32'b00000001010000000000001110010011;
ROM[27352] <= 32'b01000000011100011000001110110011;
ROM[27353] <= 32'b00000000010000111010000110000011;
ROM[27354] <= 32'b00000000100000111010001000000011;
ROM[27355] <= 32'b00000000110000111010001010000011;
ROM[27356] <= 32'b00000001000000111010001100000011;
ROM[27357] <= 32'b00000000000000001000000011100111;
ROM[27358] <= 32'b00000000000000010010000000100011;
ROM[27359] <= 32'b00000000010000010000000100010011;
ROM[27360] <= 32'b00000000010000100010001110000011;
ROM[27361] <= 32'b00000000011100010010000000100011;
ROM[27362] <= 32'b00000000010000010000000100010011;
ROM[27363] <= 32'b00000000100000100010001110000011;
ROM[27364] <= 32'b00000000011100010010000000100011;
ROM[27365] <= 32'b00000000010000010000000100010011;
ROM[27366] <= 32'b11111111110000010000000100010011;
ROM[27367] <= 32'b00000000000000010010001110000011;
ROM[27368] <= 32'b11111111110000010000000100010011;
ROM[27369] <= 32'b00000000000000010010010000000011;
ROM[27370] <= 32'b00000000011101000010001110110011;
ROM[27371] <= 32'b00000000011100010010000000100011;
ROM[27372] <= 32'b00000000010000010000000100010011;
ROM[27373] <= 32'b11111111110000010000000100010011;
ROM[27374] <= 32'b00000000000000010010001110000011;
ROM[27375] <= 32'b00000000000000111000101001100011;
ROM[27376] <= 32'b00000000000000011011001110110111;
ROM[27377] <= 32'b10111101010000111000001110010011;
ROM[27378] <= 32'b00000000111000111000001110110011;
ROM[27379] <= 32'b00000000000000111000000011100111;
ROM[27380] <= 32'b00011100100000000000000011101111;
ROM[27381] <= 32'b00000000000000100010001110000011;
ROM[27382] <= 32'b00000000011100010010000000100011;
ROM[27383] <= 32'b00000000010000010000000100010011;
ROM[27384] <= 32'b00000000010000100010001110000011;
ROM[27385] <= 32'b00000000011100010010000000100011;
ROM[27386] <= 32'b00000000010000010000000100010011;
ROM[27387] <= 32'b00000000100000100010001110000011;
ROM[27388] <= 32'b00000000011100010010000000100011;
ROM[27389] <= 32'b00000000010000010000000100010011;
ROM[27390] <= 32'b00000000000000011011001110110111;
ROM[27391] <= 32'b11000100010000111000001110010011;
ROM[27392] <= 32'b00000000111000111000001110110011;
ROM[27393] <= 32'b00000000011100010010000000100011;
ROM[27394] <= 32'b00000000010000010000000100010011;
ROM[27395] <= 32'b00000000001100010010000000100011;
ROM[27396] <= 32'b00000000010000010000000100010011;
ROM[27397] <= 32'b00000000010000010010000000100011;
ROM[27398] <= 32'b00000000010000010000000100010011;
ROM[27399] <= 32'b00000000010100010010000000100011;
ROM[27400] <= 32'b00000000010000010000000100010011;
ROM[27401] <= 32'b00000000011000010010000000100011;
ROM[27402] <= 32'b00000000010000010000000100010011;
ROM[27403] <= 32'b00000001010000000000001110010011;
ROM[27404] <= 32'b00000000110000111000001110010011;
ROM[27405] <= 32'b01000000011100010000001110110011;
ROM[27406] <= 32'b00000000011100000000001000110011;
ROM[27407] <= 32'b00000000001000000000000110110011;
ROM[27408] <= 32'b00011001110000000000000011101111;
ROM[27409] <= 32'b11111111110000010000000100010011;
ROM[27410] <= 32'b00000000000000010010001110000011;
ROM[27411] <= 32'b00000000011100011010000000100011;
ROM[27412] <= 32'b00000000000000100010001110000011;
ROM[27413] <= 32'b00000000011100010010000000100011;
ROM[27414] <= 32'b00000000010000010000000100010011;
ROM[27415] <= 32'b00000000010000100010001110000011;
ROM[27416] <= 32'b00000000011100010010000000100011;
ROM[27417] <= 32'b00000000010000010000000100010011;
ROM[27418] <= 32'b00000000000000011010001110000011;
ROM[27419] <= 32'b00000000011100010010000000100011;
ROM[27420] <= 32'b00000000010000010000000100010011;
ROM[27421] <= 32'b00000000000100000000001110010011;
ROM[27422] <= 32'b00000000011100010010000000100011;
ROM[27423] <= 32'b00000000010000010000000100010011;
ROM[27424] <= 32'b11111111110000010000000100010011;
ROM[27425] <= 32'b00000000000000010010001110000011;
ROM[27426] <= 32'b11111111110000010000000100010011;
ROM[27427] <= 32'b00000000000000010010010000000011;
ROM[27428] <= 32'b01000000011101000000001110110011;
ROM[27429] <= 32'b00000000011100010010000000100011;
ROM[27430] <= 32'b00000000010000010000000100010011;
ROM[27431] <= 32'b00000000000000011011001110110111;
ROM[27432] <= 32'b11001110100000111000001110010011;
ROM[27433] <= 32'b00000000111000111000001110110011;
ROM[27434] <= 32'b00000000011100010010000000100011;
ROM[27435] <= 32'b00000000010000010000000100010011;
ROM[27436] <= 32'b00000000001100010010000000100011;
ROM[27437] <= 32'b00000000010000010000000100010011;
ROM[27438] <= 32'b00000000010000010010000000100011;
ROM[27439] <= 32'b00000000010000010000000100010011;
ROM[27440] <= 32'b00000000010100010010000000100011;
ROM[27441] <= 32'b00000000010000010000000100010011;
ROM[27442] <= 32'b00000000011000010010000000100011;
ROM[27443] <= 32'b00000000010000010000000100010011;
ROM[27444] <= 32'b00000001010000000000001110010011;
ROM[27445] <= 32'b00000000110000111000001110010011;
ROM[27446] <= 32'b01000000011100010000001110110011;
ROM[27447] <= 32'b00000000011100000000001000110011;
ROM[27448] <= 32'b00000000001000000000000110110011;
ROM[27449] <= 32'b11101001010111111111000011101111;
ROM[27450] <= 32'b11111111110000010000000100010011;
ROM[27451] <= 32'b00000000000000010010001110000011;
ROM[27452] <= 32'b00000000011101100010000000100011;
ROM[27453] <= 32'b00000000000000100010001110000011;
ROM[27454] <= 32'b00000000011100010010000000100011;
ROM[27455] <= 32'b00000000010000010000000100010011;
ROM[27456] <= 32'b00000000000000011010001110000011;
ROM[27457] <= 32'b00000000011100010010000000100011;
ROM[27458] <= 32'b00000000010000010000000100010011;
ROM[27459] <= 32'b00000000000100000000001110010011;
ROM[27460] <= 32'b00000000011100010010000000100011;
ROM[27461] <= 32'b00000000010000010000000100010011;
ROM[27462] <= 32'b11111111110000010000000100010011;
ROM[27463] <= 32'b00000000000000010010001110000011;
ROM[27464] <= 32'b11111111110000010000000100010011;
ROM[27465] <= 32'b00000000000000010010010000000011;
ROM[27466] <= 32'b00000000011101000000001110110011;
ROM[27467] <= 32'b00000000011100010010000000100011;
ROM[27468] <= 32'b00000000010000010000000100010011;
ROM[27469] <= 32'b00000000100000100010001110000011;
ROM[27470] <= 32'b00000000011100010010000000100011;
ROM[27471] <= 32'b00000000010000010000000100010011;
ROM[27472] <= 32'b00000000000000011011001110110111;
ROM[27473] <= 32'b11011000110000111000001110010011;
ROM[27474] <= 32'b00000000111000111000001110110011;
ROM[27475] <= 32'b00000000011100010010000000100011;
ROM[27476] <= 32'b00000000010000010000000100010011;
ROM[27477] <= 32'b00000000001100010010000000100011;
ROM[27478] <= 32'b00000000010000010000000100010011;
ROM[27479] <= 32'b00000000010000010010000000100011;
ROM[27480] <= 32'b00000000010000010000000100010011;
ROM[27481] <= 32'b00000000010100010010000000100011;
ROM[27482] <= 32'b00000000010000010000000100010011;
ROM[27483] <= 32'b00000000011000010010000000100011;
ROM[27484] <= 32'b00000000010000010000000100010011;
ROM[27485] <= 32'b00000001010000000000001110010011;
ROM[27486] <= 32'b00000000110000111000001110010011;
ROM[27487] <= 32'b01000000011100010000001110110011;
ROM[27488] <= 32'b00000000011100000000001000110011;
ROM[27489] <= 32'b00000000001000000000000110110011;
ROM[27490] <= 32'b11011111000111111111000011101111;
ROM[27491] <= 32'b11111111110000010000000100010011;
ROM[27492] <= 32'b00000000000000010010001110000011;
ROM[27493] <= 32'b00000000011101100010000000100011;
ROM[27494] <= 32'b00000000000000000000001110010011;
ROM[27495] <= 32'b00000000011100010010000000100011;
ROM[27496] <= 32'b00000000010000010000000100010011;
ROM[27497] <= 32'b00000001010000000000001110010011;
ROM[27498] <= 32'b01000000011100011000001110110011;
ROM[27499] <= 32'b00000000000000111010000010000011;
ROM[27500] <= 32'b11111111110000010000000100010011;
ROM[27501] <= 32'b00000000000000010010001110000011;
ROM[27502] <= 32'b00000000011100100010000000100011;
ROM[27503] <= 32'b00000000010000100000000100010011;
ROM[27504] <= 32'b00000001010000000000001110010011;
ROM[27505] <= 32'b01000000011100011000001110110011;
ROM[27506] <= 32'b00000000010000111010000110000011;
ROM[27507] <= 32'b00000000100000111010001000000011;
ROM[27508] <= 32'b00000000110000111010001010000011;
ROM[27509] <= 32'b00000001000000111010001100000011;
ROM[27510] <= 32'b00000000000000001000000011100111;
ROM[27511] <= 32'b00000000000000010010000000100011;
ROM[27512] <= 32'b00000000010000010000000100010011;
ROM[27513] <= 32'b00000000000000010010000000100011;
ROM[27514] <= 32'b00000000010000010000000100010011;
ROM[27515] <= 32'b00000000000000010010000000100011;
ROM[27516] <= 32'b00000000010000010000000100010011;
ROM[27517] <= 32'b00000000000000010010000000100011;
ROM[27518] <= 32'b00000000010000010000000100010011;
ROM[27519] <= 32'b00000000000000100010001110000011;
ROM[27520] <= 32'b00000000011100010010000000100011;
ROM[27521] <= 32'b00000000010000010000000100010011;
ROM[27522] <= 32'b00000000100000100010001110000011;
ROM[27523] <= 32'b00000000011100010010000000100011;
ROM[27524] <= 32'b00000000010000010000000100010011;
ROM[27525] <= 32'b00000000010000000000001110010011;
ROM[27526] <= 32'b00000000011100010010000000100011;
ROM[27527] <= 32'b00000000010000010000000100010011;
ROM[27528] <= 32'b00000000000000011011001110110111;
ROM[27529] <= 32'b11100110110000111000001110010011;
ROM[27530] <= 32'b00000000111000111000001110110011;
ROM[27531] <= 32'b00000000011100010010000000100011;
ROM[27532] <= 32'b00000000010000010000000100010011;
ROM[27533] <= 32'b00000000001100010010000000100011;
ROM[27534] <= 32'b00000000010000010000000100010011;
ROM[27535] <= 32'b00000000010000010010000000100011;
ROM[27536] <= 32'b00000000010000010000000100010011;
ROM[27537] <= 32'b00000000010100010010000000100011;
ROM[27538] <= 32'b00000000010000010000000100010011;
ROM[27539] <= 32'b00000000011000010010000000100011;
ROM[27540] <= 32'b00000000010000010000000100010011;
ROM[27541] <= 32'b00000001010000000000001110010011;
ROM[27542] <= 32'b00000000100000111000001110010011;
ROM[27543] <= 32'b01000000011100010000001110110011;
ROM[27544] <= 32'b00000000011100000000001000110011;
ROM[27545] <= 32'b00000000001000000000000110110011;
ROM[27546] <= 32'b10011100010111110110000011101111;
ROM[27547] <= 32'b11111111110000010000000100010011;
ROM[27548] <= 32'b00000000000000010010001110000011;
ROM[27549] <= 32'b11111111110000010000000100010011;
ROM[27550] <= 32'b00000000000000010010010000000011;
ROM[27551] <= 32'b00000000011101000000001110110011;
ROM[27552] <= 32'b00000000011100010010000000100011;
ROM[27553] <= 32'b00000000010000010000000100010011;
ROM[27554] <= 32'b11111111110000010000000100010011;
ROM[27555] <= 32'b00000000000000010010001110000011;
ROM[27556] <= 32'b00000000000000111000001100010011;
ROM[27557] <= 32'b00000000110100110000010000110011;
ROM[27558] <= 32'b00000000000001000010001110000011;
ROM[27559] <= 32'b00000000011100010010000000100011;
ROM[27560] <= 32'b00000000010000010000000100010011;
ROM[27561] <= 32'b11111111110000010000000100010011;
ROM[27562] <= 32'b00000000000000010010001110000011;
ROM[27563] <= 32'b00000000011100011010000000100011;
ROM[27564] <= 32'b00000000010000100010001110000011;
ROM[27565] <= 32'b00000000011100010010000000100011;
ROM[27566] <= 32'b00000000010000010000000100010011;
ROM[27567] <= 32'b00000000000100000000001110010011;
ROM[27568] <= 32'b00000000011100010010000000100011;
ROM[27569] <= 32'b00000000010000010000000100010011;
ROM[27570] <= 32'b11111111110000010000000100010011;
ROM[27571] <= 32'b00000000000000010010001110000011;
ROM[27572] <= 32'b11111111110000010000000100010011;
ROM[27573] <= 32'b00000000000000010010010000000011;
ROM[27574] <= 32'b01000000011101000000001110110011;
ROM[27575] <= 32'b00000000011100010010000000100011;
ROM[27576] <= 32'b00000000010000010000000100010011;
ROM[27577] <= 32'b11111111110000010000000100010011;
ROM[27578] <= 32'b00000000000000010010001110000011;
ROM[27579] <= 32'b00000000011100011010001000100011;
ROM[27580] <= 32'b00000000010000100010001110000011;
ROM[27581] <= 32'b00000000011100010010000000100011;
ROM[27582] <= 32'b00000000010000010000000100010011;
ROM[27583] <= 32'b11111111110000010000000100010011;
ROM[27584] <= 32'b00000000000000010010001110000011;
ROM[27585] <= 32'b00000000011100011010010000100011;
ROM[27586] <= 32'b00000000100000011010001110000011;
ROM[27587] <= 32'b00000000011100010010000000100011;
ROM[27588] <= 32'b00000000010000010000000100010011;
ROM[27589] <= 32'b00000000100000100010001110000011;
ROM[27590] <= 32'b00000000011100010010000000100011;
ROM[27591] <= 32'b00000000010000010000000100010011;
ROM[27592] <= 32'b11111111110000010000000100010011;
ROM[27593] <= 32'b00000000000000010010001110000011;
ROM[27594] <= 32'b11111111110000010000000100010011;
ROM[27595] <= 32'b00000000000000010010010000000011;
ROM[27596] <= 32'b00000000011101000010001110110011;
ROM[27597] <= 32'b00000000011100010010000000100011;
ROM[27598] <= 32'b00000000010000010000000100010011;
ROM[27599] <= 32'b11111111110000010000000100010011;
ROM[27600] <= 32'b00000000000000010010001110000011;
ROM[27601] <= 32'b01000000011100000000001110110011;
ROM[27602] <= 32'b00000000000100111000001110010011;
ROM[27603] <= 32'b00000000011100010010000000100011;
ROM[27604] <= 32'b00000000010000010000000100010011;
ROM[27605] <= 32'b11111111110000010000000100010011;
ROM[27606] <= 32'b00000000000000010010001110000011;
ROM[27607] <= 32'b00000000000000111000101001100011;
ROM[27608] <= 32'b00000000000000011011001110110111;
ROM[27609] <= 32'b00111001110000111000001110010011;
ROM[27610] <= 32'b00000000111000111000001110110011;
ROM[27611] <= 32'b00000000000000111000000011100111;
ROM[27612] <= 32'b00000000000000100010001110000011;
ROM[27613] <= 32'b00000000011100010010000000100011;
ROM[27614] <= 32'b00000000010000010000000100010011;
ROM[27615] <= 32'b00000000100000011010001110000011;
ROM[27616] <= 32'b00000000011100010010000000100011;
ROM[27617] <= 32'b00000000010000010000000100010011;
ROM[27618] <= 32'b00000000010000000000001110010011;
ROM[27619] <= 32'b00000000011100010010000000100011;
ROM[27620] <= 32'b00000000010000010000000100010011;
ROM[27621] <= 32'b00000000000000011011001110110111;
ROM[27622] <= 32'b11111110000000111000001110010011;
ROM[27623] <= 32'b00000000111000111000001110110011;
ROM[27624] <= 32'b00000000011100010010000000100011;
ROM[27625] <= 32'b00000000010000010000000100010011;
ROM[27626] <= 32'b00000000001100010010000000100011;
ROM[27627] <= 32'b00000000010000010000000100010011;
ROM[27628] <= 32'b00000000010000010010000000100011;
ROM[27629] <= 32'b00000000010000010000000100010011;
ROM[27630] <= 32'b00000000010100010010000000100011;
ROM[27631] <= 32'b00000000010000010000000100010011;
ROM[27632] <= 32'b00000000011000010010000000100011;
ROM[27633] <= 32'b00000000010000010000000100010011;
ROM[27634] <= 32'b00000001010000000000001110010011;
ROM[27635] <= 32'b00000000100000111000001110010011;
ROM[27636] <= 32'b01000000011100010000001110110011;
ROM[27637] <= 32'b00000000011100000000001000110011;
ROM[27638] <= 32'b00000000001000000000000110110011;
ROM[27639] <= 32'b10000101000111110110000011101111;
ROM[27640] <= 32'b11111111110000010000000100010011;
ROM[27641] <= 32'b00000000000000010010001110000011;
ROM[27642] <= 32'b11111111110000010000000100010011;
ROM[27643] <= 32'b00000000000000010010010000000011;
ROM[27644] <= 32'b00000000011101000000001110110011;
ROM[27645] <= 32'b00000000011100010010000000100011;
ROM[27646] <= 32'b00000000010000010000000100010011;
ROM[27647] <= 32'b11111111110000010000000100010011;
ROM[27648] <= 32'b00000000000000010010001110000011;
ROM[27649] <= 32'b00000000000000111000001100010011;
ROM[27650] <= 32'b00000000110100110000010000110011;
ROM[27651] <= 32'b00000000000001000010001110000011;
ROM[27652] <= 32'b00000000011100010010000000100011;
ROM[27653] <= 32'b00000000010000010000000100010011;
ROM[27654] <= 32'b00000000000000011010001110000011;
ROM[27655] <= 32'b00000000011100010010000000100011;
ROM[27656] <= 32'b00000000010000010000000100010011;
ROM[27657] <= 32'b11111111110000010000000100010011;
ROM[27658] <= 32'b00000000000000010010001110000011;
ROM[27659] <= 32'b11111111110000010000000100010011;
ROM[27660] <= 32'b00000000000000010010010000000011;
ROM[27661] <= 32'b00000000011101000010001110110011;
ROM[27662] <= 32'b00000000011100010010000000100011;
ROM[27663] <= 32'b00000000010000010000000100010011;
ROM[27664] <= 32'b11111111110000010000000100010011;
ROM[27665] <= 32'b00000000000000010010001110000011;
ROM[27666] <= 32'b00000000000000111000101001100011;
ROM[27667] <= 32'b00000000000000011011001110110111;
ROM[27668] <= 32'b00000110000000111000001110010011;
ROM[27669] <= 32'b00000000111000111000001110110011;
ROM[27670] <= 32'b00000000000000111000000011100111;
ROM[27671] <= 32'b00101111110000000000000011101111;
ROM[27672] <= 32'b00000000010000011010001110000011;
ROM[27673] <= 32'b00000000011100010010000000100011;
ROM[27674] <= 32'b00000000010000010000000100010011;
ROM[27675] <= 32'b00000000000100000000001110010011;
ROM[27676] <= 32'b00000000011100010010000000100011;
ROM[27677] <= 32'b00000000010000010000000100010011;
ROM[27678] <= 32'b11111111110000010000000100010011;
ROM[27679] <= 32'b00000000000000010010001110000011;
ROM[27680] <= 32'b11111111110000010000000100010011;
ROM[27681] <= 32'b00000000000000010010010000000011;
ROM[27682] <= 32'b00000000011101000000001110110011;
ROM[27683] <= 32'b00000000011100010010000000100011;
ROM[27684] <= 32'b00000000010000010000000100010011;
ROM[27685] <= 32'b11111111110000010000000100010011;
ROM[27686] <= 32'b00000000000000010010001110000011;
ROM[27687] <= 32'b00000000011100011010001000100011;
ROM[27688] <= 32'b00000000000000100010001110000011;
ROM[27689] <= 32'b00000000011100010010000000100011;
ROM[27690] <= 32'b00000000010000010000000100010011;
ROM[27691] <= 32'b00000000010000011010001110000011;
ROM[27692] <= 32'b00000000011100010010000000100011;
ROM[27693] <= 32'b00000000010000010000000100010011;
ROM[27694] <= 32'b00000000010000000000001110010011;
ROM[27695] <= 32'b00000000011100010010000000100011;
ROM[27696] <= 32'b00000000010000010000000100010011;
ROM[27697] <= 32'b00000000000000011011001110110111;
ROM[27698] <= 32'b00010001000000111000001110010011;
ROM[27699] <= 32'b00000000111000111000001110110011;
ROM[27700] <= 32'b00000000011100010010000000100011;
ROM[27701] <= 32'b00000000010000010000000100010011;
ROM[27702] <= 32'b00000000001100010010000000100011;
ROM[27703] <= 32'b00000000010000010000000100010011;
ROM[27704] <= 32'b00000000010000010010000000100011;
ROM[27705] <= 32'b00000000010000010000000100010011;
ROM[27706] <= 32'b00000000010100010010000000100011;
ROM[27707] <= 32'b00000000010000010000000100010011;
ROM[27708] <= 32'b00000000011000010010000000100011;
ROM[27709] <= 32'b00000000010000010000000100010011;
ROM[27710] <= 32'b00000001010000000000001110010011;
ROM[27711] <= 32'b00000000100000111000001110010011;
ROM[27712] <= 32'b01000000011100010000001110110011;
ROM[27713] <= 32'b00000000011100000000001000110011;
ROM[27714] <= 32'b00000000001000000000000110110011;
ROM[27715] <= 32'b11110010000011110110000011101111;
ROM[27716] <= 32'b11111111110000010000000100010011;
ROM[27717] <= 32'b00000000000000010010001110000011;
ROM[27718] <= 32'b11111111110000010000000100010011;
ROM[27719] <= 32'b00000000000000010010010000000011;
ROM[27720] <= 32'b00000000011101000000001110110011;
ROM[27721] <= 32'b00000000011100010010000000100011;
ROM[27722] <= 32'b00000000010000010000000100010011;
ROM[27723] <= 32'b11111111110000010000000100010011;
ROM[27724] <= 32'b00000000000000010010001110000011;
ROM[27725] <= 32'b00000000000000111000001100010011;
ROM[27726] <= 32'b00000000110100110000010000110011;
ROM[27727] <= 32'b00000000000001000010001110000011;
ROM[27728] <= 32'b00000000011100010010000000100011;
ROM[27729] <= 32'b00000000010000010000000100010011;
ROM[27730] <= 32'b11111111110000010000000100010011;
ROM[27731] <= 32'b00000000000000010010001110000011;
ROM[27732] <= 32'b00000000011100011010011000100011;
ROM[27733] <= 32'b00000000000000100010001110000011;
ROM[27734] <= 32'b00000000011100010010000000100011;
ROM[27735] <= 32'b00000000010000010000000100010011;
ROM[27736] <= 32'b00000000100000011010001110000011;
ROM[27737] <= 32'b00000000011100010010000000100011;
ROM[27738] <= 32'b00000000010000010000000100010011;
ROM[27739] <= 32'b00000000010000000000001110010011;
ROM[27740] <= 32'b00000000011100010010000000100011;
ROM[27741] <= 32'b00000000010000010000000100010011;
ROM[27742] <= 32'b00000000000000011011001110110111;
ROM[27743] <= 32'b00011100010000111000001110010011;
ROM[27744] <= 32'b00000000111000111000001110110011;
ROM[27745] <= 32'b00000000011100010010000000100011;
ROM[27746] <= 32'b00000000010000010000000100010011;
ROM[27747] <= 32'b00000000001100010010000000100011;
ROM[27748] <= 32'b00000000010000010000000100010011;
ROM[27749] <= 32'b00000000010000010010000000100011;
ROM[27750] <= 32'b00000000010000010000000100010011;
ROM[27751] <= 32'b00000000010100010010000000100011;
ROM[27752] <= 32'b00000000010000010000000100010011;
ROM[27753] <= 32'b00000000011000010010000000100011;
ROM[27754] <= 32'b00000000010000010000000100010011;
ROM[27755] <= 32'b00000001010000000000001110010011;
ROM[27756] <= 32'b00000000100000111000001110010011;
ROM[27757] <= 32'b01000000011100010000001110110011;
ROM[27758] <= 32'b00000000011100000000001000110011;
ROM[27759] <= 32'b00000000001000000000000110110011;
ROM[27760] <= 32'b11100110110011110110000011101111;
ROM[27761] <= 32'b11111111110000010000000100010011;
ROM[27762] <= 32'b00000000000000010010001110000011;
ROM[27763] <= 32'b11111111110000010000000100010011;
ROM[27764] <= 32'b00000000000000010010010000000011;
ROM[27765] <= 32'b00000000011101000000001110110011;
ROM[27766] <= 32'b00000000011100010010000000100011;
ROM[27767] <= 32'b00000000010000010000000100010011;
ROM[27768] <= 32'b11111111110000010000000100010011;
ROM[27769] <= 32'b00000000000000010010001110000011;
ROM[27770] <= 32'b00000000000000111000001100010011;
ROM[27771] <= 32'b00000000110100110000010000110011;
ROM[27772] <= 32'b00000000000001000010001110000011;
ROM[27773] <= 32'b00000000011100010010000000100011;
ROM[27774] <= 32'b00000000010000010000000100010011;
ROM[27775] <= 32'b00000000000000100010001110000011;
ROM[27776] <= 32'b00000000011100010010000000100011;
ROM[27777] <= 32'b00000000010000010000000100010011;
ROM[27778] <= 32'b00000000010000011010001110000011;
ROM[27779] <= 32'b00000000011100010010000000100011;
ROM[27780] <= 32'b00000000010000010000000100010011;
ROM[27781] <= 32'b00000000010000000000001110010011;
ROM[27782] <= 32'b00000000011100010010000000100011;
ROM[27783] <= 32'b00000000010000010000000100010011;
ROM[27784] <= 32'b00000000000000011011001110110111;
ROM[27785] <= 32'b00100110110000111000001110010011;
ROM[27786] <= 32'b00000000111000111000001110110011;
ROM[27787] <= 32'b00000000011100010010000000100011;
ROM[27788] <= 32'b00000000010000010000000100010011;
ROM[27789] <= 32'b00000000001100010010000000100011;
ROM[27790] <= 32'b00000000010000010000000100010011;
ROM[27791] <= 32'b00000000010000010010000000100011;
ROM[27792] <= 32'b00000000010000010000000100010011;
ROM[27793] <= 32'b00000000010100010010000000100011;
ROM[27794] <= 32'b00000000010000010000000100010011;
ROM[27795] <= 32'b00000000011000010010000000100011;
ROM[27796] <= 32'b00000000010000010000000100010011;
ROM[27797] <= 32'b00000001010000000000001110010011;
ROM[27798] <= 32'b00000000100000111000001110010011;
ROM[27799] <= 32'b01000000011100010000001110110011;
ROM[27800] <= 32'b00000000011100000000001000110011;
ROM[27801] <= 32'b00000000001000000000000110110011;
ROM[27802] <= 32'b11011100010011110110000011101111;
ROM[27803] <= 32'b11111111110000010000000100010011;
ROM[27804] <= 32'b00000000000000010010001110000011;
ROM[27805] <= 32'b11111111110000010000000100010011;
ROM[27806] <= 32'b00000000000000010010010000000011;
ROM[27807] <= 32'b00000000011101000000001110110011;
ROM[27808] <= 32'b00000000011100010010000000100011;
ROM[27809] <= 32'b00000000010000010000000100010011;
ROM[27810] <= 32'b11111111110000010000000100010011;
ROM[27811] <= 32'b00000000000000010010001110000011;
ROM[27812] <= 32'b00000000000000111000001100010011;
ROM[27813] <= 32'b11111111110000010000000100010011;
ROM[27814] <= 32'b00000000000000010010001110000011;
ROM[27815] <= 32'b00000000110100110000010000110011;
ROM[27816] <= 32'b00000000011101000010000000100011;
ROM[27817] <= 32'b00000000110000011010001110000011;
ROM[27818] <= 32'b00000000011100010010000000100011;
ROM[27819] <= 32'b00000000010000010000000100010011;
ROM[27820] <= 32'b00000000000000100010001110000011;
ROM[27821] <= 32'b00000000011100010010000000100011;
ROM[27822] <= 32'b00000000010000010000000100010011;
ROM[27823] <= 32'b00000000100000011010001110000011;
ROM[27824] <= 32'b00000000011100010010000000100011;
ROM[27825] <= 32'b00000000010000010000000100010011;
ROM[27826] <= 32'b00000000010000000000001110010011;
ROM[27827] <= 32'b00000000011100010010000000100011;
ROM[27828] <= 32'b00000000010000010000000100010011;
ROM[27829] <= 32'b00000000000000011011001110110111;
ROM[27830] <= 32'b00110010000000111000001110010011;
ROM[27831] <= 32'b00000000111000111000001110110011;
ROM[27832] <= 32'b00000000011100010010000000100011;
ROM[27833] <= 32'b00000000010000010000000100010011;
ROM[27834] <= 32'b00000000001100010010000000100011;
ROM[27835] <= 32'b00000000010000010000000100010011;
ROM[27836] <= 32'b00000000010000010010000000100011;
ROM[27837] <= 32'b00000000010000010000000100010011;
ROM[27838] <= 32'b00000000010100010010000000100011;
ROM[27839] <= 32'b00000000010000010000000100010011;
ROM[27840] <= 32'b00000000011000010010000000100011;
ROM[27841] <= 32'b00000000010000010000000100010011;
ROM[27842] <= 32'b00000001010000000000001110010011;
ROM[27843] <= 32'b00000000100000111000001110010011;
ROM[27844] <= 32'b01000000011100010000001110110011;
ROM[27845] <= 32'b00000000011100000000001000110011;
ROM[27846] <= 32'b00000000001000000000000110110011;
ROM[27847] <= 32'b11010001000011110110000011101111;
ROM[27848] <= 32'b11111111110000010000000100010011;
ROM[27849] <= 32'b00000000000000010010001110000011;
ROM[27850] <= 32'b11111111110000010000000100010011;
ROM[27851] <= 32'b00000000000000010010010000000011;
ROM[27852] <= 32'b00000000011101000000001110110011;
ROM[27853] <= 32'b00000000011100010010000000100011;
ROM[27854] <= 32'b00000000010000010000000100010011;
ROM[27855] <= 32'b11111111110000010000000100010011;
ROM[27856] <= 32'b00000000000000010010001110000011;
ROM[27857] <= 32'b00000000000000111000001100010011;
ROM[27858] <= 32'b11111111110000010000000100010011;
ROM[27859] <= 32'b00000000000000010010001110000011;
ROM[27860] <= 32'b00000000110100110000010000110011;
ROM[27861] <= 32'b00000000011101000010000000100011;
ROM[27862] <= 32'b00000000100000011010001110000011;
ROM[27863] <= 32'b00000000011100010010000000100011;
ROM[27864] <= 32'b00000000010000010000000100010011;
ROM[27865] <= 32'b00000000000100000000001110010011;
ROM[27866] <= 32'b00000000011100010010000000100011;
ROM[27867] <= 32'b00000000010000010000000100010011;
ROM[27868] <= 32'b11111111110000010000000100010011;
ROM[27869] <= 32'b00000000000000010010001110000011;
ROM[27870] <= 32'b11111111110000010000000100010011;
ROM[27871] <= 32'b00000000000000010010010000000011;
ROM[27872] <= 32'b00000000011101000000001110110011;
ROM[27873] <= 32'b00000000011100010010000000100011;
ROM[27874] <= 32'b00000000010000010000000100010011;
ROM[27875] <= 32'b11111111110000010000000100010011;
ROM[27876] <= 32'b00000000000000010010001110000011;
ROM[27877] <= 32'b00000000011100011010010000100011;
ROM[27878] <= 32'b10110111000111111111000011101111;
ROM[27879] <= 32'b00000000000000100010001110000011;
ROM[27880] <= 32'b00000000011100010010000000100011;
ROM[27881] <= 32'b00000000010000010000000100010011;
ROM[27882] <= 32'b00000000010000011010001110000011;
ROM[27883] <= 32'b00000000011100010010000000100011;
ROM[27884] <= 32'b00000000010000010000000100010011;
ROM[27885] <= 32'b00000000000100000000001110010011;
ROM[27886] <= 32'b00000000011100010010000000100011;
ROM[27887] <= 32'b00000000010000010000000100010011;
ROM[27888] <= 32'b11111111110000010000000100010011;
ROM[27889] <= 32'b00000000000000010010001110000011;
ROM[27890] <= 32'b11111111110000010000000100010011;
ROM[27891] <= 32'b00000000000000010010010000000011;
ROM[27892] <= 32'b00000000011101000000001110110011;
ROM[27893] <= 32'b00000000011100010010000000100011;
ROM[27894] <= 32'b00000000010000010000000100010011;
ROM[27895] <= 32'b00000000010000000000001110010011;
ROM[27896] <= 32'b00000000011100010010000000100011;
ROM[27897] <= 32'b00000000010000010000000100010011;
ROM[27898] <= 32'b00000000000000011011001110110111;
ROM[27899] <= 32'b01000011010000111000001110010011;
ROM[27900] <= 32'b00000000111000111000001110110011;
ROM[27901] <= 32'b00000000011100010010000000100011;
ROM[27902] <= 32'b00000000010000010000000100010011;
ROM[27903] <= 32'b00000000001100010010000000100011;
ROM[27904] <= 32'b00000000010000010000000100010011;
ROM[27905] <= 32'b00000000010000010010000000100011;
ROM[27906] <= 32'b00000000010000010000000100010011;
ROM[27907] <= 32'b00000000010100010010000000100011;
ROM[27908] <= 32'b00000000010000010000000100010011;
ROM[27909] <= 32'b00000000011000010010000000100011;
ROM[27910] <= 32'b00000000010000010000000100010011;
ROM[27911] <= 32'b00000001010000000000001110010011;
ROM[27912] <= 32'b00000000100000111000001110010011;
ROM[27913] <= 32'b01000000011100010000001110110011;
ROM[27914] <= 32'b00000000011100000000001000110011;
ROM[27915] <= 32'b00000000001000000000000110110011;
ROM[27916] <= 32'b10111111110011110110000011101111;
ROM[27917] <= 32'b11111111110000010000000100010011;
ROM[27918] <= 32'b00000000000000010010001110000011;
ROM[27919] <= 32'b11111111110000010000000100010011;
ROM[27920] <= 32'b00000000000000010010010000000011;
ROM[27921] <= 32'b00000000011101000000001110110011;
ROM[27922] <= 32'b00000000011100010010000000100011;
ROM[27923] <= 32'b00000000010000010000000100010011;
ROM[27924] <= 32'b11111111110000010000000100010011;
ROM[27925] <= 32'b00000000000000010010001110000011;
ROM[27926] <= 32'b00000000000000111000001100010011;
ROM[27927] <= 32'b00000000110100110000010000110011;
ROM[27928] <= 32'b00000000000001000010001110000011;
ROM[27929] <= 32'b00000000011100010010000000100011;
ROM[27930] <= 32'b00000000010000010000000100010011;
ROM[27931] <= 32'b11111111110000010000000100010011;
ROM[27932] <= 32'b00000000000000010010001110000011;
ROM[27933] <= 32'b00000000011100011010011000100011;
ROM[27934] <= 32'b00000000000000100010001110000011;
ROM[27935] <= 32'b00000000011100010010000000100011;
ROM[27936] <= 32'b00000000010000010000000100010011;
ROM[27937] <= 32'b00000000100000100010001110000011;
ROM[27938] <= 32'b00000000011100010010000000100011;
ROM[27939] <= 32'b00000000010000010000000100010011;
ROM[27940] <= 32'b00000000010000000000001110010011;
ROM[27941] <= 32'b00000000011100010010000000100011;
ROM[27942] <= 32'b00000000010000010000000100010011;
ROM[27943] <= 32'b00000000000000011011001110110111;
ROM[27944] <= 32'b01001110100000111000001110010011;
ROM[27945] <= 32'b00000000111000111000001110110011;
ROM[27946] <= 32'b00000000011100010010000000100011;
ROM[27947] <= 32'b00000000010000010000000100010011;
ROM[27948] <= 32'b00000000001100010010000000100011;
ROM[27949] <= 32'b00000000010000010000000100010011;
ROM[27950] <= 32'b00000000010000010010000000100011;
ROM[27951] <= 32'b00000000010000010000000100010011;
ROM[27952] <= 32'b00000000010100010010000000100011;
ROM[27953] <= 32'b00000000010000010000000100010011;
ROM[27954] <= 32'b00000000011000010010000000100011;
ROM[27955] <= 32'b00000000010000010000000100010011;
ROM[27956] <= 32'b00000001010000000000001110010011;
ROM[27957] <= 32'b00000000100000111000001110010011;
ROM[27958] <= 32'b01000000011100010000001110110011;
ROM[27959] <= 32'b00000000011100000000001000110011;
ROM[27960] <= 32'b00000000001000000000000110110011;
ROM[27961] <= 32'b10110100100011110110000011101111;
ROM[27962] <= 32'b11111111110000010000000100010011;
ROM[27963] <= 32'b00000000000000010010001110000011;
ROM[27964] <= 32'b11111111110000010000000100010011;
ROM[27965] <= 32'b00000000000000010010010000000011;
ROM[27966] <= 32'b00000000011101000000001110110011;
ROM[27967] <= 32'b00000000011100010010000000100011;
ROM[27968] <= 32'b00000000010000010000000100010011;
ROM[27969] <= 32'b11111111110000010000000100010011;
ROM[27970] <= 32'b00000000000000010010001110000011;
ROM[27971] <= 32'b00000000000000111000001100010011;
ROM[27972] <= 32'b00000000110100110000010000110011;
ROM[27973] <= 32'b00000000000001000010001110000011;
ROM[27974] <= 32'b00000000011100010010000000100011;
ROM[27975] <= 32'b00000000010000010000000100010011;
ROM[27976] <= 32'b00000000000000100010001110000011;
ROM[27977] <= 32'b00000000011100010010000000100011;
ROM[27978] <= 32'b00000000010000010000000100010011;
ROM[27979] <= 32'b00000000010000011010001110000011;
ROM[27980] <= 32'b00000000011100010010000000100011;
ROM[27981] <= 32'b00000000010000010000000100010011;
ROM[27982] <= 32'b00000000000100000000001110010011;
ROM[27983] <= 32'b00000000011100010010000000100011;
ROM[27984] <= 32'b00000000010000010000000100010011;
ROM[27985] <= 32'b11111111110000010000000100010011;
ROM[27986] <= 32'b00000000000000010010001110000011;
ROM[27987] <= 32'b11111111110000010000000100010011;
ROM[27988] <= 32'b00000000000000010010010000000011;
ROM[27989] <= 32'b00000000011101000000001110110011;
ROM[27990] <= 32'b00000000011100010010000000100011;
ROM[27991] <= 32'b00000000010000010000000100010011;
ROM[27992] <= 32'b00000000010000000000001110010011;
ROM[27993] <= 32'b00000000011100010010000000100011;
ROM[27994] <= 32'b00000000010000010000000100010011;
ROM[27995] <= 32'b00000000000000011011001110110111;
ROM[27996] <= 32'b01011011100000111000001110010011;
ROM[27997] <= 32'b00000000111000111000001110110011;
ROM[27998] <= 32'b00000000011100010010000000100011;
ROM[27999] <= 32'b00000000010000010000000100010011;
ROM[28000] <= 32'b00000000001100010010000000100011;
ROM[28001] <= 32'b00000000010000010000000100010011;
ROM[28002] <= 32'b00000000010000010010000000100011;
ROM[28003] <= 32'b00000000010000010000000100010011;
ROM[28004] <= 32'b00000000010100010010000000100011;
ROM[28005] <= 32'b00000000010000010000000100010011;
ROM[28006] <= 32'b00000000011000010010000000100011;
ROM[28007] <= 32'b00000000010000010000000100010011;
ROM[28008] <= 32'b00000001010000000000001110010011;
ROM[28009] <= 32'b00000000100000111000001110010011;
ROM[28010] <= 32'b01000000011100010000001110110011;
ROM[28011] <= 32'b00000000011100000000001000110011;
ROM[28012] <= 32'b00000000001000000000000110110011;
ROM[28013] <= 32'b10100111100011110110000011101111;
ROM[28014] <= 32'b11111111110000010000000100010011;
ROM[28015] <= 32'b00000000000000010010001110000011;
ROM[28016] <= 32'b11111111110000010000000100010011;
ROM[28017] <= 32'b00000000000000010010010000000011;
ROM[28018] <= 32'b00000000011101000000001110110011;
ROM[28019] <= 32'b00000000011100010010000000100011;
ROM[28020] <= 32'b00000000010000010000000100010011;
ROM[28021] <= 32'b11111111110000010000000100010011;
ROM[28022] <= 32'b00000000000000010010001110000011;
ROM[28023] <= 32'b00000000000000111000001100010011;
ROM[28024] <= 32'b11111111110000010000000100010011;
ROM[28025] <= 32'b00000000000000010010001110000011;
ROM[28026] <= 32'b00000000110100110000010000110011;
ROM[28027] <= 32'b00000000011101000010000000100011;
ROM[28028] <= 32'b00000000110000011010001110000011;
ROM[28029] <= 32'b00000000011100010010000000100011;
ROM[28030] <= 32'b00000000010000010000000100010011;
ROM[28031] <= 32'b00000000000000100010001110000011;
ROM[28032] <= 32'b00000000011100010010000000100011;
ROM[28033] <= 32'b00000000010000010000000100010011;
ROM[28034] <= 32'b00000000100000100010001110000011;
ROM[28035] <= 32'b00000000011100010010000000100011;
ROM[28036] <= 32'b00000000010000010000000100010011;
ROM[28037] <= 32'b00000000010000000000001110010011;
ROM[28038] <= 32'b00000000011100010010000000100011;
ROM[28039] <= 32'b00000000010000010000000100010011;
ROM[28040] <= 32'b00000000000000011011001110110111;
ROM[28041] <= 32'b01100110110000111000001110010011;
ROM[28042] <= 32'b00000000111000111000001110110011;
ROM[28043] <= 32'b00000000011100010010000000100011;
ROM[28044] <= 32'b00000000010000010000000100010011;
ROM[28045] <= 32'b00000000001100010010000000100011;
ROM[28046] <= 32'b00000000010000010000000100010011;
ROM[28047] <= 32'b00000000010000010010000000100011;
ROM[28048] <= 32'b00000000010000010000000100010011;
ROM[28049] <= 32'b00000000010100010010000000100011;
ROM[28050] <= 32'b00000000010000010000000100010011;
ROM[28051] <= 32'b00000000011000010010000000100011;
ROM[28052] <= 32'b00000000010000010000000100010011;
ROM[28053] <= 32'b00000001010000000000001110010011;
ROM[28054] <= 32'b00000000100000111000001110010011;
ROM[28055] <= 32'b01000000011100010000001110110011;
ROM[28056] <= 32'b00000000011100000000001000110011;
ROM[28057] <= 32'b00000000001000000000000110110011;
ROM[28058] <= 32'b10011100010011110110000011101111;
ROM[28059] <= 32'b11111111110000010000000100010011;
ROM[28060] <= 32'b00000000000000010010001110000011;
ROM[28061] <= 32'b11111111110000010000000100010011;
ROM[28062] <= 32'b00000000000000010010010000000011;
ROM[28063] <= 32'b00000000011101000000001110110011;
ROM[28064] <= 32'b00000000011100010010000000100011;
ROM[28065] <= 32'b00000000010000010000000100010011;
ROM[28066] <= 32'b11111111110000010000000100010011;
ROM[28067] <= 32'b00000000000000010010001110000011;
ROM[28068] <= 32'b00000000000000111000001100010011;
ROM[28069] <= 32'b11111111110000010000000100010011;
ROM[28070] <= 32'b00000000000000010010001110000011;
ROM[28071] <= 32'b00000000110100110000010000110011;
ROM[28072] <= 32'b00000000011101000010000000100011;
ROM[28073] <= 32'b00000000010000011010001110000011;
ROM[28074] <= 32'b00000000011100010010000000100011;
ROM[28075] <= 32'b00000000010000010000000100010011;
ROM[28076] <= 32'b00000000000100000000001110010011;
ROM[28077] <= 32'b00000000011100010010000000100011;
ROM[28078] <= 32'b00000000010000010000000100010011;
ROM[28079] <= 32'b11111111110000010000000100010011;
ROM[28080] <= 32'b00000000000000010010001110000011;
ROM[28081] <= 32'b11111111110000010000000100010011;
ROM[28082] <= 32'b00000000000000010010010000000011;
ROM[28083] <= 32'b00000000011101000000001110110011;
ROM[28084] <= 32'b00000000011100010010000000100011;
ROM[28085] <= 32'b00000000010000010000000100010011;
ROM[28086] <= 32'b00000001010000000000001110010011;
ROM[28087] <= 32'b01000000011100011000001110110011;
ROM[28088] <= 32'b00000000000000111010000010000011;
ROM[28089] <= 32'b11111111110000010000000100010011;
ROM[28090] <= 32'b00000000000000010010001110000011;
ROM[28091] <= 32'b00000000011100100010000000100011;
ROM[28092] <= 32'b00000000010000100000000100010011;
ROM[28093] <= 32'b00000001010000000000001110010011;
ROM[28094] <= 32'b01000000011100011000001110110011;
ROM[28095] <= 32'b00000000010000111010000110000011;
ROM[28096] <= 32'b00000000100000111010001000000011;
ROM[28097] <= 32'b00000000110000111010001010000011;
ROM[28098] <= 32'b00000001000000111010001100000011;
ROM[28099] <= 32'b00000000000000001000000011100111;
ROM[28100] <= 32'b00000000000000010010000000100011;
ROM[28101] <= 32'b00000000010000010000000100010011;
ROM[28102] <= 32'b00000000000000010010000000100011;
ROM[28103] <= 32'b00000000010000010000000100010011;
ROM[28104] <= 32'b00000000000100000000001110010011;
ROM[28105] <= 32'b00000000011100010010000000100011;
ROM[28106] <= 32'b00000000010000010000000100010011;
ROM[28107] <= 32'b11111111110000010000000100010011;
ROM[28108] <= 32'b00000000000000010010001110000011;
ROM[28109] <= 32'b00000000011100011010000000100011;
ROM[28110] <= 32'b00000000000000011011001110110111;
ROM[28111] <= 32'b01111000010000111000001110010011;
ROM[28112] <= 32'b00000000111000111000001110110011;
ROM[28113] <= 32'b00000000011100010010000000100011;
ROM[28114] <= 32'b00000000010000010000000100010011;
ROM[28115] <= 32'b00000000001100010010000000100011;
ROM[28116] <= 32'b00000000010000010000000100010011;
ROM[28117] <= 32'b00000000010000010010000000100011;
ROM[28118] <= 32'b00000000010000010000000100010011;
ROM[28119] <= 32'b00000000010100010010000000100011;
ROM[28120] <= 32'b00000000010000010000000100010011;
ROM[28121] <= 32'b00000000011000010010000000100011;
ROM[28122] <= 32'b00000000010000010000000100010011;
ROM[28123] <= 32'b00000001010000000000001110010011;
ROM[28124] <= 32'b00000000000000111000001110010011;
ROM[28125] <= 32'b01000000011100010000001110110011;
ROM[28126] <= 32'b00000000011100000000001000110011;
ROM[28127] <= 32'b00000000001000000000000110110011;
ROM[28128] <= 32'b11001011110111111100000011101111;
ROM[28129] <= 32'b11111111110000010000000100010011;
ROM[28130] <= 32'b00000000000000010010001110000011;
ROM[28131] <= 32'b00000000011101100010000000100011;
ROM[28132] <= 32'b00000000000000011010001110000011;
ROM[28133] <= 32'b00000000011100010010000000100011;
ROM[28134] <= 32'b00000000010000010000000100010011;
ROM[28135] <= 32'b00000000000100000000001110010011;
ROM[28136] <= 32'b00000000011100010010000000100011;
ROM[28137] <= 32'b00000000010000010000000100010011;
ROM[28138] <= 32'b11111111110000010000000100010011;
ROM[28139] <= 32'b00000000000000010010001110000011;
ROM[28140] <= 32'b11111111110000010000000100010011;
ROM[28141] <= 32'b00000000000000010010010000000011;
ROM[28142] <= 32'b00000000011101000010010010110011;
ROM[28143] <= 32'b00000000100000111010010100110011;
ROM[28144] <= 32'b00000000101001001000001110110011;
ROM[28145] <= 32'b00000000000100111000001110010011;
ROM[28146] <= 32'b00000000000100111111001110010011;
ROM[28147] <= 32'b00000000011100010010000000100011;
ROM[28148] <= 32'b00000000010000010000000100010011;
ROM[28149] <= 32'b11111111110000010000000100010011;
ROM[28150] <= 32'b00000000000000010010001110000011;
ROM[28151] <= 32'b01000000011100000000001110110011;
ROM[28152] <= 32'b00000000000100111000001110010011;
ROM[28153] <= 32'b00000000011100010010000000100011;
ROM[28154] <= 32'b00000000010000010000000100010011;
ROM[28155] <= 32'b11111111110000010000000100010011;
ROM[28156] <= 32'b00000000000000010010001110000011;
ROM[28157] <= 32'b00000000000000111000101001100011;
ROM[28158] <= 32'b00000000000000011101001110110111;
ROM[28159] <= 32'b11011000000000111000001110010011;
ROM[28160] <= 32'b00000000111000111000001110110011;
ROM[28161] <= 32'b00000000000000111000000011100111;
ROM[28162] <= 32'b00000000000000011100001110110111;
ROM[28163] <= 32'b10000101010000111000001110010011;
ROM[28164] <= 32'b00000000111000111000001110110011;
ROM[28165] <= 32'b00000000011100010010000000100011;
ROM[28166] <= 32'b00000000010000010000000100010011;
ROM[28167] <= 32'b00000000001100010010000000100011;
ROM[28168] <= 32'b00000000010000010000000100010011;
ROM[28169] <= 32'b00000000010000010010000000100011;
ROM[28170] <= 32'b00000000010000010000000100010011;
ROM[28171] <= 32'b00000000010100010010000000100011;
ROM[28172] <= 32'b00000000010000010000000100010011;
ROM[28173] <= 32'b00000000011000010010000000100011;
ROM[28174] <= 32'b00000000010000010000000100010011;
ROM[28175] <= 32'b00000001010000000000001110010011;
ROM[28176] <= 32'b00000000000000111000001110010011;
ROM[28177] <= 32'b01000000011100010000001110110011;
ROM[28178] <= 32'b00000000011100000000001000110011;
ROM[28179] <= 32'b00000000001000000000000110110011;
ROM[28180] <= 32'b10110001100111111011000011101111;
ROM[28181] <= 32'b11111111110000010000000100010011;
ROM[28182] <= 32'b00000000000000010010001110000011;
ROM[28183] <= 32'b00000000011101100010000000100011;
ROM[28184] <= 32'b00000010100100000000001110010011;
ROM[28185] <= 32'b00000000011100010010000000100011;
ROM[28186] <= 32'b00000000010000010000000100010011;
ROM[28187] <= 32'b00000000000000011100001110110111;
ROM[28188] <= 32'b10001011100000111000001110010011;
ROM[28189] <= 32'b00000000111000111000001110110011;
ROM[28190] <= 32'b00000000011100010010000000100011;
ROM[28191] <= 32'b00000000010000010000000100010011;
ROM[28192] <= 32'b00000000001100010010000000100011;
ROM[28193] <= 32'b00000000010000010000000100010011;
ROM[28194] <= 32'b00000000010000010010000000100011;
ROM[28195] <= 32'b00000000010000010000000100010011;
ROM[28196] <= 32'b00000000010100010010000000100011;
ROM[28197] <= 32'b00000000010000010000000100010011;
ROM[28198] <= 32'b00000000011000010010000000100011;
ROM[28199] <= 32'b00000000010000010000000100010011;
ROM[28200] <= 32'b00000001010000000000001110010011;
ROM[28201] <= 32'b00000000010000111000001110010011;
ROM[28202] <= 32'b01000000011100010000001110110011;
ROM[28203] <= 32'b00000000011100000000001000110011;
ROM[28204] <= 32'b00000000001000000000000110110011;
ROM[28205] <= 32'b01101000100100001101000011101111;
ROM[28206] <= 32'b00000100010000000000001110010011;
ROM[28207] <= 32'b00000000011100010010000000100011;
ROM[28208] <= 32'b00000000010000010000000100010011;
ROM[28209] <= 32'b00000000000000011100001110110111;
ROM[28210] <= 32'b10010001000000111000001110010011;
ROM[28211] <= 32'b00000000111000111000001110110011;
ROM[28212] <= 32'b00000000011100010010000000100011;
ROM[28213] <= 32'b00000000010000010000000100010011;
ROM[28214] <= 32'b00000000001100010010000000100011;
ROM[28215] <= 32'b00000000010000010000000100010011;
ROM[28216] <= 32'b00000000010000010010000000100011;
ROM[28217] <= 32'b00000000010000010000000100010011;
ROM[28218] <= 32'b00000000010100010010000000100011;
ROM[28219] <= 32'b00000000010000010000000100010011;
ROM[28220] <= 32'b00000000011000010010000000100011;
ROM[28221] <= 32'b00000000010000010000000100010011;
ROM[28222] <= 32'b00000001010000000000001110010011;
ROM[28223] <= 32'b00000000100000111000001110010011;
ROM[28224] <= 32'b01000000011100010000001110110011;
ROM[28225] <= 32'b00000000011100000000001000110011;
ROM[28226] <= 32'b00000000001000000000000110110011;
ROM[28227] <= 32'b00101010000000001110000011101111;
ROM[28228] <= 32'b00000110111100000000001110010011;
ROM[28229] <= 32'b00000000011100010010000000100011;
ROM[28230] <= 32'b00000000010000010000000100010011;
ROM[28231] <= 32'b00000000000000011100001110110111;
ROM[28232] <= 32'b10010110100000111000001110010011;
ROM[28233] <= 32'b00000000111000111000001110110011;
ROM[28234] <= 32'b00000000011100010010000000100011;
ROM[28235] <= 32'b00000000010000010000000100010011;
ROM[28236] <= 32'b00000000001100010010000000100011;
ROM[28237] <= 32'b00000000010000010000000100010011;
ROM[28238] <= 32'b00000000010000010010000000100011;
ROM[28239] <= 32'b00000000010000010000000100010011;
ROM[28240] <= 32'b00000000010100010010000000100011;
ROM[28241] <= 32'b00000000010000010000000100010011;
ROM[28242] <= 32'b00000000011000010010000000100011;
ROM[28243] <= 32'b00000000010000010000000100010011;
ROM[28244] <= 32'b00000001010000000000001110010011;
ROM[28245] <= 32'b00000000100000111000001110010011;
ROM[28246] <= 32'b01000000011100010000001110110011;
ROM[28247] <= 32'b00000000011100000000001000110011;
ROM[28248] <= 32'b00000000001000000000000110110011;
ROM[28249] <= 32'b00100100100000001110000011101111;
ROM[28250] <= 32'b00000010000000000000001110010011;
ROM[28251] <= 32'b00000000011100010010000000100011;
ROM[28252] <= 32'b00000000010000010000000100010011;
ROM[28253] <= 32'b00000000000000011100001110110111;
ROM[28254] <= 32'b10011100000000111000001110010011;
ROM[28255] <= 32'b00000000111000111000001110110011;
ROM[28256] <= 32'b00000000011100010010000000100011;
ROM[28257] <= 32'b00000000010000010000000100010011;
ROM[28258] <= 32'b00000000001100010010000000100011;
ROM[28259] <= 32'b00000000010000010000000100010011;
ROM[28260] <= 32'b00000000010000010010000000100011;
ROM[28261] <= 32'b00000000010000010000000100010011;
ROM[28262] <= 32'b00000000010100010010000000100011;
ROM[28263] <= 32'b00000000010000010000000100010011;
ROM[28264] <= 32'b00000000011000010010000000100011;
ROM[28265] <= 32'b00000000010000010000000100010011;
ROM[28266] <= 32'b00000001010000000000001110010011;
ROM[28267] <= 32'b00000000100000111000001110010011;
ROM[28268] <= 32'b01000000011100010000001110110011;
ROM[28269] <= 32'b00000000011100000000001000110011;
ROM[28270] <= 32'b00000000001000000000000110110011;
ROM[28271] <= 32'b00011111000000001110000011101111;
ROM[28272] <= 32'b00000111100100000000001110010011;
ROM[28273] <= 32'b00000000011100010010000000100011;
ROM[28274] <= 32'b00000000010000010000000100010011;
ROM[28275] <= 32'b00000000000000011100001110110111;
ROM[28276] <= 32'b10100001100000111000001110010011;
ROM[28277] <= 32'b00000000111000111000001110110011;
ROM[28278] <= 32'b00000000011100010010000000100011;
ROM[28279] <= 32'b00000000010000010000000100010011;
ROM[28280] <= 32'b00000000001100010010000000100011;
ROM[28281] <= 32'b00000000010000010000000100010011;
ROM[28282] <= 32'b00000000010000010010000000100011;
ROM[28283] <= 32'b00000000010000010000000100010011;
ROM[28284] <= 32'b00000000010100010010000000100011;
ROM[28285] <= 32'b00000000010000010000000100010011;
ROM[28286] <= 32'b00000000011000010010000000100011;
ROM[28287] <= 32'b00000000010000010000000100010011;
ROM[28288] <= 32'b00000001010000000000001110010011;
ROM[28289] <= 32'b00000000100000111000001110010011;
ROM[28290] <= 32'b01000000011100010000001110110011;
ROM[28291] <= 32'b00000000011100000000001000110011;
ROM[28292] <= 32'b00000000001000000000000110110011;
ROM[28293] <= 32'b00011001100000001110000011101111;
ROM[28294] <= 32'b00000110111100000000001110010011;
ROM[28295] <= 32'b00000000011100010010000000100011;
ROM[28296] <= 32'b00000000010000010000000100010011;
ROM[28297] <= 32'b00000000000000011100001110110111;
ROM[28298] <= 32'b10100111000000111000001110010011;
ROM[28299] <= 32'b00000000111000111000001110110011;
ROM[28300] <= 32'b00000000011100010010000000100011;
ROM[28301] <= 32'b00000000010000010000000100010011;
ROM[28302] <= 32'b00000000001100010010000000100011;
ROM[28303] <= 32'b00000000010000010000000100010011;
ROM[28304] <= 32'b00000000010000010010000000100011;
ROM[28305] <= 32'b00000000010000010000000100010011;
ROM[28306] <= 32'b00000000010100010010000000100011;
ROM[28307] <= 32'b00000000010000010000000100010011;
ROM[28308] <= 32'b00000000011000010010000000100011;
ROM[28309] <= 32'b00000000010000010000000100010011;
ROM[28310] <= 32'b00000001010000000000001110010011;
ROM[28311] <= 32'b00000000100000111000001110010011;
ROM[28312] <= 32'b01000000011100010000001110110011;
ROM[28313] <= 32'b00000000011100000000001000110011;
ROM[28314] <= 32'b00000000001000000000000110110011;
ROM[28315] <= 32'b00010100000000001110000011101111;
ROM[28316] <= 32'b00000111010100000000001110010011;
ROM[28317] <= 32'b00000000011100010010000000100011;
ROM[28318] <= 32'b00000000010000010000000100010011;
ROM[28319] <= 32'b00000000000000011100001110110111;
ROM[28320] <= 32'b10101100100000111000001110010011;
ROM[28321] <= 32'b00000000111000111000001110110011;
ROM[28322] <= 32'b00000000011100010010000000100011;
ROM[28323] <= 32'b00000000010000010000000100010011;
ROM[28324] <= 32'b00000000001100010010000000100011;
ROM[28325] <= 32'b00000000010000010000000100010011;
ROM[28326] <= 32'b00000000010000010010000000100011;
ROM[28327] <= 32'b00000000010000010000000100010011;
ROM[28328] <= 32'b00000000010100010010000000100011;
ROM[28329] <= 32'b00000000010000010000000100010011;
ROM[28330] <= 32'b00000000011000010010000000100011;
ROM[28331] <= 32'b00000000010000010000000100010011;
ROM[28332] <= 32'b00000001010000000000001110010011;
ROM[28333] <= 32'b00000000100000111000001110010011;
ROM[28334] <= 32'b01000000011100010000001110110011;
ROM[28335] <= 32'b00000000011100000000001000110011;
ROM[28336] <= 32'b00000000001000000000000110110011;
ROM[28337] <= 32'b00001110100000001110000011101111;
ROM[28338] <= 32'b00000010000000000000001110010011;
ROM[28339] <= 32'b00000000011100010010000000100011;
ROM[28340] <= 32'b00000000010000010000000100010011;
ROM[28341] <= 32'b00000000000000011100001110110111;
ROM[28342] <= 32'b10110010000000111000001110010011;
ROM[28343] <= 32'b00000000111000111000001110110011;
ROM[28344] <= 32'b00000000011100010010000000100011;
ROM[28345] <= 32'b00000000010000010000000100010011;
ROM[28346] <= 32'b00000000001100010010000000100011;
ROM[28347] <= 32'b00000000010000010000000100010011;
ROM[28348] <= 32'b00000000010000010010000000100011;
ROM[28349] <= 32'b00000000010000010000000100010011;
ROM[28350] <= 32'b00000000010100010010000000100011;
ROM[28351] <= 32'b00000000010000010000000100010011;
ROM[28352] <= 32'b00000000011000010010000000100011;
ROM[28353] <= 32'b00000000010000010000000100010011;
ROM[28354] <= 32'b00000001010000000000001110010011;
ROM[28355] <= 32'b00000000100000111000001110010011;
ROM[28356] <= 32'b01000000011100010000001110110011;
ROM[28357] <= 32'b00000000011100000000001000110011;
ROM[28358] <= 32'b00000000001000000000000110110011;
ROM[28359] <= 32'b00001001000000001110000011101111;
ROM[28360] <= 32'b00000111011100000000001110010011;
ROM[28361] <= 32'b00000000011100010010000000100011;
ROM[28362] <= 32'b00000000010000010000000100010011;
ROM[28363] <= 32'b00000000000000011100001110110111;
ROM[28364] <= 32'b10110111100000111000001110010011;
ROM[28365] <= 32'b00000000111000111000001110110011;
ROM[28366] <= 32'b00000000011100010010000000100011;
ROM[28367] <= 32'b00000000010000010000000100010011;
ROM[28368] <= 32'b00000000001100010010000000100011;
ROM[28369] <= 32'b00000000010000010000000100010011;
ROM[28370] <= 32'b00000000010000010010000000100011;
ROM[28371] <= 32'b00000000010000010000000100010011;
ROM[28372] <= 32'b00000000010100010010000000100011;
ROM[28373] <= 32'b00000000010000010000000100010011;
ROM[28374] <= 32'b00000000011000010010000000100011;
ROM[28375] <= 32'b00000000010000010000000100010011;
ROM[28376] <= 32'b00000001010000000000001110010011;
ROM[28377] <= 32'b00000000100000111000001110010011;
ROM[28378] <= 32'b01000000011100010000001110110011;
ROM[28379] <= 32'b00000000011100000000001000110011;
ROM[28380] <= 32'b00000000001000000000000110110011;
ROM[28381] <= 32'b00000011100000001110000011101111;
ROM[28382] <= 32'b00000110000100000000001110010011;
ROM[28383] <= 32'b00000000011100010010000000100011;
ROM[28384] <= 32'b00000000010000010000000100010011;
ROM[28385] <= 32'b00000000000000011100001110110111;
ROM[28386] <= 32'b10111101000000111000001110010011;
ROM[28387] <= 32'b00000000111000111000001110110011;
ROM[28388] <= 32'b00000000011100010010000000100011;
ROM[28389] <= 32'b00000000010000010000000100010011;
ROM[28390] <= 32'b00000000001100010010000000100011;
ROM[28391] <= 32'b00000000010000010000000100010011;
ROM[28392] <= 32'b00000000010000010010000000100011;
ROM[28393] <= 32'b00000000010000010000000100010011;
ROM[28394] <= 32'b00000000010100010010000000100011;
ROM[28395] <= 32'b00000000010000010000000100010011;
ROM[28396] <= 32'b00000000011000010010000000100011;
ROM[28397] <= 32'b00000000010000010000000100010011;
ROM[28398] <= 32'b00000001010000000000001110010011;
ROM[28399] <= 32'b00000000100000111000001110010011;
ROM[28400] <= 32'b01000000011100010000001110110011;
ROM[28401] <= 32'b00000000011100000000001000110011;
ROM[28402] <= 32'b00000000001000000000000110110011;
ROM[28403] <= 32'b01111110000100001101000011101111;
ROM[28404] <= 32'b00000110111000000000001110010011;
ROM[28405] <= 32'b00000000011100010010000000100011;
ROM[28406] <= 32'b00000000010000010000000100010011;
ROM[28407] <= 32'b00000000000000011100001110110111;
ROM[28408] <= 32'b11000010100000111000001110010011;
ROM[28409] <= 32'b00000000111000111000001110110011;
ROM[28410] <= 32'b00000000011100010010000000100011;
ROM[28411] <= 32'b00000000010000010000000100010011;
ROM[28412] <= 32'b00000000001100010010000000100011;
ROM[28413] <= 32'b00000000010000010000000100010011;
ROM[28414] <= 32'b00000000010000010010000000100011;
ROM[28415] <= 32'b00000000010000010000000100010011;
ROM[28416] <= 32'b00000000010100010010000000100011;
ROM[28417] <= 32'b00000000010000010000000100010011;
ROM[28418] <= 32'b00000000011000010010000000100011;
ROM[28419] <= 32'b00000000010000010000000100010011;
ROM[28420] <= 32'b00000001010000000000001110010011;
ROM[28421] <= 32'b00000000100000111000001110010011;
ROM[28422] <= 32'b01000000011100010000001110110011;
ROM[28423] <= 32'b00000000011100000000001000110011;
ROM[28424] <= 32'b00000000001000000000000110110011;
ROM[28425] <= 32'b01111000100100001101000011101111;
ROM[28426] <= 32'b00000111010000000000001110010011;
ROM[28427] <= 32'b00000000011100010010000000100011;
ROM[28428] <= 32'b00000000010000010000000100010011;
ROM[28429] <= 32'b00000000000000011100001110110111;
ROM[28430] <= 32'b11001000000000111000001110010011;
ROM[28431] <= 32'b00000000111000111000001110110011;
ROM[28432] <= 32'b00000000011100010010000000100011;
ROM[28433] <= 32'b00000000010000010000000100010011;
ROM[28434] <= 32'b00000000001100010010000000100011;
ROM[28435] <= 32'b00000000010000010000000100010011;
ROM[28436] <= 32'b00000000010000010010000000100011;
ROM[28437] <= 32'b00000000010000010000000100010011;
ROM[28438] <= 32'b00000000010100010010000000100011;
ROM[28439] <= 32'b00000000010000010000000100010011;
ROM[28440] <= 32'b00000000011000010010000000100011;
ROM[28441] <= 32'b00000000010000010000000100010011;
ROM[28442] <= 32'b00000001010000000000001110010011;
ROM[28443] <= 32'b00000000100000111000001110010011;
ROM[28444] <= 32'b01000000011100010000001110110011;
ROM[28445] <= 32'b00000000011100000000001000110011;
ROM[28446] <= 32'b00000000001000000000000110110011;
ROM[28447] <= 32'b01110011000100001101000011101111;
ROM[28448] <= 32'b00000010000000000000001110010011;
ROM[28449] <= 32'b00000000011100010010000000100011;
ROM[28450] <= 32'b00000000010000010000000100010011;
ROM[28451] <= 32'b00000000000000011100001110110111;
ROM[28452] <= 32'b11001101100000111000001110010011;
ROM[28453] <= 32'b00000000111000111000001110110011;
ROM[28454] <= 32'b00000000011100010010000000100011;
ROM[28455] <= 32'b00000000010000010000000100010011;
ROM[28456] <= 32'b00000000001100010010000000100011;
ROM[28457] <= 32'b00000000010000010000000100010011;
ROM[28458] <= 32'b00000000010000010010000000100011;
ROM[28459] <= 32'b00000000010000010000000100010011;
ROM[28460] <= 32'b00000000010100010010000000100011;
ROM[28461] <= 32'b00000000010000010000000100010011;
ROM[28462] <= 32'b00000000011000010010000000100011;
ROM[28463] <= 32'b00000000010000010000000100010011;
ROM[28464] <= 32'b00000001010000000000001110010011;
ROM[28465] <= 32'b00000000100000111000001110010011;
ROM[28466] <= 32'b01000000011100010000001110110011;
ROM[28467] <= 32'b00000000011100000000001000110011;
ROM[28468] <= 32'b00000000001000000000000110110011;
ROM[28469] <= 32'b01101101100100001101000011101111;
ROM[28470] <= 32'b00000111010000000000001110010011;
ROM[28471] <= 32'b00000000011100010010000000100011;
ROM[28472] <= 32'b00000000010000010000000100010011;
ROM[28473] <= 32'b00000000000000011100001110110111;
ROM[28474] <= 32'b11010011000000111000001110010011;
ROM[28475] <= 32'b00000000111000111000001110110011;
ROM[28476] <= 32'b00000000011100010010000000100011;
ROM[28477] <= 32'b00000000010000010000000100010011;
ROM[28478] <= 32'b00000000001100010010000000100011;
ROM[28479] <= 32'b00000000010000010000000100010011;
ROM[28480] <= 32'b00000000010000010010000000100011;
ROM[28481] <= 32'b00000000010000010000000100010011;
ROM[28482] <= 32'b00000000010100010010000000100011;
ROM[28483] <= 32'b00000000010000010000000100010011;
ROM[28484] <= 32'b00000000011000010010000000100011;
ROM[28485] <= 32'b00000000010000010000000100010011;
ROM[28486] <= 32'b00000001010000000000001110010011;
ROM[28487] <= 32'b00000000100000111000001110010011;
ROM[28488] <= 32'b01000000011100010000001110110011;
ROM[28489] <= 32'b00000000011100000000001000110011;
ROM[28490] <= 32'b00000000001000000000000110110011;
ROM[28491] <= 32'b01101000000100001101000011101111;
ROM[28492] <= 32'b00000110111100000000001110010011;
ROM[28493] <= 32'b00000000011100010010000000100011;
ROM[28494] <= 32'b00000000010000010000000100010011;
ROM[28495] <= 32'b00000000000000011100001110110111;
ROM[28496] <= 32'b11011000100000111000001110010011;
ROM[28497] <= 32'b00000000111000111000001110110011;
ROM[28498] <= 32'b00000000011100010010000000100011;
ROM[28499] <= 32'b00000000010000010000000100010011;
ROM[28500] <= 32'b00000000001100010010000000100011;
ROM[28501] <= 32'b00000000010000010000000100010011;
ROM[28502] <= 32'b00000000010000010010000000100011;
ROM[28503] <= 32'b00000000010000010000000100010011;
ROM[28504] <= 32'b00000000010100010010000000100011;
ROM[28505] <= 32'b00000000010000010000000100010011;
ROM[28506] <= 32'b00000000011000010010000000100011;
ROM[28507] <= 32'b00000000010000010000000100010011;
ROM[28508] <= 32'b00000001010000000000001110010011;
ROM[28509] <= 32'b00000000100000111000001110010011;
ROM[28510] <= 32'b01000000011100010000001110110011;
ROM[28511] <= 32'b00000000011100000000001000110011;
ROM[28512] <= 32'b00000000001000000000000110110011;
ROM[28513] <= 32'b01100010100100001101000011101111;
ROM[28514] <= 32'b00000010000000000000001110010011;
ROM[28515] <= 32'b00000000011100010010000000100011;
ROM[28516] <= 32'b00000000010000010000000100010011;
ROM[28517] <= 32'b00000000000000011100001110110111;
ROM[28518] <= 32'b11011110000000111000001110010011;
ROM[28519] <= 32'b00000000111000111000001110110011;
ROM[28520] <= 32'b00000000011100010010000000100011;
ROM[28521] <= 32'b00000000010000010000000100010011;
ROM[28522] <= 32'b00000000001100010010000000100011;
ROM[28523] <= 32'b00000000010000010000000100010011;
ROM[28524] <= 32'b00000000010000010010000000100011;
ROM[28525] <= 32'b00000000010000010000000100010011;
ROM[28526] <= 32'b00000000010100010010000000100011;
ROM[28527] <= 32'b00000000010000010000000100010011;
ROM[28528] <= 32'b00000000011000010010000000100011;
ROM[28529] <= 32'b00000000010000010000000100010011;
ROM[28530] <= 32'b00000001010000000000001110010011;
ROM[28531] <= 32'b00000000100000111000001110010011;
ROM[28532] <= 32'b01000000011100010000001110110011;
ROM[28533] <= 32'b00000000011100000000001000110011;
ROM[28534] <= 32'b00000000001000000000000110110011;
ROM[28535] <= 32'b01011101000100001101000011101111;
ROM[28536] <= 32'b00000110001100000000001110010011;
ROM[28537] <= 32'b00000000011100010010000000100011;
ROM[28538] <= 32'b00000000010000010000000100010011;
ROM[28539] <= 32'b00000000000000011100001110110111;
ROM[28540] <= 32'b11100011100000111000001110010011;
ROM[28541] <= 32'b00000000111000111000001110110011;
ROM[28542] <= 32'b00000000011100010010000000100011;
ROM[28543] <= 32'b00000000010000010000000100010011;
ROM[28544] <= 32'b00000000001100010010000000100011;
ROM[28545] <= 32'b00000000010000010000000100010011;
ROM[28546] <= 32'b00000000010000010010000000100011;
ROM[28547] <= 32'b00000000010000010000000100010011;
ROM[28548] <= 32'b00000000010100010010000000100011;
ROM[28549] <= 32'b00000000010000010000000100010011;
ROM[28550] <= 32'b00000000011000010010000000100011;
ROM[28551] <= 32'b00000000010000010000000100010011;
ROM[28552] <= 32'b00000001010000000000001110010011;
ROM[28553] <= 32'b00000000100000111000001110010011;
ROM[28554] <= 32'b01000000011100010000001110110011;
ROM[28555] <= 32'b00000000011100000000001000110011;
ROM[28556] <= 32'b00000000001000000000000110110011;
ROM[28557] <= 32'b01010111100100001101000011101111;
ROM[28558] <= 32'b00000110111100000000001110010011;
ROM[28559] <= 32'b00000000011100010010000000100011;
ROM[28560] <= 32'b00000000010000010000000100010011;
ROM[28561] <= 32'b00000000000000011100001110110111;
ROM[28562] <= 32'b11101001000000111000001110010011;
ROM[28563] <= 32'b00000000111000111000001110110011;
ROM[28564] <= 32'b00000000011100010010000000100011;
ROM[28565] <= 32'b00000000010000010000000100010011;
ROM[28566] <= 32'b00000000001100010010000000100011;
ROM[28567] <= 32'b00000000010000010000000100010011;
ROM[28568] <= 32'b00000000010000010010000000100011;
ROM[28569] <= 32'b00000000010000010000000100010011;
ROM[28570] <= 32'b00000000010100010010000000100011;
ROM[28571] <= 32'b00000000010000010000000100010011;
ROM[28572] <= 32'b00000000011000010010000000100011;
ROM[28573] <= 32'b00000000010000010000000100010011;
ROM[28574] <= 32'b00000001010000000000001110010011;
ROM[28575] <= 32'b00000000100000111000001110010011;
ROM[28576] <= 32'b01000000011100010000001110110011;
ROM[28577] <= 32'b00000000011100000000001000110011;
ROM[28578] <= 32'b00000000001000000000000110110011;
ROM[28579] <= 32'b01010010000100001101000011101111;
ROM[28580] <= 32'b00000110111000000000001110010011;
ROM[28581] <= 32'b00000000011100010010000000100011;
ROM[28582] <= 32'b00000000010000010000000100010011;
ROM[28583] <= 32'b00000000000000011100001110110111;
ROM[28584] <= 32'b11101110100000111000001110010011;
ROM[28585] <= 32'b00000000111000111000001110110011;
ROM[28586] <= 32'b00000000011100010010000000100011;
ROM[28587] <= 32'b00000000010000010000000100010011;
ROM[28588] <= 32'b00000000001100010010000000100011;
ROM[28589] <= 32'b00000000010000010000000100010011;
ROM[28590] <= 32'b00000000010000010010000000100011;
ROM[28591] <= 32'b00000000010000010000000100010011;
ROM[28592] <= 32'b00000000010100010010000000100011;
ROM[28593] <= 32'b00000000010000010000000100010011;
ROM[28594] <= 32'b00000000011000010010000000100011;
ROM[28595] <= 32'b00000000010000010000000100010011;
ROM[28596] <= 32'b00000001010000000000001110010011;
ROM[28597] <= 32'b00000000100000111000001110010011;
ROM[28598] <= 32'b01000000011100010000001110110011;
ROM[28599] <= 32'b00000000011100000000001000110011;
ROM[28600] <= 32'b00000000001000000000000110110011;
ROM[28601] <= 32'b01001100100100001101000011101111;
ROM[28602] <= 32'b00000111010000000000001110010011;
ROM[28603] <= 32'b00000000011100010010000000100011;
ROM[28604] <= 32'b00000000010000010000000100010011;
ROM[28605] <= 32'b00000000000000011100001110110111;
ROM[28606] <= 32'b11110100000000111000001110010011;
ROM[28607] <= 32'b00000000111000111000001110110011;
ROM[28608] <= 32'b00000000011100010010000000100011;
ROM[28609] <= 32'b00000000010000010000000100010011;
ROM[28610] <= 32'b00000000001100010010000000100011;
ROM[28611] <= 32'b00000000010000010000000100010011;
ROM[28612] <= 32'b00000000010000010010000000100011;
ROM[28613] <= 32'b00000000010000010000000100010011;
ROM[28614] <= 32'b00000000010100010010000000100011;
ROM[28615] <= 32'b00000000010000010000000100010011;
ROM[28616] <= 32'b00000000011000010010000000100011;
ROM[28617] <= 32'b00000000010000010000000100010011;
ROM[28618] <= 32'b00000001010000000000001110010011;
ROM[28619] <= 32'b00000000100000111000001110010011;
ROM[28620] <= 32'b01000000011100010000001110110011;
ROM[28621] <= 32'b00000000011100000000001000110011;
ROM[28622] <= 32'b00000000001000000000000110110011;
ROM[28623] <= 32'b01000111000100001101000011101111;
ROM[28624] <= 32'b00000110100100000000001110010011;
ROM[28625] <= 32'b00000000011100010010000000100011;
ROM[28626] <= 32'b00000000010000010000000100010011;
ROM[28627] <= 32'b00000000000000011100001110110111;
ROM[28628] <= 32'b11111001100000111000001110010011;
ROM[28629] <= 32'b00000000111000111000001110110011;
ROM[28630] <= 32'b00000000011100010010000000100011;
ROM[28631] <= 32'b00000000010000010000000100010011;
ROM[28632] <= 32'b00000000001100010010000000100011;
ROM[28633] <= 32'b00000000010000010000000100010011;
ROM[28634] <= 32'b00000000010000010010000000100011;
ROM[28635] <= 32'b00000000010000010000000100010011;
ROM[28636] <= 32'b00000000010100010010000000100011;
ROM[28637] <= 32'b00000000010000010000000100010011;
ROM[28638] <= 32'b00000000011000010010000000100011;
ROM[28639] <= 32'b00000000010000010000000100010011;
ROM[28640] <= 32'b00000001010000000000001110010011;
ROM[28641] <= 32'b00000000100000111000001110010011;
ROM[28642] <= 32'b01000000011100010000001110110011;
ROM[28643] <= 32'b00000000011100000000001000110011;
ROM[28644] <= 32'b00000000001000000000000110110011;
ROM[28645] <= 32'b01000001100100001101000011101111;
ROM[28646] <= 32'b00000110111000000000001110010011;
ROM[28647] <= 32'b00000000011100010010000000100011;
ROM[28648] <= 32'b00000000010000010000000100010011;
ROM[28649] <= 32'b00000000000000011100001110110111;
ROM[28650] <= 32'b11111111000000111000001110010011;
ROM[28651] <= 32'b00000000111000111000001110110011;
ROM[28652] <= 32'b00000000011100010010000000100011;
ROM[28653] <= 32'b00000000010000010000000100010011;
ROM[28654] <= 32'b00000000001100010010000000100011;
ROM[28655] <= 32'b00000000010000010000000100010011;
ROM[28656] <= 32'b00000000010000010010000000100011;
ROM[28657] <= 32'b00000000010000010000000100010011;
ROM[28658] <= 32'b00000000010100010010000000100011;
ROM[28659] <= 32'b00000000010000010000000100010011;
ROM[28660] <= 32'b00000000011000010010000000100011;
ROM[28661] <= 32'b00000000010000010000000100010011;
ROM[28662] <= 32'b00000001010000000000001110010011;
ROM[28663] <= 32'b00000000100000111000001110010011;
ROM[28664] <= 32'b01000000011100010000001110110011;
ROM[28665] <= 32'b00000000011100000000001000110011;
ROM[28666] <= 32'b00000000001000000000000110110011;
ROM[28667] <= 32'b00111100000100001101000011101111;
ROM[28668] <= 32'b00000111010100000000001110010011;
ROM[28669] <= 32'b00000000011100010010000000100011;
ROM[28670] <= 32'b00000000010000010000000100010011;
ROM[28671] <= 32'b00000000000000011100001110110111;
ROM[28672] <= 32'b00000100100000111000001110010011;
ROM[28673] <= 32'b00000000111000111000001110110011;
ROM[28674] <= 32'b00000000011100010010000000100011;
ROM[28675] <= 32'b00000000010000010000000100010011;
ROM[28676] <= 32'b00000000001100010010000000100011;
ROM[28677] <= 32'b00000000010000010000000100010011;
ROM[28678] <= 32'b00000000010000010010000000100011;
ROM[28679] <= 32'b00000000010000010000000100010011;
ROM[28680] <= 32'b00000000010100010010000000100011;
ROM[28681] <= 32'b00000000010000010000000100010011;
ROM[28682] <= 32'b00000000011000010010000000100011;
ROM[28683] <= 32'b00000000010000010000000100010011;
ROM[28684] <= 32'b00000001010000000000001110010011;
ROM[28685] <= 32'b00000000100000111000001110010011;
ROM[28686] <= 32'b01000000011100010000001110110011;
ROM[28687] <= 32'b00000000011100000000001000110011;
ROM[28688] <= 32'b00000000001000000000000110110011;
ROM[28689] <= 32'b00110110100100001101000011101111;
ROM[28690] <= 32'b00000110010100000000001110010011;
ROM[28691] <= 32'b00000000011100010010000000100011;
ROM[28692] <= 32'b00000000010000010000000100010011;
ROM[28693] <= 32'b00000000000000011100001110110111;
ROM[28694] <= 32'b00001010000000111000001110010011;
ROM[28695] <= 32'b00000000111000111000001110110011;
ROM[28696] <= 32'b00000000011100010010000000100011;
ROM[28697] <= 32'b00000000010000010000000100010011;
ROM[28698] <= 32'b00000000001100010010000000100011;
ROM[28699] <= 32'b00000000010000010000000100010011;
ROM[28700] <= 32'b00000000010000010010000000100011;
ROM[28701] <= 32'b00000000010000010000000100010011;
ROM[28702] <= 32'b00000000010100010010000000100011;
ROM[28703] <= 32'b00000000010000010000000100010011;
ROM[28704] <= 32'b00000000011000010010000000100011;
ROM[28705] <= 32'b00000000010000010000000100010011;
ROM[28706] <= 32'b00000001010000000000001110010011;
ROM[28707] <= 32'b00000000100000111000001110010011;
ROM[28708] <= 32'b01000000011100010000001110110011;
ROM[28709] <= 32'b00000000011100000000001000110011;
ROM[28710] <= 32'b00000000001000000000000110110011;
ROM[28711] <= 32'b00110001000100001101000011101111;
ROM[28712] <= 32'b00000011111100000000001110010011;
ROM[28713] <= 32'b00000000011100010010000000100011;
ROM[28714] <= 32'b00000000010000010000000100010011;
ROM[28715] <= 32'b00000000000000011100001110110111;
ROM[28716] <= 32'b00001111100000111000001110010011;
ROM[28717] <= 32'b00000000111000111000001110110011;
ROM[28718] <= 32'b00000000011100010010000000100011;
ROM[28719] <= 32'b00000000010000010000000100010011;
ROM[28720] <= 32'b00000000001100010010000000100011;
ROM[28721] <= 32'b00000000010000010000000100010011;
ROM[28722] <= 32'b00000000010000010010000000100011;
ROM[28723] <= 32'b00000000010000010000000100010011;
ROM[28724] <= 32'b00000000010100010010000000100011;
ROM[28725] <= 32'b00000000010000010000000100010011;
ROM[28726] <= 32'b00000000011000010010000000100011;
ROM[28727] <= 32'b00000000010000010000000100010011;
ROM[28728] <= 32'b00000001010000000000001110010011;
ROM[28729] <= 32'b00000000100000111000001110010011;
ROM[28730] <= 32'b01000000011100010000001110110011;
ROM[28731] <= 32'b00000000011100000000001000110011;
ROM[28732] <= 32'b00000000001000000000000110110011;
ROM[28733] <= 32'b00101011100100001101000011101111;
ROM[28734] <= 32'b00000010000000000000001110010011;
ROM[28735] <= 32'b00000000011100010010000000100011;
ROM[28736] <= 32'b00000000010000010000000100010011;
ROM[28737] <= 32'b00000000000000011100001110110111;
ROM[28738] <= 32'b00010101000000111000001110010011;
ROM[28739] <= 32'b00000000111000111000001110110011;
ROM[28740] <= 32'b00000000011100010010000000100011;
ROM[28741] <= 32'b00000000010000010000000100010011;
ROM[28742] <= 32'b00000000001100010010000000100011;
ROM[28743] <= 32'b00000000010000010000000100010011;
ROM[28744] <= 32'b00000000010000010010000000100011;
ROM[28745] <= 32'b00000000010000010000000100010011;
ROM[28746] <= 32'b00000000010100010010000000100011;
ROM[28747] <= 32'b00000000010000010000000100010011;
ROM[28748] <= 32'b00000000011000010010000000100011;
ROM[28749] <= 32'b00000000010000010000000100010011;
ROM[28750] <= 32'b00000001010000000000001110010011;
ROM[28751] <= 32'b00000000100000111000001110010011;
ROM[28752] <= 32'b01000000011100010000001110110011;
ROM[28753] <= 32'b00000000011100000000001000110011;
ROM[28754] <= 32'b00000000001000000000000110110011;
ROM[28755] <= 32'b00100110000100001101000011101111;
ROM[28756] <= 32'b00000010100000000000001110010011;
ROM[28757] <= 32'b00000000011100010010000000100011;
ROM[28758] <= 32'b00000000010000010000000100010011;
ROM[28759] <= 32'b00000000000000011100001110110111;
ROM[28760] <= 32'b00011010100000111000001110010011;
ROM[28761] <= 32'b00000000111000111000001110110011;
ROM[28762] <= 32'b00000000011100010010000000100011;
ROM[28763] <= 32'b00000000010000010000000100010011;
ROM[28764] <= 32'b00000000001100010010000000100011;
ROM[28765] <= 32'b00000000010000010000000100010011;
ROM[28766] <= 32'b00000000010000010010000000100011;
ROM[28767] <= 32'b00000000010000010000000100010011;
ROM[28768] <= 32'b00000000010100010010000000100011;
ROM[28769] <= 32'b00000000010000010000000100010011;
ROM[28770] <= 32'b00000000011000010010000000100011;
ROM[28771] <= 32'b00000000010000010000000100010011;
ROM[28772] <= 32'b00000001010000000000001110010011;
ROM[28773] <= 32'b00000000100000111000001110010011;
ROM[28774] <= 32'b01000000011100010000001110110011;
ROM[28775] <= 32'b00000000011100000000001000110011;
ROM[28776] <= 32'b00000000001000000000000110110011;
ROM[28777] <= 32'b00100000100100001101000011101111;
ROM[28778] <= 32'b00000111100100000000001110010011;
ROM[28779] <= 32'b00000000011100010010000000100011;
ROM[28780] <= 32'b00000000010000010000000100010011;
ROM[28781] <= 32'b00000000000000011100001110110111;
ROM[28782] <= 32'b00100000000000111000001110010011;
ROM[28783] <= 32'b00000000111000111000001110110011;
ROM[28784] <= 32'b00000000011100010010000000100011;
ROM[28785] <= 32'b00000000010000010000000100010011;
ROM[28786] <= 32'b00000000001100010010000000100011;
ROM[28787] <= 32'b00000000010000010000000100010011;
ROM[28788] <= 32'b00000000010000010010000000100011;
ROM[28789] <= 32'b00000000010000010000000100010011;
ROM[28790] <= 32'b00000000010100010010000000100011;
ROM[28791] <= 32'b00000000010000010000000100010011;
ROM[28792] <= 32'b00000000011000010010000000100011;
ROM[28793] <= 32'b00000000010000010000000100010011;
ROM[28794] <= 32'b00000001010000000000001110010011;
ROM[28795] <= 32'b00000000100000111000001110010011;
ROM[28796] <= 32'b01000000011100010000001110110011;
ROM[28797] <= 32'b00000000011100000000001000110011;
ROM[28798] <= 32'b00000000001000000000000110110011;
ROM[28799] <= 32'b00011011000100001101000011101111;
ROM[28800] <= 32'b00000110010100000000001110010011;
ROM[28801] <= 32'b00000000011100010010000000100011;
ROM[28802] <= 32'b00000000010000010000000100010011;
ROM[28803] <= 32'b00000000000000011100001110110111;
ROM[28804] <= 32'b00100101100000111000001110010011;
ROM[28805] <= 32'b00000000111000111000001110110011;
ROM[28806] <= 32'b00000000011100010010000000100011;
ROM[28807] <= 32'b00000000010000010000000100010011;
ROM[28808] <= 32'b00000000001100010010000000100011;
ROM[28809] <= 32'b00000000010000010000000100010011;
ROM[28810] <= 32'b00000000010000010010000000100011;
ROM[28811] <= 32'b00000000010000010000000100010011;
ROM[28812] <= 32'b00000000010100010010000000100011;
ROM[28813] <= 32'b00000000010000010000000100010011;
ROM[28814] <= 32'b00000000011000010010000000100011;
ROM[28815] <= 32'b00000000010000010000000100010011;
ROM[28816] <= 32'b00000001010000000000001110010011;
ROM[28817] <= 32'b00000000100000111000001110010011;
ROM[28818] <= 32'b01000000011100010000001110110011;
ROM[28819] <= 32'b00000000011100000000001000110011;
ROM[28820] <= 32'b00000000001000000000000110110011;
ROM[28821] <= 32'b00010101100100001101000011101111;
ROM[28822] <= 32'b00000111001100000000001110010011;
ROM[28823] <= 32'b00000000011100010010000000100011;
ROM[28824] <= 32'b00000000010000010000000100010011;
ROM[28825] <= 32'b00000000000000011100001110110111;
ROM[28826] <= 32'b00101011000000111000001110010011;
ROM[28827] <= 32'b00000000111000111000001110110011;
ROM[28828] <= 32'b00000000011100010010000000100011;
ROM[28829] <= 32'b00000000010000010000000100010011;
ROM[28830] <= 32'b00000000001100010010000000100011;
ROM[28831] <= 32'b00000000010000010000000100010011;
ROM[28832] <= 32'b00000000010000010010000000100011;
ROM[28833] <= 32'b00000000010000010000000100010011;
ROM[28834] <= 32'b00000000010100010010000000100011;
ROM[28835] <= 32'b00000000010000010000000100010011;
ROM[28836] <= 32'b00000000011000010010000000100011;
ROM[28837] <= 32'b00000000010000010000000100010011;
ROM[28838] <= 32'b00000001010000000000001110010011;
ROM[28839] <= 32'b00000000100000111000001110010011;
ROM[28840] <= 32'b01000000011100010000001110110011;
ROM[28841] <= 32'b00000000011100000000001000110011;
ROM[28842] <= 32'b00000000001000000000000110110011;
ROM[28843] <= 32'b00010000000100001101000011101111;
ROM[28844] <= 32'b00000010100000000000001110010011;
ROM[28845] <= 32'b00000000011100010010000000100011;
ROM[28846] <= 32'b00000000010000010000000100010011;
ROM[28847] <= 32'b00000000000000011100001110110111;
ROM[28848] <= 32'b00110000100000111000001110010011;
ROM[28849] <= 32'b00000000111000111000001110110011;
ROM[28850] <= 32'b00000000011100010010000000100011;
ROM[28851] <= 32'b00000000010000010000000100010011;
ROM[28852] <= 32'b00000000001100010010000000100011;
ROM[28853] <= 32'b00000000010000010000000100010011;
ROM[28854] <= 32'b00000000010000010010000000100011;
ROM[28855] <= 32'b00000000010000010000000100010011;
ROM[28856] <= 32'b00000000010100010010000000100011;
ROM[28857] <= 32'b00000000010000010000000100010011;
ROM[28858] <= 32'b00000000011000010010000000100011;
ROM[28859] <= 32'b00000000010000010000000100010011;
ROM[28860] <= 32'b00000001010000000000001110010011;
ROM[28861] <= 32'b00000000100000111000001110010011;
ROM[28862] <= 32'b01000000011100010000001110110011;
ROM[28863] <= 32'b00000000011100000000001000110011;
ROM[28864] <= 32'b00000000001000000000000110110011;
ROM[28865] <= 32'b00001010100100001101000011101111;
ROM[28866] <= 32'b00000011000100000000001110010011;
ROM[28867] <= 32'b00000000011100010010000000100011;
ROM[28868] <= 32'b00000000010000010000000100010011;
ROM[28869] <= 32'b00000000000000011100001110110111;
ROM[28870] <= 32'b00110110000000111000001110010011;
ROM[28871] <= 32'b00000000111000111000001110110011;
ROM[28872] <= 32'b00000000011100010010000000100011;
ROM[28873] <= 32'b00000000010000010000000100010011;
ROM[28874] <= 32'b00000000001100010010000000100011;
ROM[28875] <= 32'b00000000010000010000000100010011;
ROM[28876] <= 32'b00000000010000010010000000100011;
ROM[28877] <= 32'b00000000010000010000000100010011;
ROM[28878] <= 32'b00000000010100010010000000100011;
ROM[28879] <= 32'b00000000010000010000000100010011;
ROM[28880] <= 32'b00000000011000010010000000100011;
ROM[28881] <= 32'b00000000010000010000000100010011;
ROM[28882] <= 32'b00000001010000000000001110010011;
ROM[28883] <= 32'b00000000100000111000001110010011;
ROM[28884] <= 32'b01000000011100010000001110110011;
ROM[28885] <= 32'b00000000011100000000001000110011;
ROM[28886] <= 32'b00000000001000000000000110110011;
ROM[28887] <= 32'b00000101000100001101000011101111;
ROM[28888] <= 32'b00000010100100000000001110010011;
ROM[28889] <= 32'b00000000011100010010000000100011;
ROM[28890] <= 32'b00000000010000010000000100010011;
ROM[28891] <= 32'b00000000000000011100001110110111;
ROM[28892] <= 32'b00111011100000111000001110010011;
ROM[28893] <= 32'b00000000111000111000001110110011;
ROM[28894] <= 32'b00000000011100010010000000100011;
ROM[28895] <= 32'b00000000010000010000000100010011;
ROM[28896] <= 32'b00000000001100010010000000100011;
ROM[28897] <= 32'b00000000010000010000000100010011;
ROM[28898] <= 32'b00000000010000010010000000100011;
ROM[28899] <= 32'b00000000010000010000000100010011;
ROM[28900] <= 32'b00000000010100010010000000100011;
ROM[28901] <= 32'b00000000010000010000000100010011;
ROM[28902] <= 32'b00000000011000010010000000100011;
ROM[28903] <= 32'b00000000010000010000000100010011;
ROM[28904] <= 32'b00000001010000000000001110010011;
ROM[28905] <= 32'b00000000100000111000001110010011;
ROM[28906] <= 32'b01000000011100010000001110110011;
ROM[28907] <= 32'b00000000011100000000001000110011;
ROM[28908] <= 32'b00000000001000000000000110110011;
ROM[28909] <= 32'b01111111100000001101000011101111;
ROM[28910] <= 32'b00000010111100000000001110010011;
ROM[28911] <= 32'b00000000011100010010000000100011;
ROM[28912] <= 32'b00000000010000010000000100010011;
ROM[28913] <= 32'b00000000000000011100001110110111;
ROM[28914] <= 32'b01000001000000111000001110010011;
ROM[28915] <= 32'b00000000111000111000001110110011;
ROM[28916] <= 32'b00000000011100010010000000100011;
ROM[28917] <= 32'b00000000010000010000000100010011;
ROM[28918] <= 32'b00000000001100010010000000100011;
ROM[28919] <= 32'b00000000010000010000000100010011;
ROM[28920] <= 32'b00000000010000010010000000100011;
ROM[28921] <= 32'b00000000010000010000000100010011;
ROM[28922] <= 32'b00000000010100010010000000100011;
ROM[28923] <= 32'b00000000010000010000000100010011;
ROM[28924] <= 32'b00000000011000010010000000100011;
ROM[28925] <= 32'b00000000010000010000000100010011;
ROM[28926] <= 32'b00000001010000000000001110010011;
ROM[28927] <= 32'b00000000100000111000001110010011;
ROM[28928] <= 32'b01000000011100010000001110110011;
ROM[28929] <= 32'b00000000011100000000001000110011;
ROM[28930] <= 32'b00000000001000000000000110110011;
ROM[28931] <= 32'b01111010000000001101000011101111;
ROM[28932] <= 32'b00000110111000000000001110010011;
ROM[28933] <= 32'b00000000011100010010000000100011;
ROM[28934] <= 32'b00000000010000010000000100010011;
ROM[28935] <= 32'b00000000000000011100001110110111;
ROM[28936] <= 32'b01000110100000111000001110010011;
ROM[28937] <= 32'b00000000111000111000001110110011;
ROM[28938] <= 32'b00000000011100010010000000100011;
ROM[28939] <= 32'b00000000010000010000000100010011;
ROM[28940] <= 32'b00000000001100010010000000100011;
ROM[28941] <= 32'b00000000010000010000000100010011;
ROM[28942] <= 32'b00000000010000010010000000100011;
ROM[28943] <= 32'b00000000010000010000000100010011;
ROM[28944] <= 32'b00000000010100010010000000100011;
ROM[28945] <= 32'b00000000010000010000000100010011;
ROM[28946] <= 32'b00000000011000010010000000100011;
ROM[28947] <= 32'b00000000010000010000000100010011;
ROM[28948] <= 32'b00000001010000000000001110010011;
ROM[28949] <= 32'b00000000100000111000001110010011;
ROM[28950] <= 32'b01000000011100010000001110110011;
ROM[28951] <= 32'b00000000011100000000001000110011;
ROM[28952] <= 32'b00000000001000000000000110110011;
ROM[28953] <= 32'b01110100100000001101000011101111;
ROM[28954] <= 32'b00000110111100000000001110010011;
ROM[28955] <= 32'b00000000011100010010000000100011;
ROM[28956] <= 32'b00000000010000010000000100010011;
ROM[28957] <= 32'b00000000000000011100001110110111;
ROM[28958] <= 32'b01001100000000111000001110010011;
ROM[28959] <= 32'b00000000111000111000001110110011;
ROM[28960] <= 32'b00000000011100010010000000100011;
ROM[28961] <= 32'b00000000010000010000000100010011;
ROM[28962] <= 32'b00000000001100010010000000100011;
ROM[28963] <= 32'b00000000010000010000000100010011;
ROM[28964] <= 32'b00000000010000010010000000100011;
ROM[28965] <= 32'b00000000010000010000000100010011;
ROM[28966] <= 32'b00000000010100010010000000100011;
ROM[28967] <= 32'b00000000010000010000000100010011;
ROM[28968] <= 32'b00000000011000010010000000100011;
ROM[28969] <= 32'b00000000010000010000000100010011;
ROM[28970] <= 32'b00000001010000000000001110010011;
ROM[28971] <= 32'b00000000100000111000001110010011;
ROM[28972] <= 32'b01000000011100010000001110110011;
ROM[28973] <= 32'b00000000011100000000001000110011;
ROM[28974] <= 32'b00000000001000000000000110110011;
ROM[28975] <= 32'b01101111000000001101000011101111;
ROM[28976] <= 32'b00000010100000000000001110010011;
ROM[28977] <= 32'b00000000011100010010000000100011;
ROM[28978] <= 32'b00000000010000010000000100010011;
ROM[28979] <= 32'b00000000000000011100001110110111;
ROM[28980] <= 32'b01010001100000111000001110010011;
ROM[28981] <= 32'b00000000111000111000001110110011;
ROM[28982] <= 32'b00000000011100010010000000100011;
ROM[28983] <= 32'b00000000010000010000000100010011;
ROM[28984] <= 32'b00000000001100010010000000100011;
ROM[28985] <= 32'b00000000010000010000000100010011;
ROM[28986] <= 32'b00000000010000010010000000100011;
ROM[28987] <= 32'b00000000010000010000000100010011;
ROM[28988] <= 32'b00000000010100010010000000100011;
ROM[28989] <= 32'b00000000010000010000000100010011;
ROM[28990] <= 32'b00000000011000010010000000100011;
ROM[28991] <= 32'b00000000010000010000000100010011;
ROM[28992] <= 32'b00000001010000000000001110010011;
ROM[28993] <= 32'b00000000100000111000001110010011;
ROM[28994] <= 32'b01000000011100010000001110110011;
ROM[28995] <= 32'b00000000011100000000001000110011;
ROM[28996] <= 32'b00000000001000000000000110110011;
ROM[28997] <= 32'b01101001100000001101000011101111;
ROM[28998] <= 32'b00000011000000000000001110010011;
ROM[28999] <= 32'b00000000011100010010000000100011;
ROM[29000] <= 32'b00000000010000010000000100010011;
ROM[29001] <= 32'b00000000000000011100001110110111;
ROM[29002] <= 32'b01010111000000111000001110010011;
ROM[29003] <= 32'b00000000111000111000001110110011;
ROM[29004] <= 32'b00000000011100010010000000100011;
ROM[29005] <= 32'b00000000010000010000000100010011;
ROM[29006] <= 32'b00000000001100010010000000100011;
ROM[29007] <= 32'b00000000010000010000000100010011;
ROM[29008] <= 32'b00000000010000010010000000100011;
ROM[29009] <= 32'b00000000010000010000000100010011;
ROM[29010] <= 32'b00000000010100010010000000100011;
ROM[29011] <= 32'b00000000010000010000000100010011;
ROM[29012] <= 32'b00000000011000010010000000100011;
ROM[29013] <= 32'b00000000010000010000000100010011;
ROM[29014] <= 32'b00000001010000000000001110010011;
ROM[29015] <= 32'b00000000100000111000001110010011;
ROM[29016] <= 32'b01000000011100010000001110110011;
ROM[29017] <= 32'b00000000011100000000001000110011;
ROM[29018] <= 32'b00000000001000000000000110110011;
ROM[29019] <= 32'b01100100000000001101000011101111;
ROM[29020] <= 32'b00000010100100000000001110010011;
ROM[29021] <= 32'b00000000011100010010000000100011;
ROM[29022] <= 32'b00000000010000010000000100010011;
ROM[29023] <= 32'b00000000000000011100001110110111;
ROM[29024] <= 32'b01011100100000111000001110010011;
ROM[29025] <= 32'b00000000111000111000001110110011;
ROM[29026] <= 32'b00000000011100010010000000100011;
ROM[29027] <= 32'b00000000010000010000000100010011;
ROM[29028] <= 32'b00000000001100010010000000100011;
ROM[29029] <= 32'b00000000010000010000000100010011;
ROM[29030] <= 32'b00000000010000010010000000100011;
ROM[29031] <= 32'b00000000010000010000000100010011;
ROM[29032] <= 32'b00000000010100010010000000100011;
ROM[29033] <= 32'b00000000010000010000000100010011;
ROM[29034] <= 32'b00000000011000010010000000100011;
ROM[29035] <= 32'b00000000010000010000000100010011;
ROM[29036] <= 32'b00000001010000000000001110010011;
ROM[29037] <= 32'b00000000100000111000001110010011;
ROM[29038] <= 32'b01000000011100010000001110110011;
ROM[29039] <= 32'b00000000011100000000001000110011;
ROM[29040] <= 32'b00000000001000000000000110110011;
ROM[29041] <= 32'b01011110100000001101000011101111;
ROM[29042] <= 32'b00000010100100000000001110010011;
ROM[29043] <= 32'b00000000011100010010000000100011;
ROM[29044] <= 32'b00000000010000010000000100010011;
ROM[29045] <= 32'b00000000000000011100001110110111;
ROM[29046] <= 32'b01100010000000111000001110010011;
ROM[29047] <= 32'b00000000111000111000001110110011;
ROM[29048] <= 32'b00000000011100010010000000100011;
ROM[29049] <= 32'b00000000010000010000000100010011;
ROM[29050] <= 32'b00000000001100010010000000100011;
ROM[29051] <= 32'b00000000010000010000000100010011;
ROM[29052] <= 32'b00000000010000010010000000100011;
ROM[29053] <= 32'b00000000010000010000000100010011;
ROM[29054] <= 32'b00000000010100010010000000100011;
ROM[29055] <= 32'b00000000010000010000000100010011;
ROM[29056] <= 32'b00000000011000010010000000100011;
ROM[29057] <= 32'b00000000010000010000000100010011;
ROM[29058] <= 32'b00000001010000000000001110010011;
ROM[29059] <= 32'b00000000100000111000001110010011;
ROM[29060] <= 32'b01000000011100010000001110110011;
ROM[29061] <= 32'b00000000011100000000001000110011;
ROM[29062] <= 32'b00000000001000000000000110110011;
ROM[29063] <= 32'b01011001000000001101000011101111;
ROM[29064] <= 32'b00000011101000000000001110010011;
ROM[29065] <= 32'b00000000011100010010000000100011;
ROM[29066] <= 32'b00000000010000010000000100010011;
ROM[29067] <= 32'b00000000000000011100001110110111;
ROM[29068] <= 32'b01100111100000111000001110010011;
ROM[29069] <= 32'b00000000111000111000001110110011;
ROM[29070] <= 32'b00000000011100010010000000100011;
ROM[29071] <= 32'b00000000010000010000000100010011;
ROM[29072] <= 32'b00000000001100010010000000100011;
ROM[29073] <= 32'b00000000010000010000000100010011;
ROM[29074] <= 32'b00000000010000010010000000100011;
ROM[29075] <= 32'b00000000010000010000000100010011;
ROM[29076] <= 32'b00000000010100010010000000100011;
ROM[29077] <= 32'b00000000010000010000000100010011;
ROM[29078] <= 32'b00000000011000010010000000100011;
ROM[29079] <= 32'b00000000010000010000000100010011;
ROM[29080] <= 32'b00000001010000000000001110010011;
ROM[29081] <= 32'b00000000100000111000001110010011;
ROM[29082] <= 32'b01000000011100010000001110110011;
ROM[29083] <= 32'b00000000011100000000001000110011;
ROM[29084] <= 32'b00000000001000000000000110110011;
ROM[29085] <= 32'b01010011100000001101000011101111;
ROM[29086] <= 32'b00000010000000000000001110010011;
ROM[29087] <= 32'b00000000011100010010000000100011;
ROM[29088] <= 32'b00000000010000010000000100010011;
ROM[29089] <= 32'b00000000000000011100001110110111;
ROM[29090] <= 32'b01101101000000111000001110010011;
ROM[29091] <= 32'b00000000111000111000001110110011;
ROM[29092] <= 32'b00000000011100010010000000100011;
ROM[29093] <= 32'b00000000010000010000000100010011;
ROM[29094] <= 32'b00000000001100010010000000100011;
ROM[29095] <= 32'b00000000010000010000000100010011;
ROM[29096] <= 32'b00000000010000010010000000100011;
ROM[29097] <= 32'b00000000010000010000000100010011;
ROM[29098] <= 32'b00000000010100010010000000100011;
ROM[29099] <= 32'b00000000010000010000000100010011;
ROM[29100] <= 32'b00000000011000010010000000100011;
ROM[29101] <= 32'b00000000010000010000000100010011;
ROM[29102] <= 32'b00000001010000000000001110010011;
ROM[29103] <= 32'b00000000100000111000001110010011;
ROM[29104] <= 32'b01000000011100010000001110110011;
ROM[29105] <= 32'b00000000011100000000001000110011;
ROM[29106] <= 32'b00000000001000000000000110110011;
ROM[29107] <= 32'b01001110000000001101000011101111;
ROM[29108] <= 32'b00000000000000011100001110110111;
ROM[29109] <= 32'b01110001110000111000001110010011;
ROM[29110] <= 32'b00000000111000111000001110110011;
ROM[29111] <= 32'b00000000011100010010000000100011;
ROM[29112] <= 32'b00000000010000010000000100010011;
ROM[29113] <= 32'b00000000001100010010000000100011;
ROM[29114] <= 32'b00000000010000010000000100010011;
ROM[29115] <= 32'b00000000010000010010000000100011;
ROM[29116] <= 32'b00000000010000010000000100010011;
ROM[29117] <= 32'b00000000010100010010000000100011;
ROM[29118] <= 32'b00000000010000010000000100010011;
ROM[29119] <= 32'b00000000011000010010000000100011;
ROM[29120] <= 32'b00000000010000010000000100010011;
ROM[29121] <= 32'b00000001010000000000001110010011;
ROM[29122] <= 32'b00000000010000111000001110010011;
ROM[29123] <= 32'b01000000011100010000001110110011;
ROM[29124] <= 32'b00000000011100000000001000110011;
ROM[29125] <= 32'b00000000001000000000000110110011;
ROM[29126] <= 32'b10011011000111110001000011101111;
ROM[29127] <= 32'b11111111110000010000000100010011;
ROM[29128] <= 32'b00000000000000010010001110000011;
ROM[29129] <= 32'b00000000011100011010001000100011;
ROM[29130] <= 32'b00000000010000011010001110000011;
ROM[29131] <= 32'b00000000011100010010000000100011;
ROM[29132] <= 32'b00000000010000010000000100010011;
ROM[29133] <= 32'b00000000000100000000001110010011;
ROM[29134] <= 32'b00000000011100010010000000100011;
ROM[29135] <= 32'b00000000010000010000000100010011;
ROM[29136] <= 32'b11111111110000010000000100010011;
ROM[29137] <= 32'b00000000000000010010001110000011;
ROM[29138] <= 32'b11111111110000010000000100010011;
ROM[29139] <= 32'b00000000000000010010010000000011;
ROM[29140] <= 32'b00000000011101000010010010110011;
ROM[29141] <= 32'b00000000100000111010010100110011;
ROM[29142] <= 32'b00000000101001001000001110110011;
ROM[29143] <= 32'b00000000000100111000001110010011;
ROM[29144] <= 32'b00000000000100111111001110010011;
ROM[29145] <= 32'b00000000011100010010000000100011;
ROM[29146] <= 32'b00000000010000010000000100010011;
ROM[29147] <= 32'b11111111110000010000000100010011;
ROM[29148] <= 32'b00000000000000010010001110000011;
ROM[29149] <= 32'b00000000000000111000101001100011;
ROM[29150] <= 32'b00000000000000011101001110110111;
ROM[29151] <= 32'b11010010010000111000001110010011;
ROM[29152] <= 32'b00000000111000111000001110110011;
ROM[29153] <= 32'b00000000000000111000000011100111;
ROM[29154] <= 32'b00000000000000000000001110010011;
ROM[29155] <= 32'b00000000011100010010000000100011;
ROM[29156] <= 32'b00000000010000010000000100010011;
ROM[29157] <= 32'b11111111110000010000000100010011;
ROM[29158] <= 32'b00000000000000010010001110000011;
ROM[29159] <= 32'b00000000011100011010000000100011;
ROM[29160] <= 32'b00000000111000000000001110010011;
ROM[29161] <= 32'b00000000011100010010000000100011;
ROM[29162] <= 32'b00000000010000010000000100010011;
ROM[29163] <= 32'b00000000000000011100001110110111;
ROM[29164] <= 32'b01111111100000111000001110010011;
ROM[29165] <= 32'b00000000111000111000001110110011;
ROM[29166] <= 32'b00000000011100010010000000100011;
ROM[29167] <= 32'b00000000010000010000000100010011;
ROM[29168] <= 32'b00000000001100010010000000100011;
ROM[29169] <= 32'b00000000010000010000000100010011;
ROM[29170] <= 32'b00000000010000010010000000100011;
ROM[29171] <= 32'b00000000010000010000000100010011;
ROM[29172] <= 32'b00000000010100010010000000100011;
ROM[29173] <= 32'b00000000010000010000000100010011;
ROM[29174] <= 32'b00000000011000010010000000100011;
ROM[29175] <= 32'b00000000010000010000000100010011;
ROM[29176] <= 32'b00000001010000000000001110010011;
ROM[29177] <= 32'b00000000010000111000001110010011;
ROM[29178] <= 32'b01000000011100010000001110110011;
ROM[29179] <= 32'b00000000011100000000001000110011;
ROM[29180] <= 32'b00000000001000000000000110110011;
ROM[29181] <= 32'b01110100100100001100000011101111;
ROM[29182] <= 32'b00000101000000000000001110010011;
ROM[29183] <= 32'b00000000011100010010000000100011;
ROM[29184] <= 32'b00000000010000010000000100010011;
ROM[29185] <= 32'b00000000000000011101001110110111;
ROM[29186] <= 32'b10000101000000111000001110010011;
ROM[29187] <= 32'b00000000111000111000001110110011;
ROM[29188] <= 32'b00000000011100010010000000100011;
ROM[29189] <= 32'b00000000010000010000000100010011;
ROM[29190] <= 32'b00000000001100010010000000100011;
ROM[29191] <= 32'b00000000010000010000000100010011;
ROM[29192] <= 32'b00000000010000010010000000100011;
ROM[29193] <= 32'b00000000010000010000000100010011;
ROM[29194] <= 32'b00000000010100010010000000100011;
ROM[29195] <= 32'b00000000010000010000000100010011;
ROM[29196] <= 32'b00000000011000010010000000100011;
ROM[29197] <= 32'b00000000010000010000000100010011;
ROM[29198] <= 32'b00000001010000000000001110010011;
ROM[29199] <= 32'b00000000100000111000001110010011;
ROM[29200] <= 32'b01000000011100010000001110110011;
ROM[29201] <= 32'b00000000011100000000001000110011;
ROM[29202] <= 32'b00000000001000000000000110110011;
ROM[29203] <= 32'b00110110000000001101000011101111;
ROM[29204] <= 32'b00000111001000000000001110010011;
ROM[29205] <= 32'b00000000011100010010000000100011;
ROM[29206] <= 32'b00000000010000010000000100010011;
ROM[29207] <= 32'b00000000000000011101001110110111;
ROM[29208] <= 32'b10001010100000111000001110010011;
ROM[29209] <= 32'b00000000111000111000001110110011;
ROM[29210] <= 32'b00000000011100010010000000100011;
ROM[29211] <= 32'b00000000010000010000000100010011;
ROM[29212] <= 32'b00000000001100010010000000100011;
ROM[29213] <= 32'b00000000010000010000000100010011;
ROM[29214] <= 32'b00000000010000010010000000100011;
ROM[29215] <= 32'b00000000010000010000000100010011;
ROM[29216] <= 32'b00000000010100010010000000100011;
ROM[29217] <= 32'b00000000010000010000000100010011;
ROM[29218] <= 32'b00000000011000010010000000100011;
ROM[29219] <= 32'b00000000010000010000000100010011;
ROM[29220] <= 32'b00000001010000000000001110010011;
ROM[29221] <= 32'b00000000100000111000001110010011;
ROM[29222] <= 32'b01000000011100010000001110110011;
ROM[29223] <= 32'b00000000011100000000001000110011;
ROM[29224] <= 32'b00000000001000000000000110110011;
ROM[29225] <= 32'b00110000100000001101000011101111;
ROM[29226] <= 32'b00000110111100000000001110010011;
ROM[29227] <= 32'b00000000011100010010000000100011;
ROM[29228] <= 32'b00000000010000010000000100010011;
ROM[29229] <= 32'b00000000000000011101001110110111;
ROM[29230] <= 32'b10010000000000111000001110010011;
ROM[29231] <= 32'b00000000111000111000001110110011;
ROM[29232] <= 32'b00000000011100010010000000100011;
ROM[29233] <= 32'b00000000010000010000000100010011;
ROM[29234] <= 32'b00000000001100010010000000100011;
ROM[29235] <= 32'b00000000010000010000000100010011;
ROM[29236] <= 32'b00000000010000010010000000100011;
ROM[29237] <= 32'b00000000010000010000000100010011;
ROM[29238] <= 32'b00000000010100010010000000100011;
ROM[29239] <= 32'b00000000010000010000000100010011;
ROM[29240] <= 32'b00000000011000010010000000100011;
ROM[29241] <= 32'b00000000010000010000000100010011;
ROM[29242] <= 32'b00000001010000000000001110010011;
ROM[29243] <= 32'b00000000100000111000001110010011;
ROM[29244] <= 32'b01000000011100010000001110110011;
ROM[29245] <= 32'b00000000011100000000001000110011;
ROM[29246] <= 32'b00000000001000000000000110110011;
ROM[29247] <= 32'b00101011000000001101000011101111;
ROM[29248] <= 32'b00000110011100000000001110010011;
ROM[29249] <= 32'b00000000011100010010000000100011;
ROM[29250] <= 32'b00000000010000010000000100010011;
ROM[29251] <= 32'b00000000000000011101001110110111;
ROM[29252] <= 32'b10010101100000111000001110010011;
ROM[29253] <= 32'b00000000111000111000001110110011;
ROM[29254] <= 32'b00000000011100010010000000100011;
ROM[29255] <= 32'b00000000010000010000000100010011;
ROM[29256] <= 32'b00000000001100010010000000100011;
ROM[29257] <= 32'b00000000010000010000000100010011;
ROM[29258] <= 32'b00000000010000010010000000100011;
ROM[29259] <= 32'b00000000010000010000000100010011;
ROM[29260] <= 32'b00000000010100010010000000100011;
ROM[29261] <= 32'b00000000010000010000000100010011;
ROM[29262] <= 32'b00000000011000010010000000100011;
ROM[29263] <= 32'b00000000010000010000000100010011;
ROM[29264] <= 32'b00000001010000000000001110010011;
ROM[29265] <= 32'b00000000100000111000001110010011;
ROM[29266] <= 32'b01000000011100010000001110110011;
ROM[29267] <= 32'b00000000011100000000001000110011;
ROM[29268] <= 32'b00000000001000000000000110110011;
ROM[29269] <= 32'b00100101100000001101000011101111;
ROM[29270] <= 32'b00000111001000000000001110010011;
ROM[29271] <= 32'b00000000011100010010000000100011;
ROM[29272] <= 32'b00000000010000010000000100010011;
ROM[29273] <= 32'b00000000000000011101001110110111;
ROM[29274] <= 32'b10011011000000111000001110010011;
ROM[29275] <= 32'b00000000111000111000001110110011;
ROM[29276] <= 32'b00000000011100010010000000100011;
ROM[29277] <= 32'b00000000010000010000000100010011;
ROM[29278] <= 32'b00000000001100010010000000100011;
ROM[29279] <= 32'b00000000010000010000000100010011;
ROM[29280] <= 32'b00000000010000010010000000100011;
ROM[29281] <= 32'b00000000010000010000000100010011;
ROM[29282] <= 32'b00000000010100010010000000100011;
ROM[29283] <= 32'b00000000010000010000000100010011;
ROM[29284] <= 32'b00000000011000010010000000100011;
ROM[29285] <= 32'b00000000010000010000000100010011;
ROM[29286] <= 32'b00000001010000000000001110010011;
ROM[29287] <= 32'b00000000100000111000001110010011;
ROM[29288] <= 32'b01000000011100010000001110110011;
ROM[29289] <= 32'b00000000011100000000001000110011;
ROM[29290] <= 32'b00000000001000000000000110110011;
ROM[29291] <= 32'b00100000000000001101000011101111;
ROM[29292] <= 32'b00000110000100000000001110010011;
ROM[29293] <= 32'b00000000011100010010000000100011;
ROM[29294] <= 32'b00000000010000010000000100010011;
ROM[29295] <= 32'b00000000000000011101001110110111;
ROM[29296] <= 32'b10100000100000111000001110010011;
ROM[29297] <= 32'b00000000111000111000001110110011;
ROM[29298] <= 32'b00000000011100010010000000100011;
ROM[29299] <= 32'b00000000010000010000000100010011;
ROM[29300] <= 32'b00000000001100010010000000100011;
ROM[29301] <= 32'b00000000010000010000000100010011;
ROM[29302] <= 32'b00000000010000010010000000100011;
ROM[29303] <= 32'b00000000010000010000000100010011;
ROM[29304] <= 32'b00000000010100010010000000100011;
ROM[29305] <= 32'b00000000010000010000000100010011;
ROM[29306] <= 32'b00000000011000010010000000100011;
ROM[29307] <= 32'b00000000010000010000000100010011;
ROM[29308] <= 32'b00000001010000000000001110010011;
ROM[29309] <= 32'b00000000100000111000001110010011;
ROM[29310] <= 32'b01000000011100010000001110110011;
ROM[29311] <= 32'b00000000011100000000001000110011;
ROM[29312] <= 32'b00000000001000000000000110110011;
ROM[29313] <= 32'b00011010100000001101000011101111;
ROM[29314] <= 32'b00000110110100000000001110010011;
ROM[29315] <= 32'b00000000011100010010000000100011;
ROM[29316] <= 32'b00000000010000010000000100010011;
ROM[29317] <= 32'b00000000000000011101001110110111;
ROM[29318] <= 32'b10100110000000111000001110010011;
ROM[29319] <= 32'b00000000111000111000001110110011;
ROM[29320] <= 32'b00000000011100010010000000100011;
ROM[29321] <= 32'b00000000010000010000000100010011;
ROM[29322] <= 32'b00000000001100010010000000100011;
ROM[29323] <= 32'b00000000010000010000000100010011;
ROM[29324] <= 32'b00000000010000010010000000100011;
ROM[29325] <= 32'b00000000010000010000000100010011;
ROM[29326] <= 32'b00000000010100010010000000100011;
ROM[29327] <= 32'b00000000010000010000000100010011;
ROM[29328] <= 32'b00000000011000010010000000100011;
ROM[29329] <= 32'b00000000010000010000000100010011;
ROM[29330] <= 32'b00000001010000000000001110010011;
ROM[29331] <= 32'b00000000100000111000001110010011;
ROM[29332] <= 32'b01000000011100010000001110110011;
ROM[29333] <= 32'b00000000011100000000001000110011;
ROM[29334] <= 32'b00000000001000000000000110110011;
ROM[29335] <= 32'b00010101000000001101000011101111;
ROM[29336] <= 32'b00000010000000000000001110010011;
ROM[29337] <= 32'b00000000011100010010000000100011;
ROM[29338] <= 32'b00000000010000010000000100010011;
ROM[29339] <= 32'b00000000000000011101001110110111;
ROM[29340] <= 32'b10101011100000111000001110010011;
ROM[29341] <= 32'b00000000111000111000001110110011;
ROM[29342] <= 32'b00000000011100010010000000100011;
ROM[29343] <= 32'b00000000010000010000000100010011;
ROM[29344] <= 32'b00000000001100010010000000100011;
ROM[29345] <= 32'b00000000010000010000000100010011;
ROM[29346] <= 32'b00000000010000010010000000100011;
ROM[29347] <= 32'b00000000010000010000000100010011;
ROM[29348] <= 32'b00000000010100010010000000100011;
ROM[29349] <= 32'b00000000010000010000000100010011;
ROM[29350] <= 32'b00000000011000010010000000100011;
ROM[29351] <= 32'b00000000010000010000000100010011;
ROM[29352] <= 32'b00000001010000000000001110010011;
ROM[29353] <= 32'b00000000100000111000001110010011;
ROM[29354] <= 32'b01000000011100010000001110110011;
ROM[29355] <= 32'b00000000011100000000001000110011;
ROM[29356] <= 32'b00000000001000000000000110110011;
ROM[29357] <= 32'b00001111100000001101000011101111;
ROM[29358] <= 32'b00000110010100000000001110010011;
ROM[29359] <= 32'b00000000011100010010000000100011;
ROM[29360] <= 32'b00000000010000010000000100010011;
ROM[29361] <= 32'b00000000000000011101001110110111;
ROM[29362] <= 32'b10110001000000111000001110010011;
ROM[29363] <= 32'b00000000111000111000001110110011;
ROM[29364] <= 32'b00000000011100010010000000100011;
ROM[29365] <= 32'b00000000010000010000000100010011;
ROM[29366] <= 32'b00000000001100010010000000100011;
ROM[29367] <= 32'b00000000010000010000000100010011;
ROM[29368] <= 32'b00000000010000010010000000100011;
ROM[29369] <= 32'b00000000010000010000000100010011;
ROM[29370] <= 32'b00000000010100010010000000100011;
ROM[29371] <= 32'b00000000010000010000000100010011;
ROM[29372] <= 32'b00000000011000010010000000100011;
ROM[29373] <= 32'b00000000010000010000000100010011;
ROM[29374] <= 32'b00000001010000000000001110010011;
ROM[29375] <= 32'b00000000100000111000001110010011;
ROM[29376] <= 32'b01000000011100010000001110110011;
ROM[29377] <= 32'b00000000011100000000001000110011;
ROM[29378] <= 32'b00000000001000000000000110110011;
ROM[29379] <= 32'b00001010000000001101000011101111;
ROM[29380] <= 32'b00000110111000000000001110010011;
ROM[29381] <= 32'b00000000011100010010000000100011;
ROM[29382] <= 32'b00000000010000010000000100010011;
ROM[29383] <= 32'b00000000000000011101001110110111;
ROM[29384] <= 32'b10110110100000111000001110010011;
ROM[29385] <= 32'b00000000111000111000001110110011;
ROM[29386] <= 32'b00000000011100010010000000100011;
ROM[29387] <= 32'b00000000010000010000000100010011;
ROM[29388] <= 32'b00000000001100010010000000100011;
ROM[29389] <= 32'b00000000010000010000000100010011;
ROM[29390] <= 32'b00000000010000010010000000100011;
ROM[29391] <= 32'b00000000010000010000000100010011;
ROM[29392] <= 32'b00000000010100010010000000100011;
ROM[29393] <= 32'b00000000010000010000000100010011;
ROM[29394] <= 32'b00000000011000010010000000100011;
ROM[29395] <= 32'b00000000010000010000000100010011;
ROM[29396] <= 32'b00000001010000000000001110010011;
ROM[29397] <= 32'b00000000100000111000001110010011;
ROM[29398] <= 32'b01000000011100010000001110110011;
ROM[29399] <= 32'b00000000011100000000001000110011;
ROM[29400] <= 32'b00000000001000000000000110110011;
ROM[29401] <= 32'b00000100100000001101000011101111;
ROM[29402] <= 32'b00000110010000000000001110010011;
ROM[29403] <= 32'b00000000011100010010000000100011;
ROM[29404] <= 32'b00000000010000010000000100010011;
ROM[29405] <= 32'b00000000000000011101001110110111;
ROM[29406] <= 32'b10111100000000111000001110010011;
ROM[29407] <= 32'b00000000111000111000001110110011;
ROM[29408] <= 32'b00000000011100010010000000100011;
ROM[29409] <= 32'b00000000010000010000000100010011;
ROM[29410] <= 32'b00000000001100010010000000100011;
ROM[29411] <= 32'b00000000010000010000000100010011;
ROM[29412] <= 32'b00000000010000010010000000100011;
ROM[29413] <= 32'b00000000010000010000000100010011;
ROM[29414] <= 32'b00000000010100010010000000100011;
ROM[29415] <= 32'b00000000010000010000000100010011;
ROM[29416] <= 32'b00000000011000010010000000100011;
ROM[29417] <= 32'b00000000010000010000000100010011;
ROM[29418] <= 32'b00000001010000000000001110010011;
ROM[29419] <= 32'b00000000100000111000001110010011;
ROM[29420] <= 32'b01000000011100010000001110110011;
ROM[29421] <= 32'b00000000011100000000001000110011;
ROM[29422] <= 32'b00000000001000000000000110110011;
ROM[29423] <= 32'b01111111000100001100000011101111;
ROM[29424] <= 32'b00000110010100000000001110010011;
ROM[29425] <= 32'b00000000011100010010000000100011;
ROM[29426] <= 32'b00000000010000010000000100010011;
ROM[29427] <= 32'b00000000000000011101001110110111;
ROM[29428] <= 32'b11000001100000111000001110010011;
ROM[29429] <= 32'b00000000111000111000001110110011;
ROM[29430] <= 32'b00000000011100010010000000100011;
ROM[29431] <= 32'b00000000010000010000000100010011;
ROM[29432] <= 32'b00000000001100010010000000100011;
ROM[29433] <= 32'b00000000010000010000000100010011;
ROM[29434] <= 32'b00000000010000010010000000100011;
ROM[29435] <= 32'b00000000010000010000000100010011;
ROM[29436] <= 32'b00000000010100010010000000100011;
ROM[29437] <= 32'b00000000010000010000000100010011;
ROM[29438] <= 32'b00000000011000010010000000100011;
ROM[29439] <= 32'b00000000010000010000000100010011;
ROM[29440] <= 32'b00000001010000000000001110010011;
ROM[29441] <= 32'b00000000100000111000001110010011;
ROM[29442] <= 32'b01000000011100010000001110110011;
ROM[29443] <= 32'b00000000011100000000001000110011;
ROM[29444] <= 32'b00000000001000000000000110110011;
ROM[29445] <= 32'b01111001100100001100000011101111;
ROM[29446] <= 32'b00000110010000000000001110010011;
ROM[29447] <= 32'b00000000011100010010000000100011;
ROM[29448] <= 32'b00000000010000010000000100010011;
ROM[29449] <= 32'b00000000000000011101001110110111;
ROM[29450] <= 32'b11000111000000111000001110010011;
ROM[29451] <= 32'b00000000111000111000001110110011;
ROM[29452] <= 32'b00000000011100010010000000100011;
ROM[29453] <= 32'b00000000010000010000000100010011;
ROM[29454] <= 32'b00000000001100010010000000100011;
ROM[29455] <= 32'b00000000010000010000000100010011;
ROM[29456] <= 32'b00000000010000010010000000100011;
ROM[29457] <= 32'b00000000010000010000000100010011;
ROM[29458] <= 32'b00000000010100010010000000100011;
ROM[29459] <= 32'b00000000010000010000000100010011;
ROM[29460] <= 32'b00000000011000010010000000100011;
ROM[29461] <= 32'b00000000010000010000000100010011;
ROM[29462] <= 32'b00000001010000000000001110010011;
ROM[29463] <= 32'b00000000100000111000001110010011;
ROM[29464] <= 32'b01000000011100010000001110110011;
ROM[29465] <= 32'b00000000011100000000001000110011;
ROM[29466] <= 32'b00000000001000000000000110110011;
ROM[29467] <= 32'b01110100000100001100000011101111;
ROM[29468] <= 32'b00000010111000000000001110010011;
ROM[29469] <= 32'b00000000011100010010000000100011;
ROM[29470] <= 32'b00000000010000010000000100010011;
ROM[29471] <= 32'b00000000000000011101001110110111;
ROM[29472] <= 32'b11001100100000111000001110010011;
ROM[29473] <= 32'b00000000111000111000001110110011;
ROM[29474] <= 32'b00000000011100010010000000100011;
ROM[29475] <= 32'b00000000010000010000000100010011;
ROM[29476] <= 32'b00000000001100010010000000100011;
ROM[29477] <= 32'b00000000010000010000000100010011;
ROM[29478] <= 32'b00000000010000010010000000100011;
ROM[29479] <= 32'b00000000010000010000000100010011;
ROM[29480] <= 32'b00000000010100010010000000100011;
ROM[29481] <= 32'b00000000010000010000000100010011;
ROM[29482] <= 32'b00000000011000010010000000100011;
ROM[29483] <= 32'b00000000010000010000000100010011;
ROM[29484] <= 32'b00000001010000000000001110010011;
ROM[29485] <= 32'b00000000100000111000001110010011;
ROM[29486] <= 32'b01000000011100010000001110110011;
ROM[29487] <= 32'b00000000011100000000001000110011;
ROM[29488] <= 32'b00000000001000000000000110110011;
ROM[29489] <= 32'b01101110100100001100000011101111;
ROM[29490] <= 32'b00000000000000011101001110110111;
ROM[29491] <= 32'b11010001010000111000001110010011;
ROM[29492] <= 32'b00000000111000111000001110110011;
ROM[29493] <= 32'b00000000011100010010000000100011;
ROM[29494] <= 32'b00000000010000010000000100010011;
ROM[29495] <= 32'b00000000001100010010000000100011;
ROM[29496] <= 32'b00000000010000010000000100010011;
ROM[29497] <= 32'b00000000010000010010000000100011;
ROM[29498] <= 32'b00000000010000010000000100010011;
ROM[29499] <= 32'b00000000010100010010000000100011;
ROM[29500] <= 32'b00000000010000010000000100010011;
ROM[29501] <= 32'b00000000011000010010000000100011;
ROM[29502] <= 32'b00000000010000010000000100010011;
ROM[29503] <= 32'b00000001010000000000001110010011;
ROM[29504] <= 32'b00000000010000111000001110010011;
ROM[29505] <= 32'b01000000011100010000001110110011;
ROM[29506] <= 32'b00000000011100000000001000110011;
ROM[29507] <= 32'b00000000001000000000000110110011;
ROM[29508] <= 32'b10100101100011111010000011101111;
ROM[29509] <= 32'b11111111110000010000000100010011;
ROM[29510] <= 32'b00000000000000010010001110000011;
ROM[29511] <= 32'b00000000011101100010000000100011;
ROM[29512] <= 32'b00000101110000000000000011101111;
ROM[29513] <= 32'b00000000000000011101001110110111;
ROM[29514] <= 32'b11010111000000111000001110010011;
ROM[29515] <= 32'b00000000111000111000001110110011;
ROM[29516] <= 32'b00000000011100010010000000100011;
ROM[29517] <= 32'b00000000010000010000000100010011;
ROM[29518] <= 32'b00000000001100010010000000100011;
ROM[29519] <= 32'b00000000010000010000000100010011;
ROM[29520] <= 32'b00000000010000010010000000100011;
ROM[29521] <= 32'b00000000010000010000000100010011;
ROM[29522] <= 32'b00000000010100010010000000100011;
ROM[29523] <= 32'b00000000010000010000000100010011;
ROM[29524] <= 32'b00000000011000010010000000100011;
ROM[29525] <= 32'b00000000010000010000000100010011;
ROM[29526] <= 32'b00000001010000000000001110010011;
ROM[29527] <= 32'b00000000000000111000001110010011;
ROM[29528] <= 32'b01000000011100010000001110110011;
ROM[29529] <= 32'b00000000011100000000001000110011;
ROM[29530] <= 32'b00000000001000000000000110110011;
ROM[29531] <= 32'b11101101000011111011000011101111;
ROM[29532] <= 32'b11111111110000010000000100010011;
ROM[29533] <= 32'b00000000000000010010001110000011;
ROM[29534] <= 32'b00000000011101100010000000100011;
ROM[29535] <= 32'b10100001010111111110000011101111;
ROM[29536] <= 32'b00000000000000000000001110010011;
ROM[29537] <= 32'b00000000011100010010000000100011;
ROM[29538] <= 32'b00000000010000010000000100010011;
ROM[29539] <= 32'b00000001010000000000001110010011;
ROM[29540] <= 32'b01000000011100011000001110110011;
ROM[29541] <= 32'b00000000000000111010000010000011;
ROM[29542] <= 32'b11111111110000010000000100010011;
ROM[29543] <= 32'b00000000000000010010001110000011;
ROM[29544] <= 32'b00000000011100100010000000100011;
ROM[29545] <= 32'b00000000010000100000000100010011;
ROM[29546] <= 32'b00000001010000000000001110010011;
ROM[29547] <= 32'b01000000011100011000001110110011;
ROM[29548] <= 32'b00000000010000111010000110000011;
ROM[29549] <= 32'b00000000100000111010001000000011;
ROM[29550] <= 32'b00000000110000111010001010000011;
ROM[29551] <= 32'b00000001000000111010001100000011;
ROM[29552] <= 32'b00000000000000001000000011100111;
ROM[29553] <= 32'b00000000000000100010001110000011;
ROM[29554] <= 32'b00000000011100010010000000100011;
ROM[29555] <= 32'b00000000010000010000000100010011;
ROM[29556] <= 32'b11111111110000010000000100010011;
ROM[29557] <= 32'b00000000000000010010001110000011;
ROM[29558] <= 32'b00001000011101101010011000100011;
ROM[29559] <= 32'b00000000000000000000001110010011;
ROM[29560] <= 32'b00000000011100010010000000100011;
ROM[29561] <= 32'b00000000010000010000000100010011;
ROM[29562] <= 32'b00000001010000000000001110010011;
ROM[29563] <= 32'b01000000011100011000001110110011;
ROM[29564] <= 32'b00000000000000111010000010000011;
ROM[29565] <= 32'b11111111110000010000000100010011;
ROM[29566] <= 32'b00000000000000010010001110000011;
ROM[29567] <= 32'b00000000011100100010000000100011;
ROM[29568] <= 32'b00000000010000100000000100010011;
ROM[29569] <= 32'b00000001010000000000001110010011;
ROM[29570] <= 32'b01000000011100011000001110110011;
ROM[29571] <= 32'b00000000010000111010000110000011;
ROM[29572] <= 32'b00000000100000111010001000000011;
ROM[29573] <= 32'b00000000110000111010001010000011;
ROM[29574] <= 32'b00000001000000111010001100000011;
ROM[29575] <= 32'b00000000000000001000000011100111;
ROM[29576] <= 32'b00001000110001101010001110000011;
ROM[29577] <= 32'b00000000011100010010000000100011;
ROM[29578] <= 32'b00000000010000010000000100010011;
ROM[29579] <= 32'b00000000000000000101001110110111;
ROM[29580] <= 32'b11110001101100111000001110010011;
ROM[29581] <= 32'b00000000011100010010000000100011;
ROM[29582] <= 32'b00000000010000010000000100010011;
ROM[29583] <= 32'b11111111110000010000000100010011;
ROM[29584] <= 32'b00000000000000010010001110000011;
ROM[29585] <= 32'b11111111110000010000000100010011;
ROM[29586] <= 32'b00000000000000010010010000000011;
ROM[29587] <= 32'b00000000011101000000001110110011;
ROM[29588] <= 32'b00000000011100010010000000100011;
ROM[29589] <= 32'b00000000010000010000000100010011;
ROM[29590] <= 32'b11111111110000010000000100010011;
ROM[29591] <= 32'b00000000000000010010001110000011;
ROM[29592] <= 32'b00001000011101101010011000100011;
ROM[29593] <= 32'b00001000110001101010001110000011;
ROM[29594] <= 32'b00000000011100010010000000100011;
ROM[29595] <= 32'b00000000010000010000000100010011;
ROM[29596] <= 32'b00000000000000000000001110010011;
ROM[29597] <= 32'b00000000011100010010000000100011;
ROM[29598] <= 32'b00000000010000010000000100010011;
ROM[29599] <= 32'b11111111110000010000000100010011;
ROM[29600] <= 32'b00000000000000010010001110000011;
ROM[29601] <= 32'b11111111110000010000000100010011;
ROM[29602] <= 32'b00000000000000010010010000000011;
ROM[29603] <= 32'b00000000011101000010001110110011;
ROM[29604] <= 32'b00000000011100010010000000100011;
ROM[29605] <= 32'b00000000010000010000000100010011;
ROM[29606] <= 32'b11111111110000010000000100010011;
ROM[29607] <= 32'b00000000000000010010001110000011;
ROM[29608] <= 32'b00000000000000111000101001100011;
ROM[29609] <= 32'b00000000000000011101001110110111;
ROM[29610] <= 32'b11101011100000111000001110010011;
ROM[29611] <= 32'b00000000111000111000001110110011;
ROM[29612] <= 32'b00000000000000111000000011100111;
ROM[29613] <= 32'b00000111000000000000000011101111;
ROM[29614] <= 32'b00001000110001101010001110000011;
ROM[29615] <= 32'b00000000011100010010000000100011;
ROM[29616] <= 32'b00000000010000010000000100010011;
ROM[29617] <= 32'b00000000000000001000001110110111;
ROM[29618] <= 32'b11111111111100111000001110010011;
ROM[29619] <= 32'b00000000011100010010000000100011;
ROM[29620] <= 32'b00000000010000010000000100010011;
ROM[29621] <= 32'b11111111110000010000000100010011;
ROM[29622] <= 32'b00000000000000010010001110000011;
ROM[29623] <= 32'b11111111110000010000000100010011;
ROM[29624] <= 32'b00000000000000010010010000000011;
ROM[29625] <= 32'b01000000011101000000001110110011;
ROM[29626] <= 32'b00000000011100010010000000100011;
ROM[29627] <= 32'b00000000010000010000000100010011;
ROM[29628] <= 32'b00000000000100000000001110010011;
ROM[29629] <= 32'b00000000011100010010000000100011;
ROM[29630] <= 32'b00000000010000010000000100010011;
ROM[29631] <= 32'b11111111110000010000000100010011;
ROM[29632] <= 32'b00000000000000010010001110000011;
ROM[29633] <= 32'b11111111110000010000000100010011;
ROM[29634] <= 32'b00000000000000010010010000000011;
ROM[29635] <= 32'b01000000011101000000001110110011;
ROM[29636] <= 32'b00000000011100010010000000100011;
ROM[29637] <= 32'b00000000010000010000000100010011;
ROM[29638] <= 32'b11111111110000010000000100010011;
ROM[29639] <= 32'b00000000000000010010001110000011;
ROM[29640] <= 32'b00001000011101101010011000100011;
ROM[29641] <= 32'b00001000110001101010001110000011;
ROM[29642] <= 32'b00000000011100010010000000100011;
ROM[29643] <= 32'b00000000010000010000000100010011;
ROM[29644] <= 32'b00000001010000000000001110010011;
ROM[29645] <= 32'b01000000011100011000001110110011;
ROM[29646] <= 32'b00000000000000111010000010000011;
ROM[29647] <= 32'b11111111110000010000000100010011;
ROM[29648] <= 32'b00000000000000010010001110000011;
ROM[29649] <= 32'b00000000011100100010000000100011;
ROM[29650] <= 32'b00000000010000100000000100010011;
ROM[29651] <= 32'b00000001010000000000001110010011;
ROM[29652] <= 32'b01000000011100011000001110110011;
ROM[29653] <= 32'b00000000010000111010000110000011;
ROM[29654] <= 32'b00000000100000111010001000000011;
ROM[29655] <= 32'b00000000110000111010001010000011;
ROM[29656] <= 32'b00000001000000111010001100000011;
ROM[29657] <= 32'b00000000000000001000000011100111;
ROM[29658] <= 32'b00000000000000010010000000100011;
ROM[29659] <= 32'b00000000010000010000000100010011;
ROM[29660] <= 32'b00000000000000010010000000100011;
ROM[29661] <= 32'b00000000010000010000000100010011;
ROM[29662] <= 32'b00000000000100000000001110010011;
ROM[29663] <= 32'b00000000011100010010000000100011;
ROM[29664] <= 32'b00000000010000010000000100010011;
ROM[29665] <= 32'b11111111110000010000000100010011;
ROM[29666] <= 32'b00000000000000010010001110000011;
ROM[29667] <= 32'b00000000011100011010000000100011;
ROM[29668] <= 32'b00000000000000011010001110000011;
ROM[29669] <= 32'b00000000011100010010000000100011;
ROM[29670] <= 32'b00000000010000010000000100010011;
ROM[29671] <= 32'b00000000000000100010001110000011;
ROM[29672] <= 32'b00000000011100010010000000100011;
ROM[29673] <= 32'b00000000010000010000000100010011;
ROM[29674] <= 32'b11111111110000010000000100010011;
ROM[29675] <= 32'b00000000000000010010001110000011;
ROM[29676] <= 32'b11111111110000010000000100010011;
ROM[29677] <= 32'b00000000000000010010010000000011;
ROM[29678] <= 32'b00000000011101000010001110110011;
ROM[29679] <= 32'b00000000011100010010000000100011;
ROM[29680] <= 32'b00000000010000010000000100010011;
ROM[29681] <= 32'b11111111110000010000000100010011;
ROM[29682] <= 32'b00000000000000010010001110000011;
ROM[29683] <= 32'b01000000011100000000001110110011;
ROM[29684] <= 32'b00000000000100111000001110010011;
ROM[29685] <= 32'b00000000011100010010000000100011;
ROM[29686] <= 32'b00000000010000010000000100010011;
ROM[29687] <= 32'b11111111110000010000000100010011;
ROM[29688] <= 32'b00000000000000010010001110000011;
ROM[29689] <= 32'b00000000000000111000101001100011;
ROM[29690] <= 32'b00000000000000011101001110110111;
ROM[29691] <= 32'b00001001010000111000001110010011;
ROM[29692] <= 32'b00000000111000111000001110110011;
ROM[29693] <= 32'b00000000000000111000000011100111;
ROM[29694] <= 32'b00000000000000011010001110000011;
ROM[29695] <= 32'b00000000011100010010000000100011;
ROM[29696] <= 32'b00000000010000010000000100010011;
ROM[29697] <= 32'b00000000001000000000001110010011;
ROM[29698] <= 32'b00000000011100010010000000100011;
ROM[29699] <= 32'b00000000010000010000000100010011;
ROM[29700] <= 32'b00000000000000011101001110110111;
ROM[29701] <= 32'b00000101110000111000001110010011;
ROM[29702] <= 32'b00000000111000111000001110110011;
ROM[29703] <= 32'b00000000011100010010000000100011;
ROM[29704] <= 32'b00000000010000010000000100010011;
ROM[29705] <= 32'b00000000001100010010000000100011;
ROM[29706] <= 32'b00000000010000010000000100010011;
ROM[29707] <= 32'b00000000010000010010000000100011;
ROM[29708] <= 32'b00000000010000010000000100010011;
ROM[29709] <= 32'b00000000010100010010000000100011;
ROM[29710] <= 32'b00000000010000010000000100010011;
ROM[29711] <= 32'b00000000011000010010000000100011;
ROM[29712] <= 32'b00000000010000010000000100010011;
ROM[29713] <= 32'b00000001010000000000001110010011;
ROM[29714] <= 32'b00000000100000111000001110010011;
ROM[29715] <= 32'b01000000011100010000001110110011;
ROM[29716] <= 32'b00000000011100000000001000110011;
ROM[29717] <= 32'b00000000001000000000000110110011;
ROM[29718] <= 32'b11111101010011110100000011101111;
ROM[29719] <= 32'b00000000000100000000001110010011;
ROM[29720] <= 32'b00000000011100010010000000100011;
ROM[29721] <= 32'b00000000010000010000000100010011;
ROM[29722] <= 32'b11111111110000010000000100010011;
ROM[29723] <= 32'b00000000000000010010001110000011;
ROM[29724] <= 32'b11111111110000010000000100010011;
ROM[29725] <= 32'b00000000000000010010010000000011;
ROM[29726] <= 32'b00000000011101000000001110110011;
ROM[29727] <= 32'b00000000011100010010000000100011;
ROM[29728] <= 32'b00000000010000010000000100010011;
ROM[29729] <= 32'b11111111110000010000000100010011;
ROM[29730] <= 32'b00000000000000010010001110000011;
ROM[29731] <= 32'b00000000011100011010000000100011;
ROM[29732] <= 32'b11110000000111111111000011101111;
ROM[29733] <= 32'b00000000000000011101001110110111;
ROM[29734] <= 32'b00001110000000111000001110010011;
ROM[29735] <= 32'b00000000111000111000001110110011;
ROM[29736] <= 32'b00000000011100010010000000100011;
ROM[29737] <= 32'b00000000010000010000000100010011;
ROM[29738] <= 32'b00000000001100010010000000100011;
ROM[29739] <= 32'b00000000010000010000000100010011;
ROM[29740] <= 32'b00000000010000010010000000100011;
ROM[29741] <= 32'b00000000010000010000000100010011;
ROM[29742] <= 32'b00000000010100010010000000100011;
ROM[29743] <= 32'b00000000010000010000000100010011;
ROM[29744] <= 32'b00000000011000010010000000100011;
ROM[29745] <= 32'b00000000010000010000000100010011;
ROM[29746] <= 32'b00000001010000000000001110010011;
ROM[29747] <= 32'b00000000000000111000001110010011;
ROM[29748] <= 32'b01000000011100010000001110110011;
ROM[29749] <= 32'b00000000011100000000001000110011;
ROM[29750] <= 32'b00000000001000000000000110110011;
ROM[29751] <= 32'b11010100010111111111000011101111;
ROM[29752] <= 32'b00000000000000011010001110000011;
ROM[29753] <= 32'b00000000011100010010000000100011;
ROM[29754] <= 32'b00000000010000010000000100010011;
ROM[29755] <= 32'b11111111110000010000000100010011;
ROM[29756] <= 32'b00000000000000010010001110000011;
ROM[29757] <= 32'b11111111110000010000000100010011;
ROM[29758] <= 32'b00000000000000010010010000000011;
ROM[29759] <= 32'b00000000011101000111001110110011;
ROM[29760] <= 32'b00000000011100010010000000100011;
ROM[29761] <= 32'b00000000010000010000000100010011;
ROM[29762] <= 32'b11111111110000010000000100010011;
ROM[29763] <= 32'b00000000000000010010001110000011;
ROM[29764] <= 32'b00000000011100011010001000100011;
ROM[29765] <= 32'b00000000010000011010001110000011;
ROM[29766] <= 32'b00000000011100010010000000100011;
ROM[29767] <= 32'b00000000010000010000000100010011;
ROM[29768] <= 32'b00000000000000100010001110000011;
ROM[29769] <= 32'b00000000011100010010000000100011;
ROM[29770] <= 32'b00000000010000010000000100010011;
ROM[29771] <= 32'b11111111110000010000000100010011;
ROM[29772] <= 32'b00000000000000010010001110000011;
ROM[29773] <= 32'b11111111110000010000000100010011;
ROM[29774] <= 32'b00000000000000010010010000000011;
ROM[29775] <= 32'b00000000100000111010001110110011;
ROM[29776] <= 32'b00000000011100010010000000100011;
ROM[29777] <= 32'b00000000010000010000000100010011;
ROM[29778] <= 32'b11111111110000010000000100010011;
ROM[29779] <= 32'b00000000000000010010001110000011;
ROM[29780] <= 32'b01000000011100000000001110110011;
ROM[29781] <= 32'b00000000000100111000001110010011;
ROM[29782] <= 32'b00000000011100010010000000100011;
ROM[29783] <= 32'b00000000010000010000000100010011;
ROM[29784] <= 32'b11111111110000010000000100010011;
ROM[29785] <= 32'b00000000000000010010001110000011;
ROM[29786] <= 32'b00000000000000111000101001100011;
ROM[29787] <= 32'b00000000000000011101001110110111;
ROM[29788] <= 32'b00100000000000111000001110010011;
ROM[29789] <= 32'b00000000111000111000001110110011;
ROM[29790] <= 32'b00000000000000111000000011100111;
ROM[29791] <= 32'b00000000000000011101001110110111;
ROM[29792] <= 32'b00011100100000111000001110010011;
ROM[29793] <= 32'b00000000111000111000001110110011;
ROM[29794] <= 32'b00000000011100010010000000100011;
ROM[29795] <= 32'b00000000010000010000000100010011;
ROM[29796] <= 32'b00000000001100010010000000100011;
ROM[29797] <= 32'b00000000010000010000000100010011;
ROM[29798] <= 32'b00000000010000010010000000100011;
ROM[29799] <= 32'b00000000010000010000000100010011;
ROM[29800] <= 32'b00000000010100010010000000100011;
ROM[29801] <= 32'b00000000010000010000000100010011;
ROM[29802] <= 32'b00000000011000010010000000100011;
ROM[29803] <= 32'b00000000010000010000000100010011;
ROM[29804] <= 32'b00000001010000000000001110010011;
ROM[29805] <= 32'b00000000000000111000001110010011;
ROM[29806] <= 32'b01000000011100010000001110110011;
ROM[29807] <= 32'b00000000011100000000001000110011;
ROM[29808] <= 32'b00000000001000000000000110110011;
ROM[29809] <= 32'b11000101110111111111000011101111;
ROM[29810] <= 32'b00000000000000011010001110000011;
ROM[29811] <= 32'b00000000011100010010000000100011;
ROM[29812] <= 32'b00000000010000010000000100010011;
ROM[29813] <= 32'b11111111110000010000000100010011;
ROM[29814] <= 32'b00000000000000010010001110000011;
ROM[29815] <= 32'b11111111110000010000000100010011;
ROM[29816] <= 32'b00000000000000010010010000000011;
ROM[29817] <= 32'b00000000011101000111001110110011;
ROM[29818] <= 32'b00000000011100010010000000100011;
ROM[29819] <= 32'b00000000010000010000000100010011;
ROM[29820] <= 32'b11111111110000010000000100010011;
ROM[29821] <= 32'b00000000000000010010001110000011;
ROM[29822] <= 32'b00000000011100011010001000100011;
ROM[29823] <= 32'b11110001100111111111000011101111;
ROM[29824] <= 32'b00000000010000011010001110000011;
ROM[29825] <= 32'b00000000011100010010000000100011;
ROM[29826] <= 32'b00000000010000010000000100010011;
ROM[29827] <= 32'b00000001010000000000001110010011;
ROM[29828] <= 32'b01000000011100011000001110110011;
ROM[29829] <= 32'b00000000000000111010000010000011;
ROM[29830] <= 32'b11111111110000010000000100010011;
ROM[29831] <= 32'b00000000000000010010001110000011;
ROM[29832] <= 32'b00000000011100100010000000100011;
ROM[29833] <= 32'b00000000010000100000000100010011;
ROM[29834] <= 32'b00000001010000000000001110010011;
ROM[29835] <= 32'b01000000011100011000001110110011;
ROM[29836] <= 32'b00000000010000111010000110000011;
ROM[29837] <= 32'b00000000100000111010001000000011;
ROM[29838] <= 32'b00000000110000111010001010000011;
ROM[29839] <= 32'b00000001000000111010001100000011;
ROM[29840] <= 32'b00000000000000001000000011100111;
ROM[29841] <= 32'b00000000000000010010000000100011;
ROM[29842] <= 32'b00000000010000010000000100010011;
ROM[29843] <= 32'b00000000000000010010000000100011;
ROM[29844] <= 32'b00000000010000010000000100010011;
ROM[29845] <= 32'b00000000000000000000001110010011;
ROM[29846] <= 32'b00000000011100010010000000100011;
ROM[29847] <= 32'b00000000010000010000000100010011;
ROM[29848] <= 32'b11111111110000010000000100010011;
ROM[29849] <= 32'b00000000000000010010001110000011;
ROM[29850] <= 32'b00000000011100011010000000100011;
ROM[29851] <= 32'b00000000000000000000001110010011;
ROM[29852] <= 32'b00000000011100010010000000100011;
ROM[29853] <= 32'b00000000010000010000000100010011;
ROM[29854] <= 32'b11111111110000010000000100010011;
ROM[29855] <= 32'b00000000000000010010001110000011;
ROM[29856] <= 32'b00000000011100011010001000100011;
ROM[29857] <= 32'b00000001010000000000001110010011;
ROM[29858] <= 32'b00000000011100010010000000100011;
ROM[29859] <= 32'b00000000010000010000000100010011;
ROM[29860] <= 32'b00000000000000011101001110110111;
ROM[29861] <= 32'b00101101110000111000001110010011;
ROM[29862] <= 32'b00000000111000111000001110110011;
ROM[29863] <= 32'b00000000011100010010000000100011;
ROM[29864] <= 32'b00000000010000010000000100010011;
ROM[29865] <= 32'b00000000001100010010000000100011;
ROM[29866] <= 32'b00000000010000010000000100010011;
ROM[29867] <= 32'b00000000010000010010000000100011;
ROM[29868] <= 32'b00000000010000010000000100010011;
ROM[29869] <= 32'b00000000010100010010000000100011;
ROM[29870] <= 32'b00000000010000010000000100010011;
ROM[29871] <= 32'b00000000011000010010000000100011;
ROM[29872] <= 32'b00000000010000010000000100010011;
ROM[29873] <= 32'b00000001010000000000001110010011;
ROM[29874] <= 32'b00000000010000111000001110010011;
ROM[29875] <= 32'b01000000011100010000001110110011;
ROM[29876] <= 32'b00000000011100000000001000110011;
ROM[29877] <= 32'b00000000001000000000000110110011;
ROM[29878] <= 32'b01000110010000001100000011101111;
ROM[29879] <= 32'b00000111000000000000001110010011;
ROM[29880] <= 32'b00000000011100010010000000100011;
ROM[29881] <= 32'b00000000010000010000000100010011;
ROM[29882] <= 32'b00000000000000011101001110110111;
ROM[29883] <= 32'b00110011010000111000001110010011;
ROM[29884] <= 32'b00000000111000111000001110110011;
ROM[29885] <= 32'b00000000011100010010000000100011;
ROM[29886] <= 32'b00000000010000010000000100010011;
ROM[29887] <= 32'b00000000001100010010000000100011;
ROM[29888] <= 32'b00000000010000010000000100010011;
ROM[29889] <= 32'b00000000010000010010000000100011;
ROM[29890] <= 32'b00000000010000010000000100010011;
ROM[29891] <= 32'b00000000010100010010000000100011;
ROM[29892] <= 32'b00000000010000010000000100010011;
ROM[29893] <= 32'b00000000011000010010000000100011;
ROM[29894] <= 32'b00000000010000010000000100010011;
ROM[29895] <= 32'b00000001010000000000001110010011;
ROM[29896] <= 32'b00000000100000111000001110010011;
ROM[29897] <= 32'b01000000011100010000001110110011;
ROM[29898] <= 32'b00000000011100000000001000110011;
ROM[29899] <= 32'b00000000001000000000000110110011;
ROM[29900] <= 32'b00000111110100001100000011101111;
ROM[29901] <= 32'b00000111001000000000001110010011;
ROM[29902] <= 32'b00000000011100010010000000100011;
ROM[29903] <= 32'b00000000010000010000000100010011;
ROM[29904] <= 32'b00000000000000011101001110110111;
ROM[29905] <= 32'b00111000110000111000001110010011;
ROM[29906] <= 32'b00000000111000111000001110110011;
ROM[29907] <= 32'b00000000011100010010000000100011;
ROM[29908] <= 32'b00000000010000010000000100010011;
ROM[29909] <= 32'b00000000001100010010000000100011;
ROM[29910] <= 32'b00000000010000010000000100010011;
ROM[29911] <= 32'b00000000010000010010000000100011;
ROM[29912] <= 32'b00000000010000010000000100010011;
ROM[29913] <= 32'b00000000010100010010000000100011;
ROM[29914] <= 32'b00000000010000010000000100010011;
ROM[29915] <= 32'b00000000011000010010000000100011;
ROM[29916] <= 32'b00000000010000010000000100010011;
ROM[29917] <= 32'b00000001010000000000001110010011;
ROM[29918] <= 32'b00000000100000111000001110010011;
ROM[29919] <= 32'b01000000011100010000001110110011;
ROM[29920] <= 32'b00000000011100000000001000110011;
ROM[29921] <= 32'b00000000001000000000000110110011;
ROM[29922] <= 32'b00000010010100001100000011101111;
ROM[29923] <= 32'b00000110010100000000001110010011;
ROM[29924] <= 32'b00000000011100010010000000100011;
ROM[29925] <= 32'b00000000010000010000000100010011;
ROM[29926] <= 32'b00000000000000011101001110110111;
ROM[29927] <= 32'b00111110010000111000001110010011;
ROM[29928] <= 32'b00000000111000111000001110110011;
ROM[29929] <= 32'b00000000011100010010000000100011;
ROM[29930] <= 32'b00000000010000010000000100010011;
ROM[29931] <= 32'b00000000001100010010000000100011;
ROM[29932] <= 32'b00000000010000010000000100010011;
ROM[29933] <= 32'b00000000010000010010000000100011;
ROM[29934] <= 32'b00000000010000010000000100010011;
ROM[29935] <= 32'b00000000010100010010000000100011;
ROM[29936] <= 32'b00000000010000010000000100010011;
ROM[29937] <= 32'b00000000011000010010000000100011;
ROM[29938] <= 32'b00000000010000010000000100010011;
ROM[29939] <= 32'b00000001010000000000001110010011;
ROM[29940] <= 32'b00000000100000111000001110010011;
ROM[29941] <= 32'b01000000011100010000001110110011;
ROM[29942] <= 32'b00000000011100000000001000110011;
ROM[29943] <= 32'b00000000001000000000000110110011;
ROM[29944] <= 32'b01111100110000001100000011101111;
ROM[29945] <= 32'b00000111001100000000001110010011;
ROM[29946] <= 32'b00000000011100010010000000100011;
ROM[29947] <= 32'b00000000010000010000000100010011;
ROM[29948] <= 32'b00000000000000011101001110110111;
ROM[29949] <= 32'b01000011110000111000001110010011;
ROM[29950] <= 32'b00000000111000111000001110110011;
ROM[29951] <= 32'b00000000011100010010000000100011;
ROM[29952] <= 32'b00000000010000010000000100010011;
ROM[29953] <= 32'b00000000001100010010000000100011;
ROM[29954] <= 32'b00000000010000010000000100010011;
ROM[29955] <= 32'b00000000010000010010000000100011;
ROM[29956] <= 32'b00000000010000010000000100010011;
ROM[29957] <= 32'b00000000010100010010000000100011;
ROM[29958] <= 32'b00000000010000010000000100010011;
ROM[29959] <= 32'b00000000011000010010000000100011;
ROM[29960] <= 32'b00000000010000010000000100010011;
ROM[29961] <= 32'b00000001010000000000001110010011;
ROM[29962] <= 32'b00000000100000111000001110010011;
ROM[29963] <= 32'b01000000011100010000001110110011;
ROM[29964] <= 32'b00000000011100000000001000110011;
ROM[29965] <= 32'b00000000001000000000000110110011;
ROM[29966] <= 32'b01110111010000001100000011101111;
ROM[29967] <= 32'b00000111001100000000001110010011;
ROM[29968] <= 32'b00000000011100010010000000100011;
ROM[29969] <= 32'b00000000010000010000000100010011;
ROM[29970] <= 32'b00000000000000011101001110110111;
ROM[29971] <= 32'b01001001010000111000001110010011;
ROM[29972] <= 32'b00000000111000111000001110110011;
ROM[29973] <= 32'b00000000011100010010000000100011;
ROM[29974] <= 32'b00000000010000010000000100010011;
ROM[29975] <= 32'b00000000001100010010000000100011;
ROM[29976] <= 32'b00000000010000010000000100010011;
ROM[29977] <= 32'b00000000010000010010000000100011;
ROM[29978] <= 32'b00000000010000010000000100010011;
ROM[29979] <= 32'b00000000010100010010000000100011;
ROM[29980] <= 32'b00000000010000010000000100010011;
ROM[29981] <= 32'b00000000011000010010000000100011;
ROM[29982] <= 32'b00000000010000010000000100010011;
ROM[29983] <= 32'b00000001010000000000001110010011;
ROM[29984] <= 32'b00000000100000111000001110010011;
ROM[29985] <= 32'b01000000011100010000001110110011;
ROM[29986] <= 32'b00000000011100000000001000110011;
ROM[29987] <= 32'b00000000001000000000000110110011;
ROM[29988] <= 32'b01110001110000001100000011101111;
ROM[29989] <= 32'b00000010000000000000001110010011;
ROM[29990] <= 32'b00000000011100010010000000100011;
ROM[29991] <= 32'b00000000010000010000000100010011;
ROM[29992] <= 32'b00000000000000011101001110110111;
ROM[29993] <= 32'b01001110110000111000001110010011;
ROM[29994] <= 32'b00000000111000111000001110110011;
ROM[29995] <= 32'b00000000011100010010000000100011;
ROM[29996] <= 32'b00000000010000010000000100010011;
ROM[29997] <= 32'b00000000001100010010000000100011;
ROM[29998] <= 32'b00000000010000010000000100010011;
ROM[29999] <= 32'b00000000010000010010000000100011;
ROM[30000] <= 32'b00000000010000010000000100010011;
ROM[30001] <= 32'b00000000010100010010000000100011;
ROM[30002] <= 32'b00000000010000010000000100010011;
ROM[30003] <= 32'b00000000011000010010000000100011;
ROM[30004] <= 32'b00000000010000010000000100010011;
ROM[30005] <= 32'b00000001010000000000001110010011;
ROM[30006] <= 32'b00000000100000111000001110010011;
ROM[30007] <= 32'b01000000011100010000001110110011;
ROM[30008] <= 32'b00000000011100000000001000110011;
ROM[30009] <= 32'b00000000001000000000000110110011;
ROM[30010] <= 32'b01101100010000001100000011101111;
ROM[30011] <= 32'b00000110000100000000001110010011;
ROM[30012] <= 32'b00000000011100010010000000100011;
ROM[30013] <= 32'b00000000010000010000000100010011;
ROM[30014] <= 32'b00000000000000011101001110110111;
ROM[30015] <= 32'b01010100010000111000001110010011;
ROM[30016] <= 32'b00000000111000111000001110110011;
ROM[30017] <= 32'b00000000011100010010000000100011;
ROM[30018] <= 32'b00000000010000010000000100010011;
ROM[30019] <= 32'b00000000001100010010000000100011;
ROM[30020] <= 32'b00000000010000010000000100010011;
ROM[30021] <= 32'b00000000010000010010000000100011;
ROM[30022] <= 32'b00000000010000010000000100010011;
ROM[30023] <= 32'b00000000010100010010000000100011;
ROM[30024] <= 32'b00000000010000010000000100010011;
ROM[30025] <= 32'b00000000011000010010000000100011;
ROM[30026] <= 32'b00000000010000010000000100010011;
ROM[30027] <= 32'b00000001010000000000001110010011;
ROM[30028] <= 32'b00000000100000111000001110010011;
ROM[30029] <= 32'b01000000011100010000001110110011;
ROM[30030] <= 32'b00000000011100000000001000110011;
ROM[30031] <= 32'b00000000001000000000000110110011;
ROM[30032] <= 32'b01100110110000001100000011101111;
ROM[30033] <= 32'b00000010000000000000001110010011;
ROM[30034] <= 32'b00000000011100010010000000100011;
ROM[30035] <= 32'b00000000010000010000000100010011;
ROM[30036] <= 32'b00000000000000011101001110110111;
ROM[30037] <= 32'b01011001110000111000001110010011;
ROM[30038] <= 32'b00000000111000111000001110110011;
ROM[30039] <= 32'b00000000011100010010000000100011;
ROM[30040] <= 32'b00000000010000010000000100010011;
ROM[30041] <= 32'b00000000001100010010000000100011;
ROM[30042] <= 32'b00000000010000010000000100010011;
ROM[30043] <= 32'b00000000010000010010000000100011;
ROM[30044] <= 32'b00000000010000010000000100010011;
ROM[30045] <= 32'b00000000010100010010000000100011;
ROM[30046] <= 32'b00000000010000010000000100010011;
ROM[30047] <= 32'b00000000011000010010000000100011;
ROM[30048] <= 32'b00000000010000010000000100010011;
ROM[30049] <= 32'b00000001010000000000001110010011;
ROM[30050] <= 32'b00000000100000111000001110010011;
ROM[30051] <= 32'b01000000011100010000001110110011;
ROM[30052] <= 32'b00000000011100000000001000110011;
ROM[30053] <= 32'b00000000001000000000000110110011;
ROM[30054] <= 32'b01100001010000001100000011101111;
ROM[30055] <= 32'b00000110101100000000001110010011;
ROM[30056] <= 32'b00000000011100010010000000100011;
ROM[30057] <= 32'b00000000010000010000000100010011;
ROM[30058] <= 32'b00000000000000011101001110110111;
ROM[30059] <= 32'b01011111010000111000001110010011;
ROM[30060] <= 32'b00000000111000111000001110110011;
ROM[30061] <= 32'b00000000011100010010000000100011;
ROM[30062] <= 32'b00000000010000010000000100010011;
ROM[30063] <= 32'b00000000001100010010000000100011;
ROM[30064] <= 32'b00000000010000010000000100010011;
ROM[30065] <= 32'b00000000010000010010000000100011;
ROM[30066] <= 32'b00000000010000010000000100010011;
ROM[30067] <= 32'b00000000010100010010000000100011;
ROM[30068] <= 32'b00000000010000010000000100010011;
ROM[30069] <= 32'b00000000011000010010000000100011;
ROM[30070] <= 32'b00000000010000010000000100010011;
ROM[30071] <= 32'b00000001010000000000001110010011;
ROM[30072] <= 32'b00000000100000111000001110010011;
ROM[30073] <= 32'b01000000011100010000001110110011;
ROM[30074] <= 32'b00000000011100000000001000110011;
ROM[30075] <= 32'b00000000001000000000000110110011;
ROM[30076] <= 32'b01011011110000001100000011101111;
ROM[30077] <= 32'b00000110010100000000001110010011;
ROM[30078] <= 32'b00000000011100010010000000100011;
ROM[30079] <= 32'b00000000010000010000000100010011;
ROM[30080] <= 32'b00000000000000011101001110110111;
ROM[30081] <= 32'b01100100110000111000001110010011;
ROM[30082] <= 32'b00000000111000111000001110110011;
ROM[30083] <= 32'b00000000011100010010000000100011;
ROM[30084] <= 32'b00000000010000010000000100010011;
ROM[30085] <= 32'b00000000001100010010000000100011;
ROM[30086] <= 32'b00000000010000010000000100010011;
ROM[30087] <= 32'b00000000010000010010000000100011;
ROM[30088] <= 32'b00000000010000010000000100010011;
ROM[30089] <= 32'b00000000010100010010000000100011;
ROM[30090] <= 32'b00000000010000010000000100010011;
ROM[30091] <= 32'b00000000011000010010000000100011;
ROM[30092] <= 32'b00000000010000010000000100010011;
ROM[30093] <= 32'b00000001010000000000001110010011;
ROM[30094] <= 32'b00000000100000111000001110010011;
ROM[30095] <= 32'b01000000011100010000001110110011;
ROM[30096] <= 32'b00000000011100000000001000110011;
ROM[30097] <= 32'b00000000001000000000000110110011;
ROM[30098] <= 32'b01010110010000001100000011101111;
ROM[30099] <= 32'b00000111100100000000001110010011;
ROM[30100] <= 32'b00000000011100010010000000100011;
ROM[30101] <= 32'b00000000010000010000000100010011;
ROM[30102] <= 32'b00000000000000011101001110110111;
ROM[30103] <= 32'b01101010010000111000001110010011;
ROM[30104] <= 32'b00000000111000111000001110110011;
ROM[30105] <= 32'b00000000011100010010000000100011;
ROM[30106] <= 32'b00000000010000010000000100010011;
ROM[30107] <= 32'b00000000001100010010000000100011;
ROM[30108] <= 32'b00000000010000010000000100010011;
ROM[30109] <= 32'b00000000010000010010000000100011;
ROM[30110] <= 32'b00000000010000010000000100010011;
ROM[30111] <= 32'b00000000010100010010000000100011;
ROM[30112] <= 32'b00000000010000010000000100010011;
ROM[30113] <= 32'b00000000011000010010000000100011;
ROM[30114] <= 32'b00000000010000010000000100010011;
ROM[30115] <= 32'b00000001010000000000001110010011;
ROM[30116] <= 32'b00000000100000111000001110010011;
ROM[30117] <= 32'b01000000011100010000001110110011;
ROM[30118] <= 32'b00000000011100000000001000110011;
ROM[30119] <= 32'b00000000001000000000000110110011;
ROM[30120] <= 32'b01010000110000001100000011101111;
ROM[30121] <= 32'b00000010000000000000001110010011;
ROM[30122] <= 32'b00000000011100010010000000100011;
ROM[30123] <= 32'b00000000010000010000000100010011;
ROM[30124] <= 32'b00000000000000011101001110110111;
ROM[30125] <= 32'b01101111110000111000001110010011;
ROM[30126] <= 32'b00000000111000111000001110110011;
ROM[30127] <= 32'b00000000011100010010000000100011;
ROM[30128] <= 32'b00000000010000010000000100010011;
ROM[30129] <= 32'b00000000001100010010000000100011;
ROM[30130] <= 32'b00000000010000010000000100010011;
ROM[30131] <= 32'b00000000010000010010000000100011;
ROM[30132] <= 32'b00000000010000010000000100010011;
ROM[30133] <= 32'b00000000010100010010000000100011;
ROM[30134] <= 32'b00000000010000010000000100010011;
ROM[30135] <= 32'b00000000011000010010000000100011;
ROM[30136] <= 32'b00000000010000010000000100010011;
ROM[30137] <= 32'b00000001010000000000001110010011;
ROM[30138] <= 32'b00000000100000111000001110010011;
ROM[30139] <= 32'b01000000011100010000001110110011;
ROM[30140] <= 32'b00000000011100000000001000110011;
ROM[30141] <= 32'b00000000001000000000000110110011;
ROM[30142] <= 32'b01001011010000001100000011101111;
ROM[30143] <= 32'b00000111010000000000001110010011;
ROM[30144] <= 32'b00000000011100010010000000100011;
ROM[30145] <= 32'b00000000010000010000000100010011;
ROM[30146] <= 32'b00000000000000011101001110110111;
ROM[30147] <= 32'b01110101010000111000001110010011;
ROM[30148] <= 32'b00000000111000111000001110110011;
ROM[30149] <= 32'b00000000011100010010000000100011;
ROM[30150] <= 32'b00000000010000010000000100010011;
ROM[30151] <= 32'b00000000001100010010000000100011;
ROM[30152] <= 32'b00000000010000010000000100010011;
ROM[30153] <= 32'b00000000010000010010000000100011;
ROM[30154] <= 32'b00000000010000010000000100010011;
ROM[30155] <= 32'b00000000010100010010000000100011;
ROM[30156] <= 32'b00000000010000010000000100010011;
ROM[30157] <= 32'b00000000011000010010000000100011;
ROM[30158] <= 32'b00000000010000010000000100010011;
ROM[30159] <= 32'b00000001010000000000001110010011;
ROM[30160] <= 32'b00000000100000111000001110010011;
ROM[30161] <= 32'b01000000011100010000001110110011;
ROM[30162] <= 32'b00000000011100000000001000110011;
ROM[30163] <= 32'b00000000001000000000000110110011;
ROM[30164] <= 32'b01000101110000001100000011101111;
ROM[30165] <= 32'b00000110111100000000001110010011;
ROM[30166] <= 32'b00000000011100010010000000100011;
ROM[30167] <= 32'b00000000010000010000000100010011;
ROM[30168] <= 32'b00000000000000011101001110110111;
ROM[30169] <= 32'b01111010110000111000001110010011;
ROM[30170] <= 32'b00000000111000111000001110110011;
ROM[30171] <= 32'b00000000011100010010000000100011;
ROM[30172] <= 32'b00000000010000010000000100010011;
ROM[30173] <= 32'b00000000001100010010000000100011;
ROM[30174] <= 32'b00000000010000010000000100010011;
ROM[30175] <= 32'b00000000010000010010000000100011;
ROM[30176] <= 32'b00000000010000010000000100010011;
ROM[30177] <= 32'b00000000010100010010000000100011;
ROM[30178] <= 32'b00000000010000010000000100010011;
ROM[30179] <= 32'b00000000011000010010000000100011;
ROM[30180] <= 32'b00000000010000010000000100010011;
ROM[30181] <= 32'b00000001010000000000001110010011;
ROM[30182] <= 32'b00000000100000111000001110010011;
ROM[30183] <= 32'b01000000011100010000001110110011;
ROM[30184] <= 32'b00000000011100000000001000110011;
ROM[30185] <= 32'b00000000001000000000000110110011;
ROM[30186] <= 32'b01000000010000001100000011101111;
ROM[30187] <= 32'b00000010000000000000001110010011;
ROM[30188] <= 32'b00000000011100010010000000100011;
ROM[30189] <= 32'b00000000010000010000000100010011;
ROM[30190] <= 32'b00000000000000011110001110110111;
ROM[30191] <= 32'b10000000010000111000001110010011;
ROM[30192] <= 32'b00000000111000111000001110110011;
ROM[30193] <= 32'b00000000011100010010000000100011;
ROM[30194] <= 32'b00000000010000010000000100010011;
ROM[30195] <= 32'b00000000001100010010000000100011;
ROM[30196] <= 32'b00000000010000010000000100010011;
ROM[30197] <= 32'b00000000010000010010000000100011;
ROM[30198] <= 32'b00000000010000010000000100010011;
ROM[30199] <= 32'b00000000010100010010000000100011;
ROM[30200] <= 32'b00000000010000010000000100010011;
ROM[30201] <= 32'b00000000011000010010000000100011;
ROM[30202] <= 32'b00000000010000010000000100010011;
ROM[30203] <= 32'b00000001010000000000001110010011;
ROM[30204] <= 32'b00000000100000111000001110010011;
ROM[30205] <= 32'b01000000011100010000001110110011;
ROM[30206] <= 32'b00000000011100000000001000110011;
ROM[30207] <= 32'b00000000001000000000000110110011;
ROM[30208] <= 32'b00111010110000001100000011101111;
ROM[30209] <= 32'b00000111001100000000001110010011;
ROM[30210] <= 32'b00000000011100010010000000100011;
ROM[30211] <= 32'b00000000010000010000000100010011;
ROM[30212] <= 32'b00000000000000011110001110110111;
ROM[30213] <= 32'b10000101110000111000001110010011;
ROM[30214] <= 32'b00000000111000111000001110110011;
ROM[30215] <= 32'b00000000011100010010000000100011;
ROM[30216] <= 32'b00000000010000010000000100010011;
ROM[30217] <= 32'b00000000001100010010000000100011;
ROM[30218] <= 32'b00000000010000010000000100010011;
ROM[30219] <= 32'b00000000010000010010000000100011;
ROM[30220] <= 32'b00000000010000010000000100010011;
ROM[30221] <= 32'b00000000010100010010000000100011;
ROM[30222] <= 32'b00000000010000010000000100010011;
ROM[30223] <= 32'b00000000011000010010000000100011;
ROM[30224] <= 32'b00000000010000010000000100010011;
ROM[30225] <= 32'b00000001010000000000001110010011;
ROM[30226] <= 32'b00000000100000111000001110010011;
ROM[30227] <= 32'b01000000011100010000001110110011;
ROM[30228] <= 32'b00000000011100000000001000110011;
ROM[30229] <= 32'b00000000001000000000000110110011;
ROM[30230] <= 32'b00110101010000001100000011101111;
ROM[30231] <= 32'b00000111010000000000001110010011;
ROM[30232] <= 32'b00000000011100010010000000100011;
ROM[30233] <= 32'b00000000010000010000000100010011;
ROM[30234] <= 32'b00000000000000011110001110110111;
ROM[30235] <= 32'b10001011010000111000001110010011;
ROM[30236] <= 32'b00000000111000111000001110110011;
ROM[30237] <= 32'b00000000011100010010000000100011;
ROM[30238] <= 32'b00000000010000010000000100010011;
ROM[30239] <= 32'b00000000001100010010000000100011;
ROM[30240] <= 32'b00000000010000010000000100010011;
ROM[30241] <= 32'b00000000010000010010000000100011;
ROM[30242] <= 32'b00000000010000010000000100010011;
ROM[30243] <= 32'b00000000010100010010000000100011;
ROM[30244] <= 32'b00000000010000010000000100010011;
ROM[30245] <= 32'b00000000011000010010000000100011;
ROM[30246] <= 32'b00000000010000010000000100010011;
ROM[30247] <= 32'b00000001010000000000001110010011;
ROM[30248] <= 32'b00000000100000111000001110010011;
ROM[30249] <= 32'b01000000011100010000001110110011;
ROM[30250] <= 32'b00000000011100000000001000110011;
ROM[30251] <= 32'b00000000001000000000000110110011;
ROM[30252] <= 32'b00101111110000001100000011101111;
ROM[30253] <= 32'b00000110000100000000001110010011;
ROM[30254] <= 32'b00000000011100010010000000100011;
ROM[30255] <= 32'b00000000010000010000000100010011;
ROM[30256] <= 32'b00000000000000011110001110110111;
ROM[30257] <= 32'b10010000110000111000001110010011;
ROM[30258] <= 32'b00000000111000111000001110110011;
ROM[30259] <= 32'b00000000011100010010000000100011;
ROM[30260] <= 32'b00000000010000010000000100010011;
ROM[30261] <= 32'b00000000001100010010000000100011;
ROM[30262] <= 32'b00000000010000010000000100010011;
ROM[30263] <= 32'b00000000010000010010000000100011;
ROM[30264] <= 32'b00000000010000010000000100010011;
ROM[30265] <= 32'b00000000010100010010000000100011;
ROM[30266] <= 32'b00000000010000010000000100010011;
ROM[30267] <= 32'b00000000011000010010000000100011;
ROM[30268] <= 32'b00000000010000010000000100010011;
ROM[30269] <= 32'b00000001010000000000001110010011;
ROM[30270] <= 32'b00000000100000111000001110010011;
ROM[30271] <= 32'b01000000011100010000001110110011;
ROM[30272] <= 32'b00000000011100000000001000110011;
ROM[30273] <= 32'b00000000001000000000000110110011;
ROM[30274] <= 32'b00101010010000001100000011101111;
ROM[30275] <= 32'b00000111001000000000001110010011;
ROM[30276] <= 32'b00000000011100010010000000100011;
ROM[30277] <= 32'b00000000010000010000000100010011;
ROM[30278] <= 32'b00000000000000011110001110110111;
ROM[30279] <= 32'b10010110010000111000001110010011;
ROM[30280] <= 32'b00000000111000111000001110110011;
ROM[30281] <= 32'b00000000011100010010000000100011;
ROM[30282] <= 32'b00000000010000010000000100010011;
ROM[30283] <= 32'b00000000001100010010000000100011;
ROM[30284] <= 32'b00000000010000010000000100010011;
ROM[30285] <= 32'b00000000010000010010000000100011;
ROM[30286] <= 32'b00000000010000010000000100010011;
ROM[30287] <= 32'b00000000010100010010000000100011;
ROM[30288] <= 32'b00000000010000010000000100010011;
ROM[30289] <= 32'b00000000011000010010000000100011;
ROM[30290] <= 32'b00000000010000010000000100010011;
ROM[30291] <= 32'b00000001010000000000001110010011;
ROM[30292] <= 32'b00000000100000111000001110010011;
ROM[30293] <= 32'b01000000011100010000001110110011;
ROM[30294] <= 32'b00000000011100000000001000110011;
ROM[30295] <= 32'b00000000001000000000000110110011;
ROM[30296] <= 32'b00100100110000001100000011101111;
ROM[30297] <= 32'b00000111010000000000001110010011;
ROM[30298] <= 32'b00000000011100010010000000100011;
ROM[30299] <= 32'b00000000010000010000000100010011;
ROM[30300] <= 32'b00000000000000011110001110110111;
ROM[30301] <= 32'b10011011110000111000001110010011;
ROM[30302] <= 32'b00000000111000111000001110110011;
ROM[30303] <= 32'b00000000011100010010000000100011;
ROM[30304] <= 32'b00000000010000010000000100010011;
ROM[30305] <= 32'b00000000001100010010000000100011;
ROM[30306] <= 32'b00000000010000010000000100010011;
ROM[30307] <= 32'b00000000010000010010000000100011;
ROM[30308] <= 32'b00000000010000010000000100010011;
ROM[30309] <= 32'b00000000010100010010000000100011;
ROM[30310] <= 32'b00000000010000010000000100010011;
ROM[30311] <= 32'b00000000011000010010000000100011;
ROM[30312] <= 32'b00000000010000010000000100010011;
ROM[30313] <= 32'b00000001010000000000001110010011;
ROM[30314] <= 32'b00000000100000111000001110010011;
ROM[30315] <= 32'b01000000011100010000001110110011;
ROM[30316] <= 32'b00000000011100000000001000110011;
ROM[30317] <= 32'b00000000001000000000000110110011;
ROM[30318] <= 32'b00011111010000001100000011101111;
ROM[30319] <= 32'b00000000000000011110001110110111;
ROM[30320] <= 32'b10100000100000111000001110010011;
ROM[30321] <= 32'b00000000111000111000001110110011;
ROM[30322] <= 32'b00000000011100010010000000100011;
ROM[30323] <= 32'b00000000010000010000000100010011;
ROM[30324] <= 32'b00000000001100010010000000100011;
ROM[30325] <= 32'b00000000010000010000000100010011;
ROM[30326] <= 32'b00000000010000010010000000100011;
ROM[30327] <= 32'b00000000010000010000000100010011;
ROM[30328] <= 32'b00000000010100010010000000100011;
ROM[30329] <= 32'b00000000010000010000000100010011;
ROM[30330] <= 32'b00000000011000010010000000100011;
ROM[30331] <= 32'b00000000010000010000000100010011;
ROM[30332] <= 32'b00000001010000000000001110010011;
ROM[30333] <= 32'b00000000010000111000001110010011;
ROM[30334] <= 32'b01000000011100010000001110110011;
ROM[30335] <= 32'b00000000011100000000001000110011;
ROM[30336] <= 32'b00000000001000000000000110110011;
ROM[30337] <= 32'b11010110010011111001000011101111;
ROM[30338] <= 32'b11111111110000010000000100010011;
ROM[30339] <= 32'b00000000000000010010001110000011;
ROM[30340] <= 32'b00000000011101100010000000100011;
ROM[30341] <= 32'b00000000000000011110001110110111;
ROM[30342] <= 32'b10100110000000111000001110010011;
ROM[30343] <= 32'b00000000111000111000001110110011;
ROM[30344] <= 32'b00000000011100010010000000100011;
ROM[30345] <= 32'b00000000010000010000000100010011;
ROM[30346] <= 32'b00000000001100010010000000100011;
ROM[30347] <= 32'b00000000010000010000000100010011;
ROM[30348] <= 32'b00000000010000010010000000100011;
ROM[30349] <= 32'b00000000010000010000000100010011;
ROM[30350] <= 32'b00000000010100010010000000100011;
ROM[30351] <= 32'b00000000010000010000000100010011;
ROM[30352] <= 32'b00000000011000010010000000100011;
ROM[30353] <= 32'b00000000010000010000000100010011;
ROM[30354] <= 32'b00000001010000000000001110010011;
ROM[30355] <= 32'b00000000000000111000001110010011;
ROM[30356] <= 32'b01000000011100010000001110110011;
ROM[30357] <= 32'b00000000011100000000001000110011;
ROM[30358] <= 32'b00000000001000000000000110110011;
ROM[30359] <= 32'b10010000110111111001000011101111;
ROM[30360] <= 32'b11111111110000010000000100010011;
ROM[30361] <= 32'b00000000000000010010001110000011;
ROM[30362] <= 32'b00000000011101100010000000100011;
ROM[30363] <= 32'b00000000010000011010001110000011;
ROM[30364] <= 32'b00000000011100010010000000100011;
ROM[30365] <= 32'b00000000010000010000000100010011;
ROM[30366] <= 32'b11111111110000010000000100010011;
ROM[30367] <= 32'b00000000000000010010001110000011;
ROM[30368] <= 32'b01000000011100000000001110110011;
ROM[30369] <= 32'b00000000000100111000001110010011;
ROM[30370] <= 32'b00000000011100010010000000100011;
ROM[30371] <= 32'b00000000010000010000000100010011;
ROM[30372] <= 32'b11111111110000010000000100010011;
ROM[30373] <= 32'b00000000000000010010001110000011;
ROM[30374] <= 32'b01000000011100000000001110110011;
ROM[30375] <= 32'b00000000000100111000001110010011;
ROM[30376] <= 32'b00000000011100010010000000100011;
ROM[30377] <= 32'b00000000010000010000000100010011;
ROM[30378] <= 32'b11111111110000010000000100010011;
ROM[30379] <= 32'b00000000000000010010001110000011;
ROM[30380] <= 32'b00000000000000111000101001100011;
ROM[30381] <= 32'b00000000000000011110001110110111;
ROM[30382] <= 32'b10111110000000111000001110010011;
ROM[30383] <= 32'b00000000111000111000001110110011;
ROM[30384] <= 32'b00000000000000111000000011100111;
ROM[30385] <= 32'b00000000000000011010001110000011;
ROM[30386] <= 32'b00000000011100010010000000100011;
ROM[30387] <= 32'b00000000010000010000000100010011;
ROM[30388] <= 32'b00000000000100000000001110010011;
ROM[30389] <= 32'b00000000011100010010000000100011;
ROM[30390] <= 32'b00000000010000010000000100010011;
ROM[30391] <= 32'b11111111110000010000000100010011;
ROM[30392] <= 32'b00000000000000010010001110000011;
ROM[30393] <= 32'b11111111110000010000000100010011;
ROM[30394] <= 32'b00000000000000010010010000000011;
ROM[30395] <= 32'b00000000011101000000001110110011;
ROM[30396] <= 32'b00000000011100010010000000100011;
ROM[30397] <= 32'b00000000010000010000000100010011;
ROM[30398] <= 32'b11111111110000010000000100010011;
ROM[30399] <= 32'b00000000000000010010001110000011;
ROM[30400] <= 32'b00000000011100011010000000100011;
ROM[30401] <= 32'b00000000000000011010001110000011;
ROM[30402] <= 32'b00000000011100010010000000100011;
ROM[30403] <= 32'b00000000010000010000000100010011;
ROM[30404] <= 32'b00000000000000001000001110110111;
ROM[30405] <= 32'b11111111111100111000001110010011;
ROM[30406] <= 32'b00000000011100010010000000100011;
ROM[30407] <= 32'b00000000010000010000000100010011;
ROM[30408] <= 32'b11111111110000010000000100010011;
ROM[30409] <= 32'b00000000000000010010001110000011;
ROM[30410] <= 32'b11111111110000010000000100010011;
ROM[30411] <= 32'b00000000000000010010010000000011;
ROM[30412] <= 32'b00000000011101000010010010110011;
ROM[30413] <= 32'b00000000100000111010010100110011;
ROM[30414] <= 32'b00000000101001001000001110110011;
ROM[30415] <= 32'b00000000000100111000001110010011;
ROM[30416] <= 32'b00000000000100111111001110010011;
ROM[30417] <= 32'b00000000011100010010000000100011;
ROM[30418] <= 32'b00000000010000010000000100010011;
ROM[30419] <= 32'b11111111110000010000000100010011;
ROM[30420] <= 32'b00000000000000010010001110000011;
ROM[30421] <= 32'b00000000000000111000101001100011;
ROM[30422] <= 32'b00000000000000011110001110110111;
ROM[30423] <= 32'b10110110110000111000001110010011;
ROM[30424] <= 32'b00000000111000111000001110110011;
ROM[30425] <= 32'b00000000000000111000000011100111;
ROM[30426] <= 32'b00000001110000000000000011101111;
ROM[30427] <= 32'b00000000000000000000001110010011;
ROM[30428] <= 32'b00000000011100010010000000100011;
ROM[30429] <= 32'b00000000010000010000000100010011;
ROM[30430] <= 32'b11111111110000010000000100010011;
ROM[30431] <= 32'b00000000000000010010001110000011;
ROM[30432] <= 32'b00000000011100011010000000100011;
ROM[30433] <= 32'b00000000000000011110001110110111;
ROM[30434] <= 32'b10111101000000111000001110010011;
ROM[30435] <= 32'b00000000111000111000001110110011;
ROM[30436] <= 32'b00000000011100010010000000100011;
ROM[30437] <= 32'b00000000010000010000000100010011;
ROM[30438] <= 32'b00000000001100010010000000100011;
ROM[30439] <= 32'b00000000010000010000000100010011;
ROM[30440] <= 32'b00000000010000010010000000100011;
ROM[30441] <= 32'b00000000010000010000000100010011;
ROM[30442] <= 32'b00000000010100010010000000100011;
ROM[30443] <= 32'b00000000010000010000000100010011;
ROM[30444] <= 32'b00000000011000010010000000100011;
ROM[30445] <= 32'b00000000010000010000000100010011;
ROM[30446] <= 32'b00000001010000000000001110010011;
ROM[30447] <= 32'b00000000000000111000001110010011;
ROM[30448] <= 32'b01000000011100010000001110110011;
ROM[30449] <= 32'b00000000011100000000001000110011;
ROM[30450] <= 32'b00000000001000000000000110110011;
ROM[30451] <= 32'b11001000110111101111000011101111;
ROM[30452] <= 32'b11111111110000010000000100010011;
ROM[30453] <= 32'b00000000000000010010001110000011;
ROM[30454] <= 32'b00000000011100011010001000100011;
ROM[30455] <= 32'b11101001000111111111000011101111;
ROM[30456] <= 32'b00000000000000011110001110110111;
ROM[30457] <= 32'b11000010110000111000001110010011;
ROM[30458] <= 32'b00000000111000111000001110110011;
ROM[30459] <= 32'b00000000011100010010000000100011;
ROM[30460] <= 32'b00000000010000010000000100010011;
ROM[30461] <= 32'b00000000001100010010000000100011;
ROM[30462] <= 32'b00000000010000010000000100010011;
ROM[30463] <= 32'b00000000010000010010000000100011;
ROM[30464] <= 32'b00000000010000010000000100010011;
ROM[30465] <= 32'b00000000010100010010000000100011;
ROM[30466] <= 32'b00000000010000010000000100010011;
ROM[30467] <= 32'b00000000011000010010000000100011;
ROM[30468] <= 32'b00000000010000010000000100010011;
ROM[30469] <= 32'b00000001010000000000001110010011;
ROM[30470] <= 32'b00000000000000111000001110010011;
ROM[30471] <= 32'b01000000011100010000001110110011;
ROM[30472] <= 32'b00000000011100000000001000110011;
ROM[30473] <= 32'b00000000001000000000000110110011;
ROM[30474] <= 32'b00100010000000000000000011101111;
ROM[30475] <= 32'b11111111110000010000000100010011;
ROM[30476] <= 32'b00000000000000010010001110000011;
ROM[30477] <= 32'b00000000011101100010000000100011;
ROM[30478] <= 32'b00000000000000011010001110000011;
ROM[30479] <= 32'b00000000011100010010000000100011;
ROM[30480] <= 32'b00000000010000010000000100010011;
ROM[30481] <= 32'b00000001010000000000001110010011;
ROM[30482] <= 32'b01000000011100011000001110110011;
ROM[30483] <= 32'b00000000000000111010000010000011;
ROM[30484] <= 32'b11111111110000010000000100010011;
ROM[30485] <= 32'b00000000000000010010001110000011;
ROM[30486] <= 32'b00000000011100100010000000100011;
ROM[30487] <= 32'b00000000010000100000000100010011;
ROM[30488] <= 32'b00000001010000000000001110010011;
ROM[30489] <= 32'b01000000011100011000001110110011;
ROM[30490] <= 32'b00000000010000111010000110000011;
ROM[30491] <= 32'b00000000100000111010001000000011;
ROM[30492] <= 32'b00000000110000111010001010000011;
ROM[30493] <= 32'b00000001000000111010001100000011;
ROM[30494] <= 32'b00000000000000001000000011100111;
ROM[30495] <= 32'b00000000000000010010000000100011;
ROM[30496] <= 32'b00000000010000010000000100010011;
ROM[30497] <= 32'b00000000110000000000001110010011;
ROM[30498] <= 32'b00000000011100010010000000100011;
ROM[30499] <= 32'b00000000010000010000000100010011;
ROM[30500] <= 32'b00000000000000011110001110110111;
ROM[30501] <= 32'b11001101110000111000001110010011;
ROM[30502] <= 32'b00000000111000111000001110110011;
ROM[30503] <= 32'b00000000011100010010000000100011;
ROM[30504] <= 32'b00000000010000010000000100010011;
ROM[30505] <= 32'b00000000001100010010000000100011;
ROM[30506] <= 32'b00000000010000010000000100010011;
ROM[30507] <= 32'b00000000010000010010000000100011;
ROM[30508] <= 32'b00000000010000010000000100010011;
ROM[30509] <= 32'b00000000010100010010000000100011;
ROM[30510] <= 32'b00000000010000010000000100010011;
ROM[30511] <= 32'b00000000011000010010000000100011;
ROM[30512] <= 32'b00000000010000010000000100010011;
ROM[30513] <= 32'b00000001010000000000001110010011;
ROM[30514] <= 32'b00000000010000111000001110010011;
ROM[30515] <= 32'b01000000011100010000001110110011;
ROM[30516] <= 32'b00000000011100000000001000110011;
ROM[30517] <= 32'b00000000001000000000000110110011;
ROM[30518] <= 32'b11001001010011110101000011101111;
ROM[30519] <= 32'b11111111110000010000000100010011;
ROM[30520] <= 32'b00000000000000010010001110000011;
ROM[30521] <= 32'b00000000011100011010000000100011;
ROM[30522] <= 32'b00000010001000000000001110010011;
ROM[30523] <= 32'b00000000011100010010000000100011;
ROM[30524] <= 32'b00000000010000010000000100010011;
ROM[30525] <= 32'b00000000000000011010001110000011;
ROM[30526] <= 32'b00000000011100010010000000100011;
ROM[30527] <= 32'b00000000010000010000000100010011;
ROM[30528] <= 32'b00000000000000011110001110110111;
ROM[30529] <= 32'b11010100110000111000001110010011;
ROM[30530] <= 32'b00000000111000111000001110110011;
ROM[30531] <= 32'b00000000011100010010000000100011;
ROM[30532] <= 32'b00000000010000010000000100010011;
ROM[30533] <= 32'b00000000001100010010000000100011;
ROM[30534] <= 32'b00000000010000010000000100010011;
ROM[30535] <= 32'b00000000010000010010000000100011;
ROM[30536] <= 32'b00000000010000010000000100010011;
ROM[30537] <= 32'b00000000010100010010000000100011;
ROM[30538] <= 32'b00000000010000010000000100010011;
ROM[30539] <= 32'b00000000011000010010000000100011;
ROM[30540] <= 32'b00000000010000010000000100010011;
ROM[30541] <= 32'b00000001010000000000001110010011;
ROM[30542] <= 32'b00000000100000111000001110010011;
ROM[30543] <= 32'b01000000011100010000001110110011;
ROM[30544] <= 32'b00000000011100000000001000110011;
ROM[30545] <= 32'b00000000001000000000000110110011;
ROM[30546] <= 32'b10101110010111110011000011101111;
ROM[30547] <= 32'b11111111110000010000000100010011;
ROM[30548] <= 32'b00000000000000010010001110000011;
ROM[30549] <= 32'b00000000011100011010000000100011;
ROM[30550] <= 32'b00000000000000011010001110000011;
ROM[30551] <= 32'b00000000011100010010000000100011;
ROM[30552] <= 32'b00000000010000010000000100010011;
ROM[30553] <= 32'b01011000000000000000001110010011;
ROM[30554] <= 32'b00000000011100010010000000100011;
ROM[30555] <= 32'b00000000010000010000000100010011;
ROM[30556] <= 32'b11111111110000010000000100010011;
ROM[30557] <= 32'b00000000000000010010001110000011;
ROM[30558] <= 32'b11111111110000010000000100010011;
ROM[30559] <= 32'b00000000000000010010010000000011;
ROM[30560] <= 32'b00000000011101000000001110110011;
ROM[30561] <= 32'b00000000011100010010000000100011;
ROM[30562] <= 32'b00000000010000010000000100010011;
ROM[30563] <= 32'b11111111110000010000000100010011;
ROM[30564] <= 32'b00000000000000010010001110000011;
ROM[30565] <= 32'b00000000011100011010000000100011;
ROM[30566] <= 32'b00000000000000000000001110010011;
ROM[30567] <= 32'b00000000011100010010000000100011;
ROM[30568] <= 32'b00000000010000010000000100010011;
ROM[30569] <= 32'b00000000000000011010001110000011;
ROM[30570] <= 32'b00000000011100010010000000100011;
ROM[30571] <= 32'b00000000010000010000000100010011;
ROM[30572] <= 32'b11111111110000010000000100010011;
ROM[30573] <= 32'b00000000000000010010001110000011;
ROM[30574] <= 32'b11111111110000010000000100010011;
ROM[30575] <= 32'b00000000000000010010010000000011;
ROM[30576] <= 32'b01000000011101000000001110110011;
ROM[30577] <= 32'b00000000011100010010000000100011;
ROM[30578] <= 32'b00000000010000010000000100010011;
ROM[30579] <= 32'b11111111110000010000000100010011;
ROM[30580] <= 32'b00000000000000010010001110000011;
ROM[30581] <= 32'b00001000011101101010100000100011;
ROM[30582] <= 32'b00000000000100000000001110010011;
ROM[30583] <= 32'b00000000011100010010000000100011;
ROM[30584] <= 32'b00000000010000010000000100010011;
ROM[30585] <= 32'b11111111110000010000000100010011;
ROM[30586] <= 32'b00000000000000010010001110000011;
ROM[30587] <= 32'b01000000011100000000001110110011;
ROM[30588] <= 32'b00000000011100010010000000100011;
ROM[30589] <= 32'b00000000010000010000000100010011;
ROM[30590] <= 32'b11111111110000010000000100010011;
ROM[30591] <= 32'b00000000000000010010001110000011;
ROM[30592] <= 32'b00001000011101101010101000100011;
ROM[30593] <= 32'b00000000000000000000001110010011;
ROM[30594] <= 32'b00000000011100010010000000100011;
ROM[30595] <= 32'b00000000010000010000000100010011;
ROM[30596] <= 32'b00000001010000000000001110010011;
ROM[30597] <= 32'b01000000011100011000001110110011;
ROM[30598] <= 32'b00000000000000111010000010000011;
ROM[30599] <= 32'b11111111110000010000000100010011;
ROM[30600] <= 32'b00000000000000010010001110000011;
ROM[30601] <= 32'b00000000011100100010000000100011;
ROM[30602] <= 32'b00000000010000100000000100010011;
ROM[30603] <= 32'b00000001010000000000001110010011;
ROM[30604] <= 32'b01000000011100011000001110110011;
ROM[30605] <= 32'b00000000010000111010000110000011;
ROM[30606] <= 32'b00000000100000111010001000000011;
ROM[30607] <= 32'b00000000110000111010001010000011;
ROM[30608] <= 32'b00000001000000111010001100000011;
ROM[30609] <= 32'b00000000000000001000000011100111;
ROM[30610] <= 32'b00000000000000010010000000100011;
ROM[30611] <= 32'b00000000010000010000000100010011;
ROM[30612] <= 32'b00000000000000010010000000100011;
ROM[30613] <= 32'b00000000010000010000000100010011;
ROM[30614] <= 32'b00000000000000000000001110010011;
ROM[30615] <= 32'b00000000011100010010000000100011;
ROM[30616] <= 32'b00000000010000010000000100010011;
ROM[30617] <= 32'b11111111110000010000000100010011;
ROM[30618] <= 32'b00000000000000010010001110000011;
ROM[30619] <= 32'b00000000011100011010000000100011;
ROM[30620] <= 32'b00000000000000011010001110000011;
ROM[30621] <= 32'b00000000011100010010000000100011;
ROM[30622] <= 32'b00000000010000010000000100010011;
ROM[30623] <= 32'b00000000000000000001001110110111;
ROM[30624] <= 32'b10010110000000111000001110010011;
ROM[30625] <= 32'b00000000011100010010000000100011;
ROM[30626] <= 32'b00000000010000010000000100010011;
ROM[30627] <= 32'b11111111110000010000000100010011;
ROM[30628] <= 32'b00000000000000010010001110000011;
ROM[30629] <= 32'b11111111110000010000000100010011;
ROM[30630] <= 32'b00000000000000010010010000000011;
ROM[30631] <= 32'b00000000011101000010001110110011;
ROM[30632] <= 32'b00000000011100010010000000100011;
ROM[30633] <= 32'b00000000010000010000000100010011;
ROM[30634] <= 32'b11111111110000010000000100010011;
ROM[30635] <= 32'b00000000000000010010001110000011;
ROM[30636] <= 32'b01000000011100000000001110110011;
ROM[30637] <= 32'b00000000000100111000001110010011;
ROM[30638] <= 32'b00000000011100010010000000100011;
ROM[30639] <= 32'b00000000010000010000000100010011;
ROM[30640] <= 32'b11111111110000010000000100010011;
ROM[30641] <= 32'b00000000000000010010001110000011;
ROM[30642] <= 32'b00000000000000111000101001100011;
ROM[30643] <= 32'b00000000000000011110001110110111;
ROM[30644] <= 32'b00000000110000111000001110010011;
ROM[30645] <= 32'b00000000111000111000001110110011;
ROM[30646] <= 32'b00000000000000111000000011100111;
ROM[30647] <= 32'b00000000000000011010001110000011;
ROM[30648] <= 32'b00000000011100010010000000100011;
ROM[30649] <= 32'b00000000010000010000000100010011;
ROM[30650] <= 32'b00000000000000011010001110000011;
ROM[30651] <= 32'b00000000011100010010000000100011;
ROM[30652] <= 32'b00000000010000010000000100010011;
ROM[30653] <= 32'b11111111110000010000000100010011;
ROM[30654] <= 32'b00000000000000010010001110000011;
ROM[30655] <= 32'b11111111110000010000000100010011;
ROM[30656] <= 32'b00000000000000010010010000000011;
ROM[30657] <= 32'b00000000011101000000001110110011;
ROM[30658] <= 32'b00000000011100010010000000100011;
ROM[30659] <= 32'b00000000010000010000000100010011;
ROM[30660] <= 32'b00000000000000011010001110000011;
ROM[30661] <= 32'b00000000011100010010000000100011;
ROM[30662] <= 32'b00000000010000010000000100010011;
ROM[30663] <= 32'b11111111110000010000000100010011;
ROM[30664] <= 32'b00000000000000010010001110000011;
ROM[30665] <= 32'b11111111110000010000000100010011;
ROM[30666] <= 32'b00000000000000010010010000000011;
ROM[30667] <= 32'b00000000011101000000001110110011;
ROM[30668] <= 32'b00000000011100010010000000100011;
ROM[30669] <= 32'b00000000010000010000000100010011;
ROM[30670] <= 32'b00000000000000011010001110000011;
ROM[30671] <= 32'b00000000011100010010000000100011;
ROM[30672] <= 32'b00000000010000010000000100010011;
ROM[30673] <= 32'b11111111110000010000000100010011;
ROM[30674] <= 32'b00000000000000010010001110000011;
ROM[30675] <= 32'b11111111110000010000000100010011;
ROM[30676] <= 32'b00000000000000010010010000000011;
ROM[30677] <= 32'b00000000011101000000001110110011;
ROM[30678] <= 32'b00000000011100010010000000100011;
ROM[30679] <= 32'b00000000010000010000000100010011;
ROM[30680] <= 32'b11111111110000010000000100010011;
ROM[30681] <= 32'b00000000000000010010001110000011;
ROM[30682] <= 32'b00000000011100011010001000100011;
ROM[30683] <= 32'b00000000000000000000001110010011;
ROM[30684] <= 32'b00000000011100010010000000100011;
ROM[30685] <= 32'b00000000010000010000000100010011;
ROM[30686] <= 32'b00001001000001101010001110000011;
ROM[30687] <= 32'b00000000011100010010000000100011;
ROM[30688] <= 32'b00000000010000010000000100010011;
ROM[30689] <= 32'b00000000010000011010001110000011;
ROM[30690] <= 32'b00000000011100010010000000100011;
ROM[30691] <= 32'b00000000010000010000000100010011;
ROM[30692] <= 32'b11111111110000010000000100010011;
ROM[30693] <= 32'b00000000000000010010001110000011;
ROM[30694] <= 32'b11111111110000010000000100010011;
ROM[30695] <= 32'b00000000000000010010010000000011;
ROM[30696] <= 32'b00000000011101000000001110110011;
ROM[30697] <= 32'b00000000011100010010000000100011;
ROM[30698] <= 32'b00000000010000010000000100010011;
ROM[30699] <= 32'b11111111110000010000000100010011;
ROM[30700] <= 32'b00000000000000010010001110000011;
ROM[30701] <= 32'b00000000000000111000001100010011;
ROM[30702] <= 32'b11111111110000010000000100010011;
ROM[30703] <= 32'b00000000000000010010001110000011;
ROM[30704] <= 32'b00000000110100110000010000110011;
ROM[30705] <= 32'b00000000011101000010000000100011;
ROM[30706] <= 32'b00000000000000011010001110000011;
ROM[30707] <= 32'b00000000011100010010000000100011;
ROM[30708] <= 32'b00000000010000010000000100010011;
ROM[30709] <= 32'b00000000000100000000001110010011;
ROM[30710] <= 32'b00000000011100010010000000100011;
ROM[30711] <= 32'b00000000010000010000000100010011;
ROM[30712] <= 32'b11111111110000010000000100010011;
ROM[30713] <= 32'b00000000000000010010001110000011;
ROM[30714] <= 32'b11111111110000010000000100010011;
ROM[30715] <= 32'b00000000000000010010010000000011;
ROM[30716] <= 32'b00000000011101000000001110110011;
ROM[30717] <= 32'b00000000011100010010000000100011;
ROM[30718] <= 32'b00000000010000010000000100010011;
ROM[30719] <= 32'b11111111110000010000000100010011;
ROM[30720] <= 32'b00000000000000010010001110000011;
ROM[30721] <= 32'b00000000011100011010000000100011;
ROM[30722] <= 32'b11100110100111111111000011101111;
ROM[30723] <= 32'b00000000000000000000001110010011;
ROM[30724] <= 32'b00000000011100010010000000100011;
ROM[30725] <= 32'b00000000010000010000000100010011;
ROM[30726] <= 32'b00000001010000000000001110010011;
ROM[30727] <= 32'b01000000011100011000001110110011;
ROM[30728] <= 32'b00000000000000111010000010000011;
ROM[30729] <= 32'b11111111110000010000000100010011;
ROM[30730] <= 32'b00000000000000010010001110000011;
ROM[30731] <= 32'b00000000011100100010000000100011;
ROM[30732] <= 32'b00000000010000100000000100010011;
ROM[30733] <= 32'b00000001010000000000001110010011;
ROM[30734] <= 32'b01000000011100011000001110110011;
ROM[30735] <= 32'b00000000010000111010000110000011;
ROM[30736] <= 32'b00000000100000111010001000000011;
ROM[30737] <= 32'b00000000110000111010001010000011;
ROM[30738] <= 32'b00000001000000111010001100000011;
ROM[30739] <= 32'b00000000000000001000000011100111;
ROM[30740] <= 32'b00000000000000100010001110000011;
ROM[30741] <= 32'b00000000011100010010000000100011;
ROM[30742] <= 32'b00000000010000010000000100010011;
ROM[30743] <= 32'b11111111110000010000000100010011;
ROM[30744] <= 32'b00000000000000010010001110000011;
ROM[30745] <= 32'b00001000011101101010101000100011;
ROM[30746] <= 32'b00000000000000000000001110010011;
ROM[30747] <= 32'b00000000011100010010000000100011;
ROM[30748] <= 32'b00000000010000010000000100010011;
ROM[30749] <= 32'b00000001010000000000001110010011;
ROM[30750] <= 32'b01000000011100011000001110110011;
ROM[30751] <= 32'b00000000000000111010000010000011;
ROM[30752] <= 32'b11111111110000010000000100010011;
ROM[30753] <= 32'b00000000000000010010001110000011;
ROM[30754] <= 32'b00000000011100100010000000100011;
ROM[30755] <= 32'b00000000010000100000000100010011;
ROM[30756] <= 32'b00000001010000000000001110010011;
ROM[30757] <= 32'b01000000011100011000001110110011;
ROM[30758] <= 32'b00000000010000111010000110000011;
ROM[30759] <= 32'b00000000100000111010001000000011;
ROM[30760] <= 32'b00000000110000111010001010000011;
ROM[30761] <= 32'b00000001000000111010001100000011;
ROM[30762] <= 32'b00000000000000001000000011100111;
ROM[30763] <= 32'b00000000000000010010000000100011;
ROM[30764] <= 32'b00000000010000010000000100010011;
ROM[30765] <= 32'b00000000000000010010000000100011;
ROM[30766] <= 32'b00000000010000010000000100010011;
ROM[30767] <= 32'b00000000000000010010000000100011;
ROM[30768] <= 32'b00000000010000010000000100010011;
ROM[30769] <= 32'b00000000000000010010000000100011;
ROM[30770] <= 32'b00000000010000010000000100010011;
ROM[30771] <= 32'b00000000000000100010001110000011;
ROM[30772] <= 32'b00000000011100010010000000100011;
ROM[30773] <= 32'b00000000010000010000000100010011;
ROM[30774] <= 32'b00000001111100000000001110010011;
ROM[30775] <= 32'b00000000011100010010000000100011;
ROM[30776] <= 32'b00000000010000010000000100010011;
ROM[30777] <= 32'b11111111110000010000000100010011;
ROM[30778] <= 32'b00000000000000010010001110000011;
ROM[30779] <= 32'b11111111110000010000000100010011;
ROM[30780] <= 32'b00000000000000010010010000000011;
ROM[30781] <= 32'b00000000011101000111001110110011;
ROM[30782] <= 32'b00000000011100010010000000100011;
ROM[30783] <= 32'b00000000010000010000000100010011;
ROM[30784] <= 32'b11111111110000010000000100010011;
ROM[30785] <= 32'b00000000000000010010001110000011;
ROM[30786] <= 32'b00000000011100011010010000100011;
ROM[30787] <= 32'b00000001111100000000001110010011;
ROM[30788] <= 32'b00000000011100010010000000100011;
ROM[30789] <= 32'b00000000010000010000000100010011;
ROM[30790] <= 32'b00000000100000011010001110000011;
ROM[30791] <= 32'b00000000011100010010000000100011;
ROM[30792] <= 32'b00000000010000010000000100010011;
ROM[30793] <= 32'b11111111110000010000000100010011;
ROM[30794] <= 32'b00000000000000010010001110000011;
ROM[30795] <= 32'b11111111110000010000000100010011;
ROM[30796] <= 32'b00000000000000010010010000000011;
ROM[30797] <= 32'b01000000011101000000001110110011;
ROM[30798] <= 32'b00000000011100010010000000100011;
ROM[30799] <= 32'b00000000010000010000000100010011;
ROM[30800] <= 32'b11111111110000010000000100010011;
ROM[30801] <= 32'b00000000000000010010001110000011;
ROM[30802] <= 32'b00000000011100011010010000100011;
ROM[30803] <= 32'b00000000010000100010001110000011;
ROM[30804] <= 32'b00000000011100010010000000100011;
ROM[30805] <= 32'b00000000010000010000000100010011;
ROM[30806] <= 32'b00000000101000000000001110010011;
ROM[30807] <= 32'b00000000011100010010000000100011;
ROM[30808] <= 32'b00000000010000010000000100010011;
ROM[30809] <= 32'b00000000000000011110001110110111;
ROM[30810] <= 32'b00011011000000111000001110010011;
ROM[30811] <= 32'b00000000111000111000001110110011;
ROM[30812] <= 32'b00000000011100010010000000100011;
ROM[30813] <= 32'b00000000010000010000000100010011;
ROM[30814] <= 32'b00000000001100010010000000100011;
ROM[30815] <= 32'b00000000010000010000000100010011;
ROM[30816] <= 32'b00000000010000010010000000100011;
ROM[30817] <= 32'b00000000010000010000000100010011;
ROM[30818] <= 32'b00000000010100010010000000100011;
ROM[30819] <= 32'b00000000010000010000000100010011;
ROM[30820] <= 32'b00000000011000010010000000100011;
ROM[30821] <= 32'b00000000010000010000000100010011;
ROM[30822] <= 32'b00000001010000000000001110010011;
ROM[30823] <= 32'b00000000100000111000001110010011;
ROM[30824] <= 32'b01000000011100010000001110110011;
ROM[30825] <= 32'b00000000011100000000001000110011;
ROM[30826] <= 32'b00000000001000000000000110110011;
ROM[30827] <= 32'b11101000000011110011000011101111;
ROM[30828] <= 32'b00000000000000100010001110000011;
ROM[30829] <= 32'b00000000011100010010000000100011;
ROM[30830] <= 32'b00000000010000010000000100010011;
ROM[30831] <= 32'b00000010000000000000001110010011;
ROM[30832] <= 32'b00000000011100010010000000100011;
ROM[30833] <= 32'b00000000010000010000000100010011;
ROM[30834] <= 32'b00000000000000011110001110110111;
ROM[30835] <= 32'b00100001010000111000001110010011;
ROM[30836] <= 32'b00000000111000111000001110110011;
ROM[30837] <= 32'b00000000011100010010000000100011;
ROM[30838] <= 32'b00000000010000010000000100010011;
ROM[30839] <= 32'b00000000001100010010000000100011;
ROM[30840] <= 32'b00000000010000010000000100010011;
ROM[30841] <= 32'b00000000010000010010000000100011;
ROM[30842] <= 32'b00000000010000010000000100010011;
ROM[30843] <= 32'b00000000010100010010000000100011;
ROM[30844] <= 32'b00000000010000010000000100010011;
ROM[30845] <= 32'b00000000011000010010000000100011;
ROM[30846] <= 32'b00000000010000010000000100010011;
ROM[30847] <= 32'b00000001010000000000001110010011;
ROM[30848] <= 32'b00000000100000111000001110010011;
ROM[30849] <= 32'b01000000011100010000001110110011;
ROM[30850] <= 32'b00000000011100000000001000110011;
ROM[30851] <= 32'b00000000001000000000000110110011;
ROM[30852] <= 32'b10011001100111110011000011101111;
ROM[30853] <= 32'b11111111110000010000000100010011;
ROM[30854] <= 32'b00000000000000010010001110000011;
ROM[30855] <= 32'b11111111110000010000000100010011;
ROM[30856] <= 32'b00000000000000010010010000000011;
ROM[30857] <= 32'b00000000011101000000001110110011;
ROM[30858] <= 32'b00000000011100010010000000100011;
ROM[30859] <= 32'b00000000010000010000000100010011;
ROM[30860] <= 32'b11111111110000010000000100010011;
ROM[30861] <= 32'b00000000000000010010001110000011;
ROM[30862] <= 32'b00000000011100011010000000100011;
ROM[30863] <= 32'b00000000000000011010001110000011;
ROM[30864] <= 32'b00000000011100010010000000100011;
ROM[30865] <= 32'b00000000010000010000000100010011;
ROM[30866] <= 32'b00000000000000011010001110000011;
ROM[30867] <= 32'b00000000011100010010000000100011;
ROM[30868] <= 32'b00000000010000010000000100010011;
ROM[30869] <= 32'b11111111110000010000000100010011;
ROM[30870] <= 32'b00000000000000010010001110000011;
ROM[30871] <= 32'b11111111110000010000000100010011;
ROM[30872] <= 32'b00000000000000010010010000000011;
ROM[30873] <= 32'b00000000011101000000001110110011;
ROM[30874] <= 32'b00000000011100010010000000100011;
ROM[30875] <= 32'b00000000010000010000000100010011;
ROM[30876] <= 32'b00000000000000011010001110000011;
ROM[30877] <= 32'b00000000011100010010000000100011;
ROM[30878] <= 32'b00000000010000010000000100010011;
ROM[30879] <= 32'b11111111110000010000000100010011;
ROM[30880] <= 32'b00000000000000010010001110000011;
ROM[30881] <= 32'b11111111110000010000000100010011;
ROM[30882] <= 32'b00000000000000010010010000000011;
ROM[30883] <= 32'b00000000011101000000001110110011;
ROM[30884] <= 32'b00000000011100010010000000100011;
ROM[30885] <= 32'b00000000010000010000000100010011;
ROM[30886] <= 32'b00000000000000011010001110000011;
ROM[30887] <= 32'b00000000011100010010000000100011;
ROM[30888] <= 32'b00000000010000010000000100010011;
ROM[30889] <= 32'b11111111110000010000000100010011;
ROM[30890] <= 32'b00000000000000010010001110000011;
ROM[30891] <= 32'b11111111110000010000000100010011;
ROM[30892] <= 32'b00000000000000010010010000000011;
ROM[30893] <= 32'b00000000011101000000001110110011;
ROM[30894] <= 32'b00000000011100010010000000100011;
ROM[30895] <= 32'b00000000010000010000000100010011;
ROM[30896] <= 32'b11111111110000010000000100010011;
ROM[30897] <= 32'b00000000000000010010001110000011;
ROM[30898] <= 32'b00000000011100011010011000100011;
ROM[30899] <= 32'b00000000100000011010001110000011;
ROM[30900] <= 32'b00000000011100010010000000100011;
ROM[30901] <= 32'b00000000010000010000000100010011;
ROM[30902] <= 32'b00000000000000011110001110110111;
ROM[30903] <= 32'b00110010010000111000001110010011;
ROM[30904] <= 32'b00000000111000111000001110110011;
ROM[30905] <= 32'b00000000011100010010000000100011;
ROM[30906] <= 32'b00000000010000010000000100010011;
ROM[30907] <= 32'b00000000001100010010000000100011;
ROM[30908] <= 32'b00000000010000010000000100010011;
ROM[30909] <= 32'b00000000010000010010000000100011;
ROM[30910] <= 32'b00000000010000010000000100010011;
ROM[30911] <= 32'b00000000010100010010000000100011;
ROM[30912] <= 32'b00000000010000010000000100010011;
ROM[30913] <= 32'b00000000011000010010000000100011;
ROM[30914] <= 32'b00000000010000010000000100010011;
ROM[30915] <= 32'b00000001010000000000001110010011;
ROM[30916] <= 32'b00000000010000111000001110010011;
ROM[30917] <= 32'b01000000011100010000001110110011;
ROM[30918] <= 32'b00000000011100000000001000110011;
ROM[30919] <= 32'b00000000001000000000000110110011;
ROM[30920] <= 32'b11100100110111110100000011101111;
ROM[30921] <= 32'b11111111110000010000000100010011;
ROM[30922] <= 32'b00000000000000010010001110000011;
ROM[30923] <= 32'b00000000011100011010001000100011;
ROM[30924] <= 32'b00001001010001101010001110000011;
ROM[30925] <= 32'b00000000011100010010000000100011;
ROM[30926] <= 32'b00000000010000010000000100010011;
ROM[30927] <= 32'b11111111110000010000000100010011;
ROM[30928] <= 32'b00000000000000010010001110000011;
ROM[30929] <= 32'b00000000000000111000101001100011;
ROM[30930] <= 32'b00000000000000011110001110110111;
ROM[30931] <= 32'b01000011110000111000001110010011;
ROM[30932] <= 32'b00000000111000111000001110110011;
ROM[30933] <= 32'b00000000000000111000000011100111;
ROM[30934] <= 32'b00001001000001101010001110000011;
ROM[30935] <= 32'b00000000011100010010000000100011;
ROM[30936] <= 32'b00000000010000010000000100010011;
ROM[30937] <= 32'b00000000110000011010001110000011;
ROM[30938] <= 32'b00000000011100010010000000100011;
ROM[30939] <= 32'b00000000010000010000000100010011;
ROM[30940] <= 32'b11111111110000010000000100010011;
ROM[30941] <= 32'b00000000000000010010001110000011;
ROM[30942] <= 32'b11111111110000010000000100010011;
ROM[30943] <= 32'b00000000000000010010010000000011;
ROM[30944] <= 32'b00000000011101000000001110110011;
ROM[30945] <= 32'b00000000011100010010000000100011;
ROM[30946] <= 32'b00000000010000010000000100010011;
ROM[30947] <= 32'b11111111110000010000000100010011;
ROM[30948] <= 32'b00000000000000010010001110000011;
ROM[30949] <= 32'b00000000000000111000001100010011;
ROM[30950] <= 32'b00000000110100110000010000110011;
ROM[30951] <= 32'b00000000000001000010001110000011;
ROM[30952] <= 32'b00000000011100010010000000100011;
ROM[30953] <= 32'b00000000010000010000000100010011;
ROM[30954] <= 32'b00000000010000011010001110000011;
ROM[30955] <= 32'b00000000011100010010000000100011;
ROM[30956] <= 32'b00000000010000010000000100010011;
ROM[30957] <= 32'b11111111110000010000000100010011;
ROM[30958] <= 32'b00000000000000010010001110000011;
ROM[30959] <= 32'b01000000011100000000001110110011;
ROM[30960] <= 32'b00000000000100111000001110010011;
ROM[30961] <= 32'b00000000011100010010000000100011;
ROM[30962] <= 32'b00000000010000010000000100010011;
ROM[30963] <= 32'b11111111110000010000000100010011;
ROM[30964] <= 32'b00000000000000010010001110000011;
ROM[30965] <= 32'b11111111110000010000000100010011;
ROM[30966] <= 32'b00000000000000010010010000000011;
ROM[30967] <= 32'b00000000011101000111001110110011;
ROM[30968] <= 32'b00000000011100010010000000100011;
ROM[30969] <= 32'b00000000010000010000000100010011;
ROM[30970] <= 32'b00001001000001101010001110000011;
ROM[30971] <= 32'b00000000011100010010000000100011;
ROM[30972] <= 32'b00000000010000010000000100010011;
ROM[30973] <= 32'b00000000110000011010001110000011;
ROM[30974] <= 32'b00000000011100010010000000100011;
ROM[30975] <= 32'b00000000010000010000000100010011;
ROM[30976] <= 32'b11111111110000010000000100010011;
ROM[30977] <= 32'b00000000000000010010001110000011;
ROM[30978] <= 32'b11111111110000010000000100010011;
ROM[30979] <= 32'b00000000000000010010010000000011;
ROM[30980] <= 32'b00000000011101000000001110110011;
ROM[30981] <= 32'b00000000011100010010000000100011;
ROM[30982] <= 32'b00000000010000010000000100010011;
ROM[30983] <= 32'b11111111110000010000000100010011;
ROM[30984] <= 32'b00000000000000010010001110000011;
ROM[30985] <= 32'b00000000000000111000001100010011;
ROM[30986] <= 32'b11111111110000010000000100010011;
ROM[30987] <= 32'b00000000000000010010001110000011;
ROM[30988] <= 32'b00000000110100110000010000110011;
ROM[30989] <= 32'b00000000011101000010000000100011;
ROM[30990] <= 32'b00001100110000000000000011101111;
ROM[30991] <= 32'b00001001000001101010001110000011;
ROM[30992] <= 32'b00000000011100010010000000100011;
ROM[30993] <= 32'b00000000010000010000000100010011;
ROM[30994] <= 32'b00000000110000011010001110000011;
ROM[30995] <= 32'b00000000011100010010000000100011;
ROM[30996] <= 32'b00000000010000010000000100010011;
ROM[30997] <= 32'b11111111110000010000000100010011;
ROM[30998] <= 32'b00000000000000010010001110000011;
ROM[30999] <= 32'b11111111110000010000000100010011;
ROM[31000] <= 32'b00000000000000010010010000000011;
ROM[31001] <= 32'b00000000011101000000001110110011;
ROM[31002] <= 32'b00000000011100010010000000100011;
ROM[31003] <= 32'b00000000010000010000000100010011;
ROM[31004] <= 32'b11111111110000010000000100010011;
ROM[31005] <= 32'b00000000000000010010001110000011;
ROM[31006] <= 32'b00000000000000111000001100010011;
ROM[31007] <= 32'b00000000110100110000010000110011;
ROM[31008] <= 32'b00000000000001000010001110000011;
ROM[31009] <= 32'b00000000011100010010000000100011;
ROM[31010] <= 32'b00000000010000010000000100010011;
ROM[31011] <= 32'b00000000010000011010001110000011;
ROM[31012] <= 32'b00000000011100010010000000100011;
ROM[31013] <= 32'b00000000010000010000000100010011;
ROM[31014] <= 32'b11111111110000010000000100010011;
ROM[31015] <= 32'b00000000000000010010001110000011;
ROM[31016] <= 32'b11111111110000010000000100010011;
ROM[31017] <= 32'b00000000000000010010010000000011;
ROM[31018] <= 32'b00000000011101000110001110110011;
ROM[31019] <= 32'b00000000011100010010000000100011;
ROM[31020] <= 32'b00000000010000010000000100010011;
ROM[31021] <= 32'b00001001000001101010001110000011;
ROM[31022] <= 32'b00000000011100010010000000100011;
ROM[31023] <= 32'b00000000010000010000000100010011;
ROM[31024] <= 32'b00000000110000011010001110000011;
ROM[31025] <= 32'b00000000011100010010000000100011;
ROM[31026] <= 32'b00000000010000010000000100010011;
ROM[31027] <= 32'b11111111110000010000000100010011;
ROM[31028] <= 32'b00000000000000010010001110000011;
ROM[31029] <= 32'b11111111110000010000000100010011;
ROM[31030] <= 32'b00000000000000010010010000000011;
ROM[31031] <= 32'b00000000011101000000001110110011;
ROM[31032] <= 32'b00000000011100010010000000100011;
ROM[31033] <= 32'b00000000010000010000000100010011;
ROM[31034] <= 32'b11111111110000010000000100010011;
ROM[31035] <= 32'b00000000000000010010001110000011;
ROM[31036] <= 32'b00000000000000111000001100010011;
ROM[31037] <= 32'b11111111110000010000000100010011;
ROM[31038] <= 32'b00000000000000010010001110000011;
ROM[31039] <= 32'b00000000110100110000010000110011;
ROM[31040] <= 32'b00000000011101000010000000100011;
ROM[31041] <= 32'b00000000000000000000001110010011;
ROM[31042] <= 32'b00000000011100010010000000100011;
ROM[31043] <= 32'b00000000010000010000000100010011;
ROM[31044] <= 32'b00000001010000000000001110010011;
ROM[31045] <= 32'b01000000011100011000001110110011;
ROM[31046] <= 32'b00000000000000111010000010000011;
ROM[31047] <= 32'b11111111110000010000000100010011;
ROM[31048] <= 32'b00000000000000010010001110000011;
ROM[31049] <= 32'b00000000011100100010000000100011;
ROM[31050] <= 32'b00000000010000100000000100010011;
ROM[31051] <= 32'b00000001010000000000001110010011;
ROM[31052] <= 32'b01000000011100011000001110110011;
ROM[31053] <= 32'b00000000010000111010000110000011;
ROM[31054] <= 32'b00000000100000111010001000000011;
ROM[31055] <= 32'b00000000110000111010001010000011;
ROM[31056] <= 32'b00000001000000111010001100000011;
ROM[31057] <= 32'b00000000000000001000000011100111;
ROM[31058] <= 32'b00000000000000010010000000100011;
ROM[31059] <= 32'b00000000010000010000000100010011;
ROM[31060] <= 32'b00000000000000010010000000100011;
ROM[31061] <= 32'b00000000010000010000000100010011;
ROM[31062] <= 32'b00000000000000010010000000100011;
ROM[31063] <= 32'b00000000010000010000000100010011;
ROM[31064] <= 32'b00000000000000010010000000100011;
ROM[31065] <= 32'b00000000010000010000000100010011;
ROM[31066] <= 32'b00000000000000010010000000100011;
ROM[31067] <= 32'b00000000010000010000000100010011;
ROM[31068] <= 32'b00000000000000010010000000100011;
ROM[31069] <= 32'b00000000010000010000000100010011;
ROM[31070] <= 32'b00000000000000100010001110000011;
ROM[31071] <= 32'b00000000011100010010000000100011;
ROM[31072] <= 32'b00000000010000010000000100010011;
ROM[31073] <= 32'b00000000100000100010001110000011;
ROM[31074] <= 32'b00000000011100010010000000100011;
ROM[31075] <= 32'b00000000010000010000000100010011;
ROM[31076] <= 32'b11111111110000010000000100010011;
ROM[31077] <= 32'b00000000000000010010001110000011;
ROM[31078] <= 32'b11111111110000010000000100010011;
ROM[31079] <= 32'b00000000000000010010010000000011;
ROM[31080] <= 32'b00000000100000111010001110110011;
ROM[31081] <= 32'b00000000011100010010000000100011;
ROM[31082] <= 32'b00000000010000010000000100010011;
ROM[31083] <= 32'b11111111110000010000000100010011;
ROM[31084] <= 32'b00000000000000010010001110000011;
ROM[31085] <= 32'b00000000000000111000101001100011;
ROM[31086] <= 32'b00000000000000011110001110110111;
ROM[31087] <= 32'b01011100110000111000001110010011;
ROM[31088] <= 32'b00000000111000111000001110110011;
ROM[31089] <= 32'b00000000000000111000000011100111;
ROM[31090] <= 32'b00001001010000000000000011101111;
ROM[31091] <= 32'b00000000000000100010001110000011;
ROM[31092] <= 32'b00000000011100010010000000100011;
ROM[31093] <= 32'b00000000010000010000000100010011;
ROM[31094] <= 32'b11111111110000010000000100010011;
ROM[31095] <= 32'b00000000000000010010001110000011;
ROM[31096] <= 32'b00000000011100011010100000100011;
ROM[31097] <= 32'b00000000100000100010001110000011;
ROM[31098] <= 32'b00000000011100010010000000100011;
ROM[31099] <= 32'b00000000010000010000000100010011;
ROM[31100] <= 32'b11111111110000010000000100010011;
ROM[31101] <= 32'b00000000000000010010001110000011;
ROM[31102] <= 32'b00000000011100100010000000100011;
ROM[31103] <= 32'b00000001000000011010001110000011;
ROM[31104] <= 32'b00000000011100010010000000100011;
ROM[31105] <= 32'b00000000010000010000000100010011;
ROM[31106] <= 32'b11111111110000010000000100010011;
ROM[31107] <= 32'b00000000000000010010001110000011;
ROM[31108] <= 32'b00000000011100100010010000100011;
ROM[31109] <= 32'b00000000010000100010001110000011;
ROM[31110] <= 32'b00000000011100010010000000100011;
ROM[31111] <= 32'b00000000010000010000000100010011;
ROM[31112] <= 32'b11111111110000010000000100010011;
ROM[31113] <= 32'b00000000000000010010001110000011;
ROM[31114] <= 32'b00000000011100011010100000100011;
ROM[31115] <= 32'b00000000110000100010001110000011;
ROM[31116] <= 32'b00000000011100010010000000100011;
ROM[31117] <= 32'b00000000010000010000000100010011;
ROM[31118] <= 32'b11111111110000010000000100010011;
ROM[31119] <= 32'b00000000000000010010001110000011;
ROM[31120] <= 32'b00000000011100100010001000100011;
ROM[31121] <= 32'b00000001000000011010001110000011;
ROM[31122] <= 32'b00000000011100010010000000100011;
ROM[31123] <= 32'b00000000010000010000000100010011;
ROM[31124] <= 32'b11111111110000010000000100010011;
ROM[31125] <= 32'b00000000000000010010001110000011;
ROM[31126] <= 32'b00000000011100100010011000100011;
ROM[31127] <= 32'b00000000100000100010001110000011;
ROM[31128] <= 32'b00000000011100010010000000100011;
ROM[31129] <= 32'b00000000010000010000000100010011;
ROM[31130] <= 32'b00000000000000100010001110000011;
ROM[31131] <= 32'b00000000011100010010000000100011;
ROM[31132] <= 32'b00000000010000010000000100010011;
ROM[31133] <= 32'b11111111110000010000000100010011;
ROM[31134] <= 32'b00000000000000010010001110000011;
ROM[31135] <= 32'b11111111110000010000000100010011;
ROM[31136] <= 32'b00000000000000010010010000000011;
ROM[31137] <= 32'b01000000011101000000001110110011;
ROM[31138] <= 32'b00000000011100010010000000100011;
ROM[31139] <= 32'b00000000010000010000000100010011;
ROM[31140] <= 32'b11111111110000010000000100010011;
ROM[31141] <= 32'b00000000000000010010001110000011;
ROM[31142] <= 32'b00000000011100011010000000100011;
ROM[31143] <= 32'b00000000110000100010001110000011;
ROM[31144] <= 32'b00000000011100010010000000100011;
ROM[31145] <= 32'b00000000010000010000000100010011;
ROM[31146] <= 32'b00000000010000100010001110000011;
ROM[31147] <= 32'b00000000011100010010000000100011;
ROM[31148] <= 32'b00000000010000010000000100010011;
ROM[31149] <= 32'b11111111110000010000000100010011;
ROM[31150] <= 32'b00000000000000010010001110000011;
ROM[31151] <= 32'b11111111110000010000000100010011;
ROM[31152] <= 32'b00000000000000010010010000000011;
ROM[31153] <= 32'b01000000011101000000001110110011;
ROM[31154] <= 32'b00000000011100010010000000100011;
ROM[31155] <= 32'b00000000010000010000000100010011;
ROM[31156] <= 32'b11111111110000010000000100010011;
ROM[31157] <= 32'b00000000000000010010001110000011;
ROM[31158] <= 32'b00000000011100011010001000100011;
ROM[31159] <= 32'b00000000000000000000001110010011;
ROM[31160] <= 32'b00000000011100010010000000100011;
ROM[31161] <= 32'b00000000010000010000000100010011;
ROM[31162] <= 32'b11111111110000010000000100010011;
ROM[31163] <= 32'b00000000000000010010001110000011;
ROM[31164] <= 32'b00000000011100011010010000100011;
ROM[31165] <= 32'b00000000000000000000001110010011;
ROM[31166] <= 32'b00000000011100010010000000100011;
ROM[31167] <= 32'b00000000010000010000000100010011;
ROM[31168] <= 32'b11111111110000010000000100010011;
ROM[31169] <= 32'b00000000000000010010001110000011;
ROM[31170] <= 32'b00000000011100011010011000100011;
ROM[31171] <= 32'b00000000010000011010001110000011;
ROM[31172] <= 32'b00000000011100010010000000100011;
ROM[31173] <= 32'b00000000010000010000000100010011;
ROM[31174] <= 32'b00000000000000000000001110010011;
ROM[31175] <= 32'b00000000011100010010000000100011;
ROM[31176] <= 32'b00000000010000010000000100010011;
ROM[31177] <= 32'b11111111110000010000000100010011;
ROM[31178] <= 32'b00000000000000010010001110000011;
ROM[31179] <= 32'b11111111110000010000000100010011;
ROM[31180] <= 32'b00000000000000010010010000000011;
ROM[31181] <= 32'b00000000011101000010010010110011;
ROM[31182] <= 32'b00000000100000111010010100110011;
ROM[31183] <= 32'b00000000101001001000001110110011;
ROM[31184] <= 32'b00000000000100111000001110010011;
ROM[31185] <= 32'b00000000000100111111001110010011;
ROM[31186] <= 32'b00000000011100010010000000100011;
ROM[31187] <= 32'b00000000010000010000000100010011;
ROM[31188] <= 32'b11111111110000010000000100010011;
ROM[31189] <= 32'b00000000000000010010001110000011;
ROM[31190] <= 32'b00000000000000111000101001100011;
ROM[31191] <= 32'b00000000000000011111001110110111;
ROM[31192] <= 32'b11101110110000111000001110010011;
ROM[31193] <= 32'b00000000111000111000001110110011;
ROM[31194] <= 32'b00000000000000111000000011100111;
ROM[31195] <= 32'b00000000000000011010001110000011;
ROM[31196] <= 32'b00000000011100010010000000100011;
ROM[31197] <= 32'b00000000010000010000000100010011;
ROM[31198] <= 32'b00000000000000000000001110010011;
ROM[31199] <= 32'b00000000011100010010000000100011;
ROM[31200] <= 32'b00000000010000010000000100010011;
ROM[31201] <= 32'b11111111110000010000000100010011;
ROM[31202] <= 32'b00000000000000010010001110000011;
ROM[31203] <= 32'b11111111110000010000000100010011;
ROM[31204] <= 32'b00000000000000010010010000000011;
ROM[31205] <= 32'b00000000011101000010010010110011;
ROM[31206] <= 32'b00000000100000111010010100110011;
ROM[31207] <= 32'b00000000101001001000001110110011;
ROM[31208] <= 32'b00000000000100111000001110010011;
ROM[31209] <= 32'b00000000000100111111001110010011;
ROM[31210] <= 32'b00000000011100010010000000100011;
ROM[31211] <= 32'b00000000010000010000000100010011;
ROM[31212] <= 32'b11111111110000010000000100010011;
ROM[31213] <= 32'b00000000000000010010001110000011;
ROM[31214] <= 32'b00000000000000111000101001100011;
ROM[31215] <= 32'b00000000000000011111001110110111;
ROM[31216] <= 32'b11100110110000111000001110010011;
ROM[31217] <= 32'b00000000111000111000001110110011;
ROM[31218] <= 32'b00000000000000111000000011100111;
ROM[31219] <= 32'b00000000000000000000001110010011;
ROM[31220] <= 32'b00000000011100010010000000100011;
ROM[31221] <= 32'b00000000010000010000000100010011;
ROM[31222] <= 32'b11111111110000010000000100010011;
ROM[31223] <= 32'b00000000000000010010001110000011;
ROM[31224] <= 32'b00000000011100011010101000100011;
ROM[31225] <= 32'b00000000010000100010001110000011;
ROM[31226] <= 32'b00000000011100010010000000100011;
ROM[31227] <= 32'b00000000010000010000000100010011;
ROM[31228] <= 32'b00000000110000100010001110000011;
ROM[31229] <= 32'b00000000011100010010000000100011;
ROM[31230] <= 32'b00000000010000010000000100010011;
ROM[31231] <= 32'b11111111110000010000000100010011;
ROM[31232] <= 32'b00000000000000010010001110000011;
ROM[31233] <= 32'b11111111110000010000000100010011;
ROM[31234] <= 32'b00000000000000010010010000000011;
ROM[31235] <= 32'b00000000011101000010001110110011;
ROM[31236] <= 32'b00000000011100010010000000100011;
ROM[31237] <= 32'b00000000010000010000000100010011;
ROM[31238] <= 32'b11111111110000010000000100010011;
ROM[31239] <= 32'b00000000000000010010001110000011;
ROM[31240] <= 32'b00000000000000111000101001100011;
ROM[31241] <= 32'b00000000000000011111001110110111;
ROM[31242] <= 32'b10110011100000111000001110010011;
ROM[31243] <= 32'b00000000111000111000001110110011;
ROM[31244] <= 32'b00000000000000111000000011100111;
ROM[31245] <= 32'b00000000100000011010001110000011;
ROM[31246] <= 32'b00000000011100010010000000100011;
ROM[31247] <= 32'b00000000010000010000000100010011;
ROM[31248] <= 32'b00000000000000011010001110000011;
ROM[31249] <= 32'b00000000011100010010000000100011;
ROM[31250] <= 32'b00000000010000010000000100010011;
ROM[31251] <= 32'b11111111110000010000000100010011;
ROM[31252] <= 32'b00000000000000010010001110000011;
ROM[31253] <= 32'b11111111110000010000000100010011;
ROM[31254] <= 32'b00000000000000010010010000000011;
ROM[31255] <= 32'b00000000100000111010001110110011;
ROM[31256] <= 32'b00000000011100010010000000100011;
ROM[31257] <= 32'b00000000010000010000000100010011;
ROM[31258] <= 32'b11111111110000010000000100010011;
ROM[31259] <= 32'b00000000000000010010001110000011;
ROM[31260] <= 32'b01000000011100000000001110110011;
ROM[31261] <= 32'b00000000000100111000001110010011;
ROM[31262] <= 32'b00000000011100010010000000100011;
ROM[31263] <= 32'b00000000010000010000000100010011;
ROM[31264] <= 32'b00000000110000011010001110000011;
ROM[31265] <= 32'b00000000011100010010000000100011;
ROM[31266] <= 32'b00000000010000010000000100010011;
ROM[31267] <= 32'b00000000010000011010001110000011;
ROM[31268] <= 32'b00000000011100010010000000100011;
ROM[31269] <= 32'b00000000010000010000000100010011;
ROM[31270] <= 32'b11111111110000010000000100010011;
ROM[31271] <= 32'b00000000000000010010001110000011;
ROM[31272] <= 32'b11111111110000010000000100010011;
ROM[31273] <= 32'b00000000000000010010010000000011;
ROM[31274] <= 32'b00000000011101000010001110110011;
ROM[31275] <= 32'b00000000011100010010000000100011;
ROM[31276] <= 32'b00000000010000010000000100010011;
ROM[31277] <= 32'b11111111110000010000000100010011;
ROM[31278] <= 32'b00000000000000010010001110000011;
ROM[31279] <= 32'b01000000011100000000001110110011;
ROM[31280] <= 32'b00000000000100111000001110010011;
ROM[31281] <= 32'b00000000011100010010000000100011;
ROM[31282] <= 32'b00000000010000010000000100010011;
ROM[31283] <= 32'b11111111110000010000000100010011;
ROM[31284] <= 32'b00000000000000010010001110000011;
ROM[31285] <= 32'b11111111110000010000000100010011;
ROM[31286] <= 32'b00000000000000010010010000000011;
ROM[31287] <= 32'b00000000011101000111001110110011;
ROM[31288] <= 32'b00000000011100010010000000100011;
ROM[31289] <= 32'b00000000010000010000000100010011;
ROM[31290] <= 32'b11111111110000010000000100010011;
ROM[31291] <= 32'b00000000000000010010001110000011;
ROM[31292] <= 32'b01000000011100000000001110110011;
ROM[31293] <= 32'b00000000000100111000001110010011;
ROM[31294] <= 32'b00000000011100010010000000100011;
ROM[31295] <= 32'b00000000010000010000000100010011;
ROM[31296] <= 32'b11111111110000010000000100010011;
ROM[31297] <= 32'b00000000000000010010001110000011;
ROM[31298] <= 32'b00000000000000111000101001100011;
ROM[31299] <= 32'b00000000000000011111001110110111;
ROM[31300] <= 32'b10110011010000111000001110010011;
ROM[31301] <= 32'b00000000111000111000001110110011;
ROM[31302] <= 32'b00000000000000111000000011100111;
ROM[31303] <= 32'b00000000000000100010001110000011;
ROM[31304] <= 32'b00000000011100010010000000100011;
ROM[31305] <= 32'b00000000010000010000000100010011;
ROM[31306] <= 32'b00000000100000011010001110000011;
ROM[31307] <= 32'b00000000011100010010000000100011;
ROM[31308] <= 32'b00000000010000010000000100010011;
ROM[31309] <= 32'b11111111110000010000000100010011;
ROM[31310] <= 32'b00000000000000010010001110000011;
ROM[31311] <= 32'b11111111110000010000000100010011;
ROM[31312] <= 32'b00000000000000010010010000000011;
ROM[31313] <= 32'b00000000011101000000001110110011;
ROM[31314] <= 32'b00000000011100010010000000100011;
ROM[31315] <= 32'b00000000010000010000000100010011;
ROM[31316] <= 32'b00000000010000100010001110000011;
ROM[31317] <= 32'b00000000011100010010000000100011;
ROM[31318] <= 32'b00000000010000010000000100010011;
ROM[31319] <= 32'b00000000110000011010001110000011;
ROM[31320] <= 32'b00000000011100010010000000100011;
ROM[31321] <= 32'b00000000010000010000000100010011;
ROM[31322] <= 32'b11111111110000010000000100010011;
ROM[31323] <= 32'b00000000000000010010001110000011;
ROM[31324] <= 32'b11111111110000010000000100010011;
ROM[31325] <= 32'b00000000000000010010010000000011;
ROM[31326] <= 32'b01000000011101000000001110110011;
ROM[31327] <= 32'b00000000011100010010000000100011;
ROM[31328] <= 32'b00000000010000010000000100010011;
ROM[31329] <= 32'b00000000000000011111001110110111;
ROM[31330] <= 32'b10011101000000111000001110010011;
ROM[31331] <= 32'b00000000111000111000001110110011;
ROM[31332] <= 32'b00000000011100010010000000100011;
ROM[31333] <= 32'b00000000010000010000000100010011;
ROM[31334] <= 32'b00000000001100010010000000100011;
ROM[31335] <= 32'b00000000010000010000000100010011;
ROM[31336] <= 32'b00000000010000010010000000100011;
ROM[31337] <= 32'b00000000010000010000000100010011;
ROM[31338] <= 32'b00000000010100010010000000100011;
ROM[31339] <= 32'b00000000010000010000000100010011;
ROM[31340] <= 32'b00000000011000010010000000100011;
ROM[31341] <= 32'b00000000010000010000000100010011;
ROM[31342] <= 32'b00000001010000000000001110010011;
ROM[31343] <= 32'b00000000100000111000001110010011;
ROM[31344] <= 32'b01000000011100010000001110110011;
ROM[31345] <= 32'b00000000011100000000001000110011;
ROM[31346] <= 32'b00000000001000000000000110110011;
ROM[31347] <= 32'b11101110000011111111000011101111;
ROM[31348] <= 32'b11111111110000010000000100010011;
ROM[31349] <= 32'b00000000000000010010001110000011;
ROM[31350] <= 32'b00000000011101100010000000100011;
ROM[31351] <= 32'b00000001010000011010001110000011;
ROM[31352] <= 32'b00000000011100010010000000100011;
ROM[31353] <= 32'b00000000010000010000000100010011;
ROM[31354] <= 32'b00000000000000000000001110010011;
ROM[31355] <= 32'b00000000011100010010000000100011;
ROM[31356] <= 32'b00000000010000010000000100010011;
ROM[31357] <= 32'b11111111110000010000000100010011;
ROM[31358] <= 32'b00000000000000010010001110000011;
ROM[31359] <= 32'b11111111110000010000000100010011;
ROM[31360] <= 32'b00000000000000010010010000000011;
ROM[31361] <= 32'b00000000100000111010001110110011;
ROM[31362] <= 32'b00000000011100010010000000100011;
ROM[31363] <= 32'b00000000010000010000000100010011;
ROM[31364] <= 32'b11111111110000010000000100010011;
ROM[31365] <= 32'b00000000000000010010001110000011;
ROM[31366] <= 32'b00000000000000111000101001100011;
ROM[31367] <= 32'b00000000000000011111001110110111;
ROM[31368] <= 32'b10101011000000111000001110010011;
ROM[31369] <= 32'b00000000111000111000001110110011;
ROM[31370] <= 32'b00000000000000111000000011100111;
ROM[31371] <= 32'b00000000110000011010001110000011;
ROM[31372] <= 32'b00000000011100010010000000100011;
ROM[31373] <= 32'b00000000010000010000000100010011;
ROM[31374] <= 32'b00000000000100000000001110010011;
ROM[31375] <= 32'b00000000011100010010000000100011;
ROM[31376] <= 32'b00000000010000010000000100010011;
ROM[31377] <= 32'b11111111110000010000000100010011;
ROM[31378] <= 32'b00000000000000010010001110000011;
ROM[31379] <= 32'b11111111110000010000000100010011;
ROM[31380] <= 32'b00000000000000010010010000000011;
ROM[31381] <= 32'b00000000011101000000001110110011;
ROM[31382] <= 32'b00000000011100010010000000100011;
ROM[31383] <= 32'b00000000010000010000000100010011;
ROM[31384] <= 32'b11111111110000010000000100010011;
ROM[31385] <= 32'b00000000000000010010001110000011;
ROM[31386] <= 32'b00000000011100011010011000100011;
ROM[31387] <= 32'b00000001010000011010001110000011;
ROM[31388] <= 32'b00000000011100010010000000100011;
ROM[31389] <= 32'b00000000010000010000000100010011;
ROM[31390] <= 32'b00000000010000011010001110000011;
ROM[31391] <= 32'b00000000011100010010000000100011;
ROM[31392] <= 32'b00000000010000010000000100010011;
ROM[31393] <= 32'b11111111110000010000000100010011;
ROM[31394] <= 32'b00000000000000010010001110000011;
ROM[31395] <= 32'b11111111110000010000000100010011;
ROM[31396] <= 32'b00000000000000010010010000000011;
ROM[31397] <= 32'b00000000011101000000001110110011;
ROM[31398] <= 32'b00000000011100010010000000100011;
ROM[31399] <= 32'b00000000010000010000000100010011;
ROM[31400] <= 32'b11111111110000010000000100010011;
ROM[31401] <= 32'b00000000000000010010001110000011;
ROM[31402] <= 32'b00000000011100011010101000100011;
ROM[31403] <= 32'b00001000010000000000000011101111;
ROM[31404] <= 32'b00000000100000011010001110000011;
ROM[31405] <= 32'b00000000011100010010000000100011;
ROM[31406] <= 32'b00000000010000010000000100010011;
ROM[31407] <= 32'b00000000000100000000001110010011;
ROM[31408] <= 32'b00000000011100010010000000100011;
ROM[31409] <= 32'b00000000010000010000000100010011;
ROM[31410] <= 32'b11111111110000010000000100010011;
ROM[31411] <= 32'b00000000000000010010001110000011;
ROM[31412] <= 32'b11111111110000010000000100010011;
ROM[31413] <= 32'b00000000000000010010010000000011;
ROM[31414] <= 32'b00000000011101000000001110110011;
ROM[31415] <= 32'b00000000011100010010000000100011;
ROM[31416] <= 32'b00000000010000010000000100010011;
ROM[31417] <= 32'b11111111110000010000000100010011;
ROM[31418] <= 32'b00000000000000010010001110000011;
ROM[31419] <= 32'b00000000011100011010010000100011;
ROM[31420] <= 32'b00000001010000011010001110000011;
ROM[31421] <= 32'b00000000011100010010000000100011;
ROM[31422] <= 32'b00000000010000010000000100010011;
ROM[31423] <= 32'b00000000000000011010001110000011;
ROM[31424] <= 32'b00000000011100010010000000100011;
ROM[31425] <= 32'b00000000010000010000000100010011;
ROM[31426] <= 32'b11111111110000010000000100010011;
ROM[31427] <= 32'b00000000000000010010001110000011;
ROM[31428] <= 32'b11111111110000010000000100010011;
ROM[31429] <= 32'b00000000000000010010010000000011;
ROM[31430] <= 32'b01000000011101000000001110110011;
ROM[31431] <= 32'b00000000011100010010000000100011;
ROM[31432] <= 32'b00000000010000010000000100010011;
ROM[31433] <= 32'b11111111110000010000000100010011;
ROM[31434] <= 32'b00000000000000010010001110000011;
ROM[31435] <= 32'b00000000011100011010101000100011;
ROM[31436] <= 32'b11010000010111111111000011101111;
ROM[31437] <= 32'b00110011010000000000000011101111;
ROM[31438] <= 32'b00000000000000000000001110010011;
ROM[31439] <= 32'b00000000011100010010000000100011;
ROM[31440] <= 32'b00000000010000010000000100010011;
ROM[31441] <= 32'b11111111110000010000000100010011;
ROM[31442] <= 32'b00000000000000010010001110000011;
ROM[31443] <= 32'b00000000011100011010010000100011;
ROM[31444] <= 32'b00000000000000000000001110010011;
ROM[31445] <= 32'b00000000011100010010000000100011;
ROM[31446] <= 32'b00000000010000010000000100010011;
ROM[31447] <= 32'b11111111110000010000000100010011;
ROM[31448] <= 32'b00000000000000010010001110000011;
ROM[31449] <= 32'b00000000011100011010011000100011;
ROM[31450] <= 32'b00000000100000011010001110000011;
ROM[31451] <= 32'b00000000011100010010000000100011;
ROM[31452] <= 32'b00000000010000010000000100010011;
ROM[31453] <= 32'b00000000000000011010001110000011;
ROM[31454] <= 32'b00000000011100010010000000100011;
ROM[31455] <= 32'b00000000010000010000000100010011;
ROM[31456] <= 32'b11111111110000010000000100010011;
ROM[31457] <= 32'b00000000000000010010001110000011;
ROM[31458] <= 32'b11111111110000010000000100010011;
ROM[31459] <= 32'b00000000000000010010010000000011;
ROM[31460] <= 32'b00000000100000111010001110110011;
ROM[31461] <= 32'b00000000011100010010000000100011;
ROM[31462] <= 32'b00000000010000010000000100010011;
ROM[31463] <= 32'b11111111110000010000000100010011;
ROM[31464] <= 32'b00000000000000010010001110000011;
ROM[31465] <= 32'b01000000011100000000001110110011;
ROM[31466] <= 32'b00000000000100111000001110010011;
ROM[31467] <= 32'b00000000011100010010000000100011;
ROM[31468] <= 32'b00000000010000010000000100010011;
ROM[31469] <= 32'b00000000110000011010001110000011;
ROM[31470] <= 32'b00000000011100010010000000100011;
ROM[31471] <= 32'b00000000010000010000000100010011;
ROM[31472] <= 32'b00000000010000011010001110000011;
ROM[31473] <= 32'b00000000011100010010000000100011;
ROM[31474] <= 32'b00000000010000010000000100010011;
ROM[31475] <= 32'b11111111110000010000000100010011;
ROM[31476] <= 32'b00000000000000010010001110000011;
ROM[31477] <= 32'b11111111110000010000000100010011;
ROM[31478] <= 32'b00000000000000010010010000000011;
ROM[31479] <= 32'b00000000100000111010001110110011;
ROM[31480] <= 32'b00000000011100010010000000100011;
ROM[31481] <= 32'b00000000010000010000000100010011;
ROM[31482] <= 32'b11111111110000010000000100010011;
ROM[31483] <= 32'b00000000000000010010001110000011;
ROM[31484] <= 32'b01000000011100000000001110110011;
ROM[31485] <= 32'b00000000000100111000001110010011;
ROM[31486] <= 32'b00000000011100010010000000100011;
ROM[31487] <= 32'b00000000010000010000000100010011;
ROM[31488] <= 32'b11111111110000010000000100010011;
ROM[31489] <= 32'b00000000000000010010001110000011;
ROM[31490] <= 32'b11111111110000010000000100010011;
ROM[31491] <= 32'b00000000000000010010010000000011;
ROM[31492] <= 32'b00000000011101000111001110110011;
ROM[31493] <= 32'b00000000011100010010000000100011;
ROM[31494] <= 32'b00000000010000010000000100010011;
ROM[31495] <= 32'b11111111110000010000000100010011;
ROM[31496] <= 32'b00000000000000010010001110000011;
ROM[31497] <= 32'b01000000011100000000001110110011;
ROM[31498] <= 32'b00000000000100111000001110010011;
ROM[31499] <= 32'b00000000011100010010000000100011;
ROM[31500] <= 32'b00000000010000010000000100010011;
ROM[31501] <= 32'b11111111110000010000000100010011;
ROM[31502] <= 32'b00000000000000010010001110000011;
ROM[31503] <= 32'b00000000000000111000101001100011;
ROM[31504] <= 32'b00000000000000011111001110110111;
ROM[31505] <= 32'b11100110100000111000001110010011;
ROM[31506] <= 32'b00000000111000111000001110110011;
ROM[31507] <= 32'b00000000000000111000000011100111;
ROM[31508] <= 32'b00000000000000100010001110000011;
ROM[31509] <= 32'b00000000011100010010000000100011;
ROM[31510] <= 32'b00000000010000010000000100010011;
ROM[31511] <= 32'b00000000100000011010001110000011;
ROM[31512] <= 32'b00000000011100010010000000100011;
ROM[31513] <= 32'b00000000010000010000000100010011;
ROM[31514] <= 32'b11111111110000010000000100010011;
ROM[31515] <= 32'b00000000000000010010001110000011;
ROM[31516] <= 32'b11111111110000010000000100010011;
ROM[31517] <= 32'b00000000000000010010010000000011;
ROM[31518] <= 32'b00000000011101000000001110110011;
ROM[31519] <= 32'b00000000011100010010000000100011;
ROM[31520] <= 32'b00000000010000010000000100010011;
ROM[31521] <= 32'b00000000010000100010001110000011;
ROM[31522] <= 32'b00000000011100010010000000100011;
ROM[31523] <= 32'b00000000010000010000000100010011;
ROM[31524] <= 32'b00000000110000011010001110000011;
ROM[31525] <= 32'b00000000011100010010000000100011;
ROM[31526] <= 32'b00000000010000010000000100010011;
ROM[31527] <= 32'b11111111110000010000000100010011;
ROM[31528] <= 32'b00000000000000010010001110000011;
ROM[31529] <= 32'b11111111110000010000000100010011;
ROM[31530] <= 32'b00000000000000010010010000000011;
ROM[31531] <= 32'b00000000011101000000001110110011;
ROM[31532] <= 32'b00000000011100010010000000100011;
ROM[31533] <= 32'b00000000010000010000000100010011;
ROM[31534] <= 32'b00000000000000011111001110110111;
ROM[31535] <= 32'b11010000010000111000001110010011;
ROM[31536] <= 32'b00000000111000111000001110110011;
ROM[31537] <= 32'b00000000011100010010000000100011;
ROM[31538] <= 32'b00000000010000010000000100010011;
ROM[31539] <= 32'b00000000001100010010000000100011;
ROM[31540] <= 32'b00000000010000010000000100010011;
ROM[31541] <= 32'b00000000010000010010000000100011;
ROM[31542] <= 32'b00000000010000010000000100010011;
ROM[31543] <= 32'b00000000010100010010000000100011;
ROM[31544] <= 32'b00000000010000010000000100010011;
ROM[31545] <= 32'b00000000011000010010000000100011;
ROM[31546] <= 32'b00000000010000010000000100010011;
ROM[31547] <= 32'b00000001010000000000001110010011;
ROM[31548] <= 32'b00000000100000111000001110010011;
ROM[31549] <= 32'b01000000011100010000001110110011;
ROM[31550] <= 32'b00000000011100000000001000110011;
ROM[31551] <= 32'b00000000001000000000000110110011;
ROM[31552] <= 32'b10111010110011111111000011101111;
ROM[31553] <= 32'b11111111110000010000000100010011;
ROM[31554] <= 32'b00000000000000010010001110000011;
ROM[31555] <= 32'b00000000011101100010000000100011;
ROM[31556] <= 32'b00000001010000011010001110000011;
ROM[31557] <= 32'b00000000011100010010000000100011;
ROM[31558] <= 32'b00000000010000010000000100010011;
ROM[31559] <= 32'b00000000000000000000001110010011;
ROM[31560] <= 32'b00000000011100010010000000100011;
ROM[31561] <= 32'b00000000010000010000000100010011;
ROM[31562] <= 32'b11111111110000010000000100010011;
ROM[31563] <= 32'b00000000000000010010001110000011;
ROM[31564] <= 32'b11111111110000010000000100010011;
ROM[31565] <= 32'b00000000000000010010010000000011;
ROM[31566] <= 32'b00000000100000111010001110110011;
ROM[31567] <= 32'b00000000011100010010000000100011;
ROM[31568] <= 32'b00000000010000010000000100010011;
ROM[31569] <= 32'b11111111110000010000000100010011;
ROM[31570] <= 32'b00000000000000010010001110000011;
ROM[31571] <= 32'b00000000000000111000101001100011;
ROM[31572] <= 32'b00000000000000011111001110110111;
ROM[31573] <= 32'b11011110010000111000001110010011;
ROM[31574] <= 32'b00000000111000111000001110110011;
ROM[31575] <= 32'b00000000000000111000000011100111;
ROM[31576] <= 32'b00000000110000011010001110000011;
ROM[31577] <= 32'b00000000011100010010000000100011;
ROM[31578] <= 32'b00000000010000010000000100010011;
ROM[31579] <= 32'b00000000000100000000001110010011;
ROM[31580] <= 32'b00000000011100010010000000100011;
ROM[31581] <= 32'b00000000010000010000000100010011;
ROM[31582] <= 32'b11111111110000010000000100010011;
ROM[31583] <= 32'b00000000000000010010001110000011;
ROM[31584] <= 32'b11111111110000010000000100010011;
ROM[31585] <= 32'b00000000000000010010010000000011;
ROM[31586] <= 32'b00000000011101000000001110110011;
ROM[31587] <= 32'b00000000011100010010000000100011;
ROM[31588] <= 32'b00000000010000010000000100010011;
ROM[31589] <= 32'b11111111110000010000000100010011;
ROM[31590] <= 32'b00000000000000010010001110000011;
ROM[31591] <= 32'b00000000011100011010011000100011;
ROM[31592] <= 32'b00000001010000011010001110000011;
ROM[31593] <= 32'b00000000011100010010000000100011;
ROM[31594] <= 32'b00000000010000010000000100010011;
ROM[31595] <= 32'b00000000010000011010001110000011;
ROM[31596] <= 32'b00000000011100010010000000100011;
ROM[31597] <= 32'b00000000010000010000000100010011;
ROM[31598] <= 32'b11111111110000010000000100010011;
ROM[31599] <= 32'b00000000000000010010001110000011;
ROM[31600] <= 32'b11111111110000010000000100010011;
ROM[31601] <= 32'b00000000000000010010010000000011;
ROM[31602] <= 32'b00000000011101000000001110110011;
ROM[31603] <= 32'b00000000011100010010000000100011;
ROM[31604] <= 32'b00000000010000010000000100010011;
ROM[31605] <= 32'b11111111110000010000000100010011;
ROM[31606] <= 32'b00000000000000010010001110000011;
ROM[31607] <= 32'b00000000011100011010101000100011;
ROM[31608] <= 32'b00001000010000000000000011101111;
ROM[31609] <= 32'b00000000100000011010001110000011;
ROM[31610] <= 32'b00000000011100010010000000100011;
ROM[31611] <= 32'b00000000010000010000000100010011;
ROM[31612] <= 32'b00000000000100000000001110010011;
ROM[31613] <= 32'b00000000011100010010000000100011;
ROM[31614] <= 32'b00000000010000010000000100010011;
ROM[31615] <= 32'b11111111110000010000000100010011;
ROM[31616] <= 32'b00000000000000010010001110000011;
ROM[31617] <= 32'b11111111110000010000000100010011;
ROM[31618] <= 32'b00000000000000010010010000000011;
ROM[31619] <= 32'b00000000011101000000001110110011;
ROM[31620] <= 32'b00000000011100010010000000100011;
ROM[31621] <= 32'b00000000010000010000000100010011;
ROM[31622] <= 32'b11111111110000010000000100010011;
ROM[31623] <= 32'b00000000000000010010001110000011;
ROM[31624] <= 32'b00000000011100011010010000100011;
ROM[31625] <= 32'b00000001010000011010001110000011;
ROM[31626] <= 32'b00000000011100010010000000100011;
ROM[31627] <= 32'b00000000010000010000000100010011;
ROM[31628] <= 32'b00000000000000011010001110000011;
ROM[31629] <= 32'b00000000011100010010000000100011;
ROM[31630] <= 32'b00000000010000010000000100010011;
ROM[31631] <= 32'b11111111110000010000000100010011;
ROM[31632] <= 32'b00000000000000010010001110000011;
ROM[31633] <= 32'b11111111110000010000000100010011;
ROM[31634] <= 32'b00000000000000010010010000000011;
ROM[31635] <= 32'b01000000011101000000001110110011;
ROM[31636] <= 32'b00000000011100010010000000100011;
ROM[31637] <= 32'b00000000010000010000000100010011;
ROM[31638] <= 32'b11111111110000010000000100010011;
ROM[31639] <= 32'b00000000000000010010001110000011;
ROM[31640] <= 32'b00000000011100011010101000100011;
ROM[31641] <= 32'b11010000010111111111000011101111;
ROM[31642] <= 32'b00001000000000000000000011101111;
ROM[31643] <= 32'b00000000000000100010001110000011;
ROM[31644] <= 32'b00000000011100010010000000100011;
ROM[31645] <= 32'b00000000010000010000000100010011;
ROM[31646] <= 32'b00000000010000100010001110000011;
ROM[31647] <= 32'b00000000011100010010000000100011;
ROM[31648] <= 32'b00000000010000010000000100010011;
ROM[31649] <= 32'b00000000110000100010001110000011;
ROM[31650] <= 32'b00000000011100010010000000100011;
ROM[31651] <= 32'b00000000010000010000000100010011;
ROM[31652] <= 32'b00000000000000011111001110110111;
ROM[31653] <= 32'b11101101110000111000001110010011;
ROM[31654] <= 32'b00000000111000111000001110110011;
ROM[31655] <= 32'b00000000011100010010000000100011;
ROM[31656] <= 32'b00000000010000010000000100010011;
ROM[31657] <= 32'b00000000001100010010000000100011;
ROM[31658] <= 32'b00000000010000010000000100010011;
ROM[31659] <= 32'b00000000010000010010000000100011;
ROM[31660] <= 32'b00000000010000010000000100010011;
ROM[31661] <= 32'b00000000010100010010000000100011;
ROM[31662] <= 32'b00000000010000010000000100010011;
ROM[31663] <= 32'b00000000011000010010000000100011;
ROM[31664] <= 32'b00000000010000010000000100010011;
ROM[31665] <= 32'b00000001010000000000001110010011;
ROM[31666] <= 32'b00000000110000111000001110010011;
ROM[31667] <= 32'b01000000011100010000001110110011;
ROM[31668] <= 32'b00000000011100000000001000110011;
ROM[31669] <= 32'b00000000001000000000000110110011;
ROM[31670] <= 32'b00101111000000000000000011101111;
ROM[31671] <= 32'b11111111110000010000000100010011;
ROM[31672] <= 32'b00000000000000010010001110000011;
ROM[31673] <= 32'b00000000011101100010000000100011;
ROM[31674] <= 32'b00001000000000000000000011101111;
ROM[31675] <= 32'b00000000000000100010001110000011;
ROM[31676] <= 32'b00000000011100010010000000100011;
ROM[31677] <= 32'b00000000010000010000000100010011;
ROM[31678] <= 32'b00000000100000100010001110000011;
ROM[31679] <= 32'b00000000011100010010000000100011;
ROM[31680] <= 32'b00000000010000010000000100010011;
ROM[31681] <= 32'b00000000010000100010001110000011;
ROM[31682] <= 32'b00000000011100010010000000100011;
ROM[31683] <= 32'b00000000010000010000000100010011;
ROM[31684] <= 32'b00000000000000011111001110110111;
ROM[31685] <= 32'b11110101110000111000001110010011;
ROM[31686] <= 32'b00000000111000111000001110110011;
ROM[31687] <= 32'b00000000011100010010000000100011;
ROM[31688] <= 32'b00000000010000010000000100010011;
ROM[31689] <= 32'b00000000001100010010000000100011;
ROM[31690] <= 32'b00000000010000010000000100010011;
ROM[31691] <= 32'b00000000010000010010000000100011;
ROM[31692] <= 32'b00000000010000010000000100010011;
ROM[31693] <= 32'b00000000010100010010000000100011;
ROM[31694] <= 32'b00000000010000010000000100010011;
ROM[31695] <= 32'b00000000011000010010000000100011;
ROM[31696] <= 32'b00000000010000010000000100010011;
ROM[31697] <= 32'b00000001010000000000001110010011;
ROM[31698] <= 32'b00000000110000111000001110010011;
ROM[31699] <= 32'b01000000011100010000001110110011;
ROM[31700] <= 32'b00000000011100000000001000110011;
ROM[31701] <= 32'b00000000001000000000000110110011;
ROM[31702] <= 32'b00000101010000000000000011101111;
ROM[31703] <= 32'b11111111110000010000000100010011;
ROM[31704] <= 32'b00000000000000010010001110000011;
ROM[31705] <= 32'b00000000011101100010000000100011;
ROM[31706] <= 32'b00000000000000000000001110010011;
ROM[31707] <= 32'b00000000011100010010000000100011;
ROM[31708] <= 32'b00000000010000010000000100010011;
ROM[31709] <= 32'b00000001010000000000001110010011;
ROM[31710] <= 32'b01000000011100011000001110110011;
ROM[31711] <= 32'b00000000000000111010000010000011;
ROM[31712] <= 32'b11111111110000010000000100010011;
ROM[31713] <= 32'b00000000000000010010001110000011;
ROM[31714] <= 32'b00000000011100100010000000100011;
ROM[31715] <= 32'b00000000010000100000000100010011;
ROM[31716] <= 32'b00000001010000000000001110010011;
ROM[31717] <= 32'b01000000011100011000001110110011;
ROM[31718] <= 32'b00000000010000111010000110000011;
ROM[31719] <= 32'b00000000100000111010001000000011;
ROM[31720] <= 32'b00000000110000111010001010000011;
ROM[31721] <= 32'b00000001000000111010001100000011;
ROM[31722] <= 32'b00000000000000001000000011100111;
ROM[31723] <= 32'b00000000000000010010000000100011;
ROM[31724] <= 32'b00000000010000010000000100010011;
ROM[31725] <= 32'b00000000000000100010001110000011;
ROM[31726] <= 32'b00000000011100010010000000100011;
ROM[31727] <= 32'b00000000010000010000000100010011;
ROM[31728] <= 32'b00000000010000100010001110000011;
ROM[31729] <= 32'b00000000011100010010000000100011;
ROM[31730] <= 32'b00000000010000010000000100010011;
ROM[31731] <= 32'b11111111110000010000000100010011;
ROM[31732] <= 32'b00000000000000010010001110000011;
ROM[31733] <= 32'b11111111110000010000000100010011;
ROM[31734] <= 32'b00000000000000010010010000000011;
ROM[31735] <= 32'b00000000100000111010001110110011;
ROM[31736] <= 32'b00000000011100010010000000100011;
ROM[31737] <= 32'b00000000010000010000000100010011;
ROM[31738] <= 32'b11111111110000010000000100010011;
ROM[31739] <= 32'b00000000000000010010001110000011;
ROM[31740] <= 32'b00000000000000111000101001100011;
ROM[31741] <= 32'b00000000000000011111001110110111;
ROM[31742] <= 32'b00000000100000111000001110010011;
ROM[31743] <= 32'b00000000111000111000001110110011;
ROM[31744] <= 32'b00000000000000111000000011100111;
ROM[31745] <= 32'b00000100110000000000000011101111;
ROM[31746] <= 32'b00000000000000100010001110000011;
ROM[31747] <= 32'b00000000011100010010000000100011;
ROM[31748] <= 32'b00000000010000010000000100010011;
ROM[31749] <= 32'b11111111110000010000000100010011;
ROM[31750] <= 32'b00000000000000010010001110000011;
ROM[31751] <= 32'b00000000011100011010000000100011;
ROM[31752] <= 32'b00000000010000100010001110000011;
ROM[31753] <= 32'b00000000011100010010000000100011;
ROM[31754] <= 32'b00000000010000010000000100010011;
ROM[31755] <= 32'b11111111110000010000000100010011;
ROM[31756] <= 32'b00000000000000010010001110000011;
ROM[31757] <= 32'b00000000011100100010000000100011;
ROM[31758] <= 32'b00000000000000011010001110000011;
ROM[31759] <= 32'b00000000011100010010000000100011;
ROM[31760] <= 32'b00000000010000010000000100010011;
ROM[31761] <= 32'b11111111110000010000000100010011;
ROM[31762] <= 32'b00000000000000010010001110000011;
ROM[31763] <= 32'b00000000011100100010001000100011;
ROM[31764] <= 32'b00000000010000100010001110000011;
ROM[31765] <= 32'b00000000011100010010000000100011;
ROM[31766] <= 32'b00000000010000010000000100010011;
ROM[31767] <= 32'b00000000000000100010001110000011;
ROM[31768] <= 32'b00000000011100010010000000100011;
ROM[31769] <= 32'b00000000010000010000000100010011;
ROM[31770] <= 32'b11111111110000010000000100010011;
ROM[31771] <= 32'b00000000000000010010001110000011;
ROM[31772] <= 32'b11111111110000010000000100010011;
ROM[31773] <= 32'b00000000000000010010010000000011;
ROM[31774] <= 32'b00000000011101000010001110110011;
ROM[31775] <= 32'b00000000011100010010000000100011;
ROM[31776] <= 32'b00000000010000010000000100010011;
ROM[31777] <= 32'b11111111110000010000000100010011;
ROM[31778] <= 32'b00000000000000010010001110000011;
ROM[31779] <= 32'b01000000011100000000001110110011;
ROM[31780] <= 32'b00000000000100111000001110010011;
ROM[31781] <= 32'b00000000011100010010000000100011;
ROM[31782] <= 32'b00000000010000010000000100010011;
ROM[31783] <= 32'b11111111110000010000000100010011;
ROM[31784] <= 32'b00000000000000010010001110000011;
ROM[31785] <= 32'b01000000011100000000001110110011;
ROM[31786] <= 32'b00000000000100111000001110010011;
ROM[31787] <= 32'b00000000011100010010000000100011;
ROM[31788] <= 32'b00000000010000010000000100010011;
ROM[31789] <= 32'b11111111110000010000000100010011;
ROM[31790] <= 32'b00000000000000010010001110000011;
ROM[31791] <= 32'b00000000000000111000101001100011;
ROM[31792] <= 32'b00000000000000011111001110110111;
ROM[31793] <= 32'b00011000010000111000001110010011;
ROM[31794] <= 32'b00000000111000111000001110110011;
ROM[31795] <= 32'b00000000000000111000000011100111;
ROM[31796] <= 32'b00000000000000100010001110000011;
ROM[31797] <= 32'b00000000011100010010000000100011;
ROM[31798] <= 32'b00000000010000010000000100010011;
ROM[31799] <= 32'b00000000100000100010001110000011;
ROM[31800] <= 32'b00000000011100010010000000100011;
ROM[31801] <= 32'b00000000010000010000000100010011;
ROM[31802] <= 32'b00000000000000011111001110110111;
ROM[31803] <= 32'b00010011010000111000001110010011;
ROM[31804] <= 32'b00000000111000111000001110110011;
ROM[31805] <= 32'b00000000011100010010000000100011;
ROM[31806] <= 32'b00000000010000010000000100010011;
ROM[31807] <= 32'b00000000001100010010000000100011;
ROM[31808] <= 32'b00000000010000010000000100010011;
ROM[31809] <= 32'b00000000010000010010000000100011;
ROM[31810] <= 32'b00000000010000010000000100010011;
ROM[31811] <= 32'b00000000010100010010000000100011;
ROM[31812] <= 32'b00000000010000010000000100010011;
ROM[31813] <= 32'b00000000011000010010000000100011;
ROM[31814] <= 32'b00000000010000010000000100010011;
ROM[31815] <= 32'b00000001010000000000001110010011;
ROM[31816] <= 32'b00000000100000111000001110010011;
ROM[31817] <= 32'b01000000011100010000001110110011;
ROM[31818] <= 32'b00000000011100000000001000110011;
ROM[31819] <= 32'b00000000001000000000000110110011;
ROM[31820] <= 32'b11110111110111111110000011101111;
ROM[31821] <= 32'b11111111110000010000000100010011;
ROM[31822] <= 32'b00000000000000010010001110000011;
ROM[31823] <= 32'b00000000011101100010000000100011;
ROM[31824] <= 32'b00000000000000100010001110000011;
ROM[31825] <= 32'b00000000011100010010000000100011;
ROM[31826] <= 32'b00000000010000010000000100010011;
ROM[31827] <= 32'b00000000000100000000001110010011;
ROM[31828] <= 32'b00000000011100010010000000100011;
ROM[31829] <= 32'b00000000010000010000000100010011;
ROM[31830] <= 32'b11111111110000010000000100010011;
ROM[31831] <= 32'b00000000000000010010001110000011;
ROM[31832] <= 32'b11111111110000010000000100010011;
ROM[31833] <= 32'b00000000000000010010010000000011;
ROM[31834] <= 32'b00000000011101000000001110110011;
ROM[31835] <= 32'b00000000011100010010000000100011;
ROM[31836] <= 32'b00000000010000010000000100010011;
ROM[31837] <= 32'b11111111110000010000000100010011;
ROM[31838] <= 32'b00000000000000010010001110000011;
ROM[31839] <= 32'b00000000011100100010000000100011;
ROM[31840] <= 32'b11101101000111111111000011101111;
ROM[31841] <= 32'b00000000000000000000001110010011;
ROM[31842] <= 32'b00000000011100010010000000100011;
ROM[31843] <= 32'b00000000010000010000000100010011;
ROM[31844] <= 32'b00000001010000000000001110010011;
ROM[31845] <= 32'b01000000011100011000001110110011;
ROM[31846] <= 32'b00000000000000111010000010000011;
ROM[31847] <= 32'b11111111110000010000000100010011;
ROM[31848] <= 32'b00000000000000010010001110000011;
ROM[31849] <= 32'b00000000011100100010000000100011;
ROM[31850] <= 32'b00000000010000100000000100010011;
ROM[31851] <= 32'b00000001010000000000001110010011;
ROM[31852] <= 32'b01000000011100011000001110110011;
ROM[31853] <= 32'b00000000010000111010000110000011;
ROM[31854] <= 32'b00000000100000111010001000000011;
ROM[31855] <= 32'b00000000110000111010001010000011;
ROM[31856] <= 32'b00000001000000111010001100000011;
ROM[31857] <= 32'b00000000000000001000000011100111;
ROM[31858] <= 32'b00000000000000010010000000100011;
ROM[31859] <= 32'b00000000010000010000000100010011;
ROM[31860] <= 32'b00000000010000100010001110000011;
ROM[31861] <= 32'b00000000011100010010000000100011;
ROM[31862] <= 32'b00000000010000010000000100010011;
ROM[31863] <= 32'b00000000100000100010001110000011;
ROM[31864] <= 32'b00000000011100010010000000100011;
ROM[31865] <= 32'b00000000010000010000000100010011;
ROM[31866] <= 32'b11111111110000010000000100010011;
ROM[31867] <= 32'b00000000000000010010001110000011;
ROM[31868] <= 32'b11111111110000010000000100010011;
ROM[31869] <= 32'b00000000000000010010010000000011;
ROM[31870] <= 32'b00000000100000111010001110110011;
ROM[31871] <= 32'b00000000011100010010000000100011;
ROM[31872] <= 32'b00000000010000010000000100010011;
ROM[31873] <= 32'b11111111110000010000000100010011;
ROM[31874] <= 32'b00000000000000010010001110000011;
ROM[31875] <= 32'b00000000000000111000101001100011;
ROM[31876] <= 32'b00000000000000011111001110110111;
ROM[31877] <= 32'b00100010010000111000001110010011;
ROM[31878] <= 32'b00000000111000111000001110110011;
ROM[31879] <= 32'b00000000000000111000000011100111;
ROM[31880] <= 32'b00000100110000000000000011101111;
ROM[31881] <= 32'b00000000010000100010001110000011;
ROM[31882] <= 32'b00000000011100010010000000100011;
ROM[31883] <= 32'b00000000010000010000000100010011;
ROM[31884] <= 32'b11111111110000010000000100010011;
ROM[31885] <= 32'b00000000000000010010001110000011;
ROM[31886] <= 32'b00000000011100011010000000100011;
ROM[31887] <= 32'b00000000100000100010001110000011;
ROM[31888] <= 32'b00000000011100010010000000100011;
ROM[31889] <= 32'b00000000010000010000000100010011;
ROM[31890] <= 32'b11111111110000010000000100010011;
ROM[31891] <= 32'b00000000000000010010001110000011;
ROM[31892] <= 32'b00000000011100100010001000100011;
ROM[31893] <= 32'b00000000000000011010001110000011;
ROM[31894] <= 32'b00000000011100010010000000100011;
ROM[31895] <= 32'b00000000010000010000000100010011;
ROM[31896] <= 32'b11111111110000010000000100010011;
ROM[31897] <= 32'b00000000000000010010001110000011;
ROM[31898] <= 32'b00000000011100100010010000100011;
ROM[31899] <= 32'b00000000100000100010001110000011;
ROM[31900] <= 32'b00000000011100010010000000100011;
ROM[31901] <= 32'b00000000010000010000000100010011;
ROM[31902] <= 32'b00000000010000100010001110000011;
ROM[31903] <= 32'b00000000011100010010000000100011;
ROM[31904] <= 32'b00000000010000010000000100010011;
ROM[31905] <= 32'b11111111110000010000000100010011;
ROM[31906] <= 32'b00000000000000010010001110000011;
ROM[31907] <= 32'b11111111110000010000000100010011;
ROM[31908] <= 32'b00000000000000010010010000000011;
ROM[31909] <= 32'b00000000011101000010001110110011;
ROM[31910] <= 32'b00000000011100010010000000100011;
ROM[31911] <= 32'b00000000010000010000000100010011;
ROM[31912] <= 32'b11111111110000010000000100010011;
ROM[31913] <= 32'b00000000000000010010001110000011;
ROM[31914] <= 32'b01000000011100000000001110110011;
ROM[31915] <= 32'b00000000000100111000001110010011;
ROM[31916] <= 32'b00000000011100010010000000100011;
ROM[31917] <= 32'b00000000010000010000000100010011;
ROM[31918] <= 32'b11111111110000010000000100010011;
ROM[31919] <= 32'b00000000000000010010001110000011;
ROM[31920] <= 32'b01000000011100000000001110110011;
ROM[31921] <= 32'b00000000000100111000001110010011;
ROM[31922] <= 32'b00000000011100010010000000100011;
ROM[31923] <= 32'b00000000010000010000000100010011;
ROM[31924] <= 32'b11111111110000010000000100010011;
ROM[31925] <= 32'b00000000000000010010001110000011;
ROM[31926] <= 32'b00000000000000111000101001100011;
ROM[31927] <= 32'b00000000000000011111001110110111;
ROM[31928] <= 32'b00111010000000111000001110010011;
ROM[31929] <= 32'b00000000111000111000001110110011;
ROM[31930] <= 32'b00000000000000111000000011100111;
ROM[31931] <= 32'b00000000000000100010001110000011;
ROM[31932] <= 32'b00000000011100010010000000100011;
ROM[31933] <= 32'b00000000010000010000000100010011;
ROM[31934] <= 32'b00000000010000100010001110000011;
ROM[31935] <= 32'b00000000011100010010000000100011;
ROM[31936] <= 32'b00000000010000010000000100010011;
ROM[31937] <= 32'b00000000000000011111001110110111;
ROM[31938] <= 32'b00110101000000111000001110010011;
ROM[31939] <= 32'b00000000111000111000001110110011;
ROM[31940] <= 32'b00000000011100010010000000100011;
ROM[31941] <= 32'b00000000010000010000000100010011;
ROM[31942] <= 32'b00000000001100010010000000100011;
ROM[31943] <= 32'b00000000010000010000000100010011;
ROM[31944] <= 32'b00000000010000010010000000100011;
ROM[31945] <= 32'b00000000010000010000000100010011;
ROM[31946] <= 32'b00000000010100010010000000100011;
ROM[31947] <= 32'b00000000010000010000000100010011;
ROM[31948] <= 32'b00000000011000010010000000100011;
ROM[31949] <= 32'b00000000010000010000000100010011;
ROM[31950] <= 32'b00000001010000000000001110010011;
ROM[31951] <= 32'b00000000100000111000001110010011;
ROM[31952] <= 32'b01000000011100010000001110110011;
ROM[31953] <= 32'b00000000011100000000001000110011;
ROM[31954] <= 32'b00000000001000000000000110110011;
ROM[31955] <= 32'b11010110000111111110000011101111;
ROM[31956] <= 32'b11111111110000010000000100010011;
ROM[31957] <= 32'b00000000000000010010001110000011;
ROM[31958] <= 32'b00000000011101100010000000100011;
ROM[31959] <= 32'b00000000010000100010001110000011;
ROM[31960] <= 32'b00000000011100010010000000100011;
ROM[31961] <= 32'b00000000010000010000000100010011;
ROM[31962] <= 32'b00000000000100000000001110010011;
ROM[31963] <= 32'b00000000011100010010000000100011;
ROM[31964] <= 32'b00000000010000010000000100010011;
ROM[31965] <= 32'b11111111110000010000000100010011;
ROM[31966] <= 32'b00000000000000010010001110000011;
ROM[31967] <= 32'b11111111110000010000000100010011;
ROM[31968] <= 32'b00000000000000010010010000000011;
ROM[31969] <= 32'b00000000011101000000001110110011;
ROM[31970] <= 32'b00000000011100010010000000100011;
ROM[31971] <= 32'b00000000010000010000000100010011;
ROM[31972] <= 32'b11111111110000010000000100010011;
ROM[31973] <= 32'b00000000000000010010001110000011;
ROM[31974] <= 32'b00000000011100100010001000100011;
ROM[31975] <= 32'b11101101000111111111000011101111;
ROM[31976] <= 32'b00000000000000000000001110010011;
ROM[31977] <= 32'b00000000011100010010000000100011;
ROM[31978] <= 32'b00000000010000010000000100010011;
ROM[31979] <= 32'b00000001010000000000001110010011;
ROM[31980] <= 32'b01000000011100011000001110110011;
ROM[31981] <= 32'b00000000000000111010000010000011;
ROM[31982] <= 32'b11111111110000010000000100010011;
ROM[31983] <= 32'b00000000000000010010001110000011;
ROM[31984] <= 32'b00000000011100100010000000100011;
ROM[31985] <= 32'b00000000010000100000000100010011;
ROM[31986] <= 32'b00000001010000000000001110010011;
ROM[31987] <= 32'b01000000011100011000001110110011;
ROM[31988] <= 32'b00000000010000111010000110000011;
ROM[31989] <= 32'b00000000100000111010001000000011;
ROM[31990] <= 32'b00000000110000111010001010000011;
ROM[31991] <= 32'b00000001000000111010001100000011;
ROM[31992] <= 32'b00000000000000001000000011100111;
ROM[31993] <= 32'b00000000010000100010001110000011;
ROM[31994] <= 32'b00000000011100010010000000100011;
ROM[31995] <= 32'b00000000010000010000000100010011;
ROM[31996] <= 32'b00000000110000100010001110000011;
ROM[31997] <= 32'b00000000011100010010000000100011;
ROM[31998] <= 32'b00000000010000010000000100010011;
ROM[31999] <= 32'b11111111110000010000000100010011;
ROM[32000] <= 32'b00000000000000010010001110000011;
ROM[32001] <= 32'b11111111110000010000000100010011;
ROM[32002] <= 32'b00000000000000010010010000000011;
ROM[32003] <= 32'b00000000100000111010001110110011;
ROM[32004] <= 32'b00000000011100010010000000100011;
ROM[32005] <= 32'b00000000010000010000000100010011;
ROM[32006] <= 32'b11111111110000010000000100010011;
ROM[32007] <= 32'b00000000000000010010001110000011;
ROM[32008] <= 32'b01000000011100000000001110110011;
ROM[32009] <= 32'b00000000000100111000001110010011;
ROM[32010] <= 32'b00000000011100010010000000100011;
ROM[32011] <= 32'b00000000010000010000000100010011;
ROM[32012] <= 32'b11111111110000010000000100010011;
ROM[32013] <= 32'b00000000000000010010001110000011;
ROM[32014] <= 32'b01000000011100000000001110110011;
ROM[32015] <= 32'b00000000000100111000001110010011;
ROM[32016] <= 32'b00000000011100010010000000100011;
ROM[32017] <= 32'b00000000010000010000000100010011;
ROM[32018] <= 32'b11111111110000010000000100010011;
ROM[32019] <= 32'b00000000000000010010001110000011;
ROM[32020] <= 32'b00000000000000111000101001100011;
ROM[32021] <= 32'b00000000000000011111001110110111;
ROM[32022] <= 32'b01010010010000111000001110010011;
ROM[32023] <= 32'b00000000111000111000001110110011;
ROM[32024] <= 32'b00000000000000111000000011100111;
ROM[32025] <= 32'b00000000000000100010001110000011;
ROM[32026] <= 32'b00000000011100010010000000100011;
ROM[32027] <= 32'b00000000010000010000000100010011;
ROM[32028] <= 32'b00000000100000100010001110000011;
ROM[32029] <= 32'b00000000011100010010000000100011;
ROM[32030] <= 32'b00000000010000010000000100010011;
ROM[32031] <= 32'b00000000010000100010001110000011;
ROM[32032] <= 32'b00000000011100010010000000100011;
ROM[32033] <= 32'b00000000010000010000000100010011;
ROM[32034] <= 32'b00000000000000011111001110110111;
ROM[32035] <= 32'b01001101010000111000001110010011;
ROM[32036] <= 32'b00000000111000111000001110110011;
ROM[32037] <= 32'b00000000011100010010000000100011;
ROM[32038] <= 32'b00000000010000010000000100010011;
ROM[32039] <= 32'b00000000001100010010000000100011;
ROM[32040] <= 32'b00000000010000010000000100010011;
ROM[32041] <= 32'b00000000010000010010000000100011;
ROM[32042] <= 32'b00000000010000010000000100010011;
ROM[32043] <= 32'b00000000010100010010000000100011;
ROM[32044] <= 32'b00000000010000010000000100010011;
ROM[32045] <= 32'b00000000011000010010000000100011;
ROM[32046] <= 32'b00000000010000010000000100010011;
ROM[32047] <= 32'b00000001010000000000001110010011;
ROM[32048] <= 32'b00000000110000111000001110010011;
ROM[32049] <= 32'b01000000011100010000001110110011;
ROM[32050] <= 32'b00000000011100000000001000110011;
ROM[32051] <= 32'b00000000001000000000000110110011;
ROM[32052] <= 32'b10101101110111111111000011101111;
ROM[32053] <= 32'b11111111110000010000000100010011;
ROM[32054] <= 32'b00000000000000010010001110000011;
ROM[32055] <= 32'b00000000011101100010000000100011;
ROM[32056] <= 32'b00000000010000100010001110000011;
ROM[32057] <= 32'b00000000011100010010000000100011;
ROM[32058] <= 32'b00000000010000010000000100010011;
ROM[32059] <= 32'b00000000000100000000001110010011;
ROM[32060] <= 32'b00000000011100010010000000100011;
ROM[32061] <= 32'b00000000010000010000000100010011;
ROM[32062] <= 32'b11111111110000010000000100010011;
ROM[32063] <= 32'b00000000000000010010001110000011;
ROM[32064] <= 32'b11111111110000010000000100010011;
ROM[32065] <= 32'b00000000000000010010010000000011;
ROM[32066] <= 32'b00000000011101000000001110110011;
ROM[32067] <= 32'b00000000011100010010000000100011;
ROM[32068] <= 32'b00000000010000010000000100010011;
ROM[32069] <= 32'b11111111110000010000000100010011;
ROM[32070] <= 32'b00000000000000010010001110000011;
ROM[32071] <= 32'b00000000011100100010001000100011;
ROM[32072] <= 32'b11101100010111111111000011101111;
ROM[32073] <= 32'b00000000000000000000001110010011;
ROM[32074] <= 32'b00000000011100010010000000100011;
ROM[32075] <= 32'b00000000010000010000000100010011;
ROM[32076] <= 32'b00000001010000000000001110010011;
ROM[32077] <= 32'b01000000011100011000001110110011;
ROM[32078] <= 32'b00000000000000111010000010000011;
ROM[32079] <= 32'b11111111110000010000000100010011;
ROM[32080] <= 32'b00000000000000010010001110000011;
ROM[32081] <= 32'b00000000011100100010000000100011;
ROM[32082] <= 32'b00000000010000100000000100010011;
ROM[32083] <= 32'b00000001010000000000001110010011;
ROM[32084] <= 32'b01000000011100011000001110110011;
ROM[32085] <= 32'b00000000010000111010000110000011;
ROM[32086] <= 32'b00000000100000111010001000000011;
ROM[32087] <= 32'b00000000110000111010001010000011;
ROM[32088] <= 32'b00000001000000111010001100000011;
ROM[32089] <= 32'b00000000000000001000000011100111;
ROM[32090] <= 32'b00000000000000010010000000100011;
ROM[32091] <= 32'b00000000010000010000000100010011;
ROM[32092] <= 32'b00000000000000010010000000100011;
ROM[32093] <= 32'b00000000010000010000000100010011;
ROM[32094] <= 32'b00000000000000010010000000100011;
ROM[32095] <= 32'b00000000010000010000000100010011;
ROM[32096] <= 32'b00000000100000100010001110000011;
ROM[32097] <= 32'b00000000011100010010000000100011;
ROM[32098] <= 32'b00000000010000010000000100010011;
ROM[32099] <= 32'b11111111110000010000000100010011;
ROM[32100] <= 32'b00000000000000010010001110000011;
ROM[32101] <= 32'b01000000011100000000001110110011;
ROM[32102] <= 32'b00000000011100010010000000100011;
ROM[32103] <= 32'b00000000010000010000000100010011;
ROM[32104] <= 32'b11111111110000010000000100010011;
ROM[32105] <= 32'b00000000000000010010001110000011;
ROM[32106] <= 32'b00000000011100011010001000100011;
ROM[32107] <= 32'b00000000100000100010001110000011;
ROM[32108] <= 32'b00000000011100010010000000100011;
ROM[32109] <= 32'b00000000010000010000000100010011;
ROM[32110] <= 32'b00000000100000100010001110000011;
ROM[32111] <= 32'b00000000011100010010000000100011;
ROM[32112] <= 32'b00000000010000010000000100010011;
ROM[32113] <= 32'b00000000000000011111001110110111;
ROM[32114] <= 32'b01100001000000111000001110010011;
ROM[32115] <= 32'b00000000111000111000001110110011;
ROM[32116] <= 32'b00000000011100010010000000100011;
ROM[32117] <= 32'b00000000010000010000000100010011;
ROM[32118] <= 32'b00000000001100010010000000100011;
ROM[32119] <= 32'b00000000010000010000000100010011;
ROM[32120] <= 32'b00000000010000010010000000100011;
ROM[32121] <= 32'b00000000010000010000000100010011;
ROM[32122] <= 32'b00000000010100010010000000100011;
ROM[32123] <= 32'b00000000010000010000000100010011;
ROM[32124] <= 32'b00000000011000010010000000100011;
ROM[32125] <= 32'b00000000010000010000000100010011;
ROM[32126] <= 32'b00000001010000000000001110010011;
ROM[32127] <= 32'b00000000100000111000001110010011;
ROM[32128] <= 32'b01000000011100010000001110110011;
ROM[32129] <= 32'b00000000011100000000001000110011;
ROM[32130] <= 32'b00000000001000000000000110110011;
ROM[32131] <= 32'b10100010000011110010000011101111;
ROM[32132] <= 32'b11111111110000010000000100010011;
ROM[32133] <= 32'b00000000000000010010001110000011;
ROM[32134] <= 32'b00000000011100011010010000100011;
ROM[32135] <= 32'b00000000010000011010001110000011;
ROM[32136] <= 32'b00000000011100010010000000100011;
ROM[32137] <= 32'b00000000010000010000000100010011;
ROM[32138] <= 32'b00000000100000100010001110000011;
ROM[32139] <= 32'b00000000011100010010000000100011;
ROM[32140] <= 32'b00000000010000010000000100010011;
ROM[32141] <= 32'b11111111110000010000000100010011;
ROM[32142] <= 32'b00000000000000010010001110000011;
ROM[32143] <= 32'b11111111110000010000000100010011;
ROM[32144] <= 32'b00000000000000010010010000000011;
ROM[32145] <= 32'b00000000100000111010001110110011;
ROM[32146] <= 32'b00000000011100010010000000100011;
ROM[32147] <= 32'b00000000010000010000000100010011;
ROM[32148] <= 32'b11111111110000010000000100010011;
ROM[32149] <= 32'b00000000000000010010001110000011;
ROM[32150] <= 32'b01000000011100000000001110110011;
ROM[32151] <= 32'b00000000000100111000001110010011;
ROM[32152] <= 32'b00000000011100010010000000100011;
ROM[32153] <= 32'b00000000010000010000000100010011;
ROM[32154] <= 32'b11111111110000010000000100010011;
ROM[32155] <= 32'b00000000000000010010001110000011;
ROM[32156] <= 32'b01000000011100000000001110110011;
ROM[32157] <= 32'b00000000000100111000001110010011;
ROM[32158] <= 32'b00000000011100010010000000100011;
ROM[32159] <= 32'b00000000010000010000000100010011;
ROM[32160] <= 32'b11111111110000010000000100010011;
ROM[32161] <= 32'b00000000000000010010001110000011;
ROM[32162] <= 32'b00000000000000111000101001100011;
ROM[32163] <= 32'b00000000000000100000001110110111;
ROM[32164] <= 32'b10001011100000111000001110010011;
ROM[32165] <= 32'b00000000111000111000001110110011;
ROM[32166] <= 32'b00000000000000111000000011100111;
ROM[32167] <= 32'b00000000100000011010001110000011;
ROM[32168] <= 32'b00000000011100010010000000100011;
ROM[32169] <= 32'b00000000010000010000000100010011;
ROM[32170] <= 32'b00000000010000011010001110000011;
ROM[32171] <= 32'b00000000011100010010000000100011;
ROM[32172] <= 32'b00000000010000010000000100010011;
ROM[32173] <= 32'b00000000010000011010001110000011;
ROM[32174] <= 32'b00000000011100010010000000100011;
ROM[32175] <= 32'b00000000010000010000000100010011;
ROM[32176] <= 32'b00000000000000011111001110110111;
ROM[32177] <= 32'b01110000110000111000001110010011;
ROM[32178] <= 32'b00000000111000111000001110110011;
ROM[32179] <= 32'b00000000011100010010000000100011;
ROM[32180] <= 32'b00000000010000010000000100010011;
ROM[32181] <= 32'b00000000001100010010000000100011;
ROM[32182] <= 32'b00000000010000010000000100010011;
ROM[32183] <= 32'b00000000010000010010000000100011;
ROM[32184] <= 32'b00000000010000010000000100010011;
ROM[32185] <= 32'b00000000010100010010000000100011;
ROM[32186] <= 32'b00000000010000010000000100010011;
ROM[32187] <= 32'b00000000011000010010000000100011;
ROM[32188] <= 32'b00000000010000010000000100010011;
ROM[32189] <= 32'b00000001010000000000001110010011;
ROM[32190] <= 32'b00000000100000111000001110010011;
ROM[32191] <= 32'b01000000011100010000001110110011;
ROM[32192] <= 32'b00000000011100000000001000110011;
ROM[32193] <= 32'b00000000001000000000000110110011;
ROM[32194] <= 32'b10010010010011110010000011101111;
ROM[32195] <= 32'b11111111110000010000000100010011;
ROM[32196] <= 32'b00000000000000010010001110000011;
ROM[32197] <= 32'b11111111110000010000000100010011;
ROM[32198] <= 32'b00000000000000010010010000000011;
ROM[32199] <= 32'b01000000011101000000001110110011;
ROM[32200] <= 32'b00000000011100010010000000100011;
ROM[32201] <= 32'b00000000010000010000000100010011;
ROM[32202] <= 32'b00000000000000011111001110110111;
ROM[32203] <= 32'b01110111010000111000001110010011;
ROM[32204] <= 32'b00000000111000111000001110110011;
ROM[32205] <= 32'b00000000011100010010000000100011;
ROM[32206] <= 32'b00000000010000010000000100010011;
ROM[32207] <= 32'b00000000001100010010000000100011;
ROM[32208] <= 32'b00000000010000010000000100010011;
ROM[32209] <= 32'b00000000010000010010000000100011;
ROM[32210] <= 32'b00000000010000010000000100010011;
ROM[32211] <= 32'b00000000010100010010000000100011;
ROM[32212] <= 32'b00000000010000010000000100010011;
ROM[32213] <= 32'b00000000011000010010000000100011;
ROM[32214] <= 32'b00000000010000010000000100010011;
ROM[32215] <= 32'b00000001010000000000001110010011;
ROM[32216] <= 32'b00000000010000111000001110010011;
ROM[32217] <= 32'b01000000011100010000001110110011;
ROM[32218] <= 32'b00000000011100000000001000110011;
ROM[32219] <= 32'b00000000001000000000000110110011;
ROM[32220] <= 32'b10001011010111110010000011101111;
ROM[32221] <= 32'b11111111110000010000000100010011;
ROM[32222] <= 32'b00000000000000010010001110000011;
ROM[32223] <= 32'b00000000011100011010000000100011;
ROM[32224] <= 32'b00000000000000100010001110000011;
ROM[32225] <= 32'b00000000011100010010000000100011;
ROM[32226] <= 32'b00000000010000010000000100010011;
ROM[32227] <= 32'b00000000000000011010001110000011;
ROM[32228] <= 32'b00000000011100010010000000100011;
ROM[32229] <= 32'b00000000010000010000000100010011;
ROM[32230] <= 32'b11111111110000010000000100010011;
ROM[32231] <= 32'b00000000000000010010001110000011;
ROM[32232] <= 32'b11111111110000010000000100010011;
ROM[32233] <= 32'b00000000000000010010010000000011;
ROM[32234] <= 32'b01000000011101000000001110110011;
ROM[32235] <= 32'b00000000011100010010000000100011;
ROM[32236] <= 32'b00000000010000010000000100010011;
ROM[32237] <= 32'b00000000000000100010001110000011;
ROM[32238] <= 32'b00000000011100010010000000100011;
ROM[32239] <= 32'b00000000010000010000000100010011;
ROM[32240] <= 32'b00000000000000011010001110000011;
ROM[32241] <= 32'b00000000011100010010000000100011;
ROM[32242] <= 32'b00000000010000010000000100010011;
ROM[32243] <= 32'b11111111110000010000000100010011;
ROM[32244] <= 32'b00000000000000010010001110000011;
ROM[32245] <= 32'b11111111110000010000000100010011;
ROM[32246] <= 32'b00000000000000010010010000000011;
ROM[32247] <= 32'b00000000011101000000001110110011;
ROM[32248] <= 32'b00000000011100010010000000100011;
ROM[32249] <= 32'b00000000010000010000000100010011;
ROM[32250] <= 32'b00000000010000100010001110000011;
ROM[32251] <= 32'b00000000011100010010000000100011;
ROM[32252] <= 32'b00000000010000010000000100010011;
ROM[32253] <= 32'b00000000010000011010001110000011;
ROM[32254] <= 32'b00000000011100010010000000100011;
ROM[32255] <= 32'b00000000010000010000000100010011;
ROM[32256] <= 32'b11111111110000010000000100010011;
ROM[32257] <= 32'b00000000000000010010001110000011;
ROM[32258] <= 32'b11111111110000010000000100010011;
ROM[32259] <= 32'b00000000000000010010010000000011;
ROM[32260] <= 32'b00000000011101000000001110110011;
ROM[32261] <= 32'b00000000011100010010000000100011;
ROM[32262] <= 32'b00000000010000010000000100010011;
ROM[32263] <= 32'b00000000000000100000001110110111;
ROM[32264] <= 32'b10000110100000111000001110010011;
ROM[32265] <= 32'b00000000111000111000001110110011;
ROM[32266] <= 32'b00000000011100010010000000100011;
ROM[32267] <= 32'b00000000010000010000000100010011;
ROM[32268] <= 32'b00000000001100010010000000100011;
ROM[32269] <= 32'b00000000010000010000000100010011;
ROM[32270] <= 32'b00000000010000010010000000100011;
ROM[32271] <= 32'b00000000010000010000000100010011;
ROM[32272] <= 32'b00000000010100010010000000100011;
ROM[32273] <= 32'b00000000010000010000000100010011;
ROM[32274] <= 32'b00000000011000010010000000100011;
ROM[32275] <= 32'b00000000010000010000000100010011;
ROM[32276] <= 32'b00000001010000000000001110010011;
ROM[32277] <= 32'b00000000110000111000001110010011;
ROM[32278] <= 32'b01000000011100010000001110110011;
ROM[32279] <= 32'b00000000011100000000001000110011;
ROM[32280] <= 32'b00000000001000000000000110110011;
ROM[32281] <= 32'b11110100100011111111000011101111;
ROM[32282] <= 32'b11111111110000010000000100010011;
ROM[32283] <= 32'b00000000000000010010001110000011;
ROM[32284] <= 32'b00000000011101100010000000100011;
ROM[32285] <= 32'b00000000010000011010001110000011;
ROM[32286] <= 32'b00000000011100010010000000100011;
ROM[32287] <= 32'b00000000010000010000000100010011;
ROM[32288] <= 32'b00000000000100000000001110010011;
ROM[32289] <= 32'b00000000011100010010000000100011;
ROM[32290] <= 32'b00000000010000010000000100010011;
ROM[32291] <= 32'b11111111110000010000000100010011;
ROM[32292] <= 32'b00000000000000010010001110000011;
ROM[32293] <= 32'b11111111110000010000000100010011;
ROM[32294] <= 32'b00000000000000010010010000000011;
ROM[32295] <= 32'b00000000011101000000001110110011;
ROM[32296] <= 32'b00000000011100010010000000100011;
ROM[32297] <= 32'b00000000010000010000000100010011;
ROM[32298] <= 32'b11111111110000010000000100010011;
ROM[32299] <= 32'b00000000000000010010001110000011;
ROM[32300] <= 32'b00000000011100011010001000100011;
ROM[32301] <= 32'b11010110100111111111000011101111;
ROM[32302] <= 32'b00000000000000000000001110010011;
ROM[32303] <= 32'b00000000011100010010000000100011;
ROM[32304] <= 32'b00000000010000010000000100010011;
ROM[32305] <= 32'b00000001010000000000001110010011;
ROM[32306] <= 32'b01000000011100011000001110110011;
ROM[32307] <= 32'b00000000000000111010000010000011;
ROM[32308] <= 32'b11111111110000010000000100010011;
ROM[32309] <= 32'b00000000000000010010001110000011;
ROM[32310] <= 32'b00000000011100100010000000100011;
ROM[32311] <= 32'b00000000010000100000000100010011;
ROM[32312] <= 32'b00000001010000000000001110010011;
ROM[32313] <= 32'b01000000011100011000001110110011;
ROM[32314] <= 32'b00000000010000111010000110000011;
ROM[32315] <= 32'b00000000100000111010001000000011;
ROM[32316] <= 32'b00000000110000111010001010000011;
ROM[32317] <= 32'b00000001000000111010001100000011;
ROM[32318] <= 32'b00000000000000001000000011100111;
ROM[32319] <= 32'b00000000000000010010000000100011;
ROM[32320] <= 32'b00000000010000010000000100010011;
ROM[32321] <= 32'b00000000101100000000001110010011;
ROM[32322] <= 32'b00000000011100010010000000100011;
ROM[32323] <= 32'b00000000010000010000000100010011;
ROM[32324] <= 32'b00000000000000100000001110110111;
ROM[32325] <= 32'b10010101110000111000001110010011;
ROM[32326] <= 32'b00000000111000111000001110110011;
ROM[32327] <= 32'b00000000011100010010000000100011;
ROM[32328] <= 32'b00000000010000010000000100010011;
ROM[32329] <= 32'b00000000001100010010000000100011;
ROM[32330] <= 32'b00000000010000010000000100010011;
ROM[32331] <= 32'b00000000010000010010000000100011;
ROM[32332] <= 32'b00000000010000010000000100010011;
ROM[32333] <= 32'b00000000010100010010000000100011;
ROM[32334] <= 32'b00000000010000010000000100010011;
ROM[32335] <= 32'b00000000011000010010000000100011;
ROM[32336] <= 32'b00000000010000010000000100010011;
ROM[32337] <= 32'b00000001010000000000001110010011;
ROM[32338] <= 32'b00000000010000111000001110010011;
ROM[32339] <= 32'b01000000011100010000001110110011;
ROM[32340] <= 32'b00000000011100000000001000110011;
ROM[32341] <= 32'b00000000001000000000000110110011;
ROM[32342] <= 32'b11010111110111110100000011101111;
ROM[32343] <= 32'b11111111110000010000000100010011;
ROM[32344] <= 32'b00000000000000010010001110000011;
ROM[32345] <= 32'b00000000000000111000001010010011;
ROM[32346] <= 32'b00000000000000100010001110000011;
ROM[32347] <= 32'b00000000011100010010000000100011;
ROM[32348] <= 32'b00000000010000010000000100010011;
ROM[32349] <= 32'b11111111110000010000000100010011;
ROM[32350] <= 32'b00000000000000010010001110000011;
ROM[32351] <= 32'b00000000110100101000010000110011;
ROM[32352] <= 32'b00000000011101000010000000100011;
ROM[32353] <= 32'b00000000010000100010001110000011;
ROM[32354] <= 32'b00000000011100010010000000100011;
ROM[32355] <= 32'b00000000010000010000000100010011;
ROM[32356] <= 32'b00000000110000100010001110000011;
ROM[32357] <= 32'b00000000011100010010000000100011;
ROM[32358] <= 32'b00000000010000010000000100010011;
ROM[32359] <= 32'b11111111110000010000000100010011;
ROM[32360] <= 32'b00000000000000010010001110000011;
ROM[32361] <= 32'b11111111110000010000000100010011;
ROM[32362] <= 32'b00000000000000010010010000000011;
ROM[32363] <= 32'b01000000011101000000001110110011;
ROM[32364] <= 32'b00000000011100010010000000100011;
ROM[32365] <= 32'b00000000010000010000000100010011;
ROM[32366] <= 32'b11111111110000010000000100010011;
ROM[32367] <= 32'b00000000000000010010001110000011;
ROM[32368] <= 32'b00000000110100101000010000110011;
ROM[32369] <= 32'b00000000011101000010001000100011;
ROM[32370] <= 32'b00000000100000100010001110000011;
ROM[32371] <= 32'b00000000011100010010000000100011;
ROM[32372] <= 32'b00000000010000010000000100010011;
ROM[32373] <= 32'b11111111110000010000000100010011;
ROM[32374] <= 32'b00000000000000010010001110000011;
ROM[32375] <= 32'b00000000110100101000010000110011;
ROM[32376] <= 32'b00000000011101000010010000100011;
ROM[32377] <= 32'b00000000110000100010001110000011;
ROM[32378] <= 32'b00000000011100010010000000100011;
ROM[32379] <= 32'b00000000010000010000000100010011;
ROM[32380] <= 32'b11111111110000010000000100010011;
ROM[32381] <= 32'b00000000000000010010001110000011;
ROM[32382] <= 32'b00000000110100101000010000110011;
ROM[32383] <= 32'b00000000011101000010011000100011;
ROM[32384] <= 32'b00000001000000100010001110000011;
ROM[32385] <= 32'b00000000011100010010000000100011;
ROM[32386] <= 32'b00000000010000010000000100010011;
ROM[32387] <= 32'b11111111110000010000000100010011;
ROM[32388] <= 32'b00000000000000010010001110000011;
ROM[32389] <= 32'b00000000110100101000010000110011;
ROM[32390] <= 32'b00000000011101000010100000100011;
ROM[32391] <= 32'b00000000000000000000001110010011;
ROM[32392] <= 32'b00000000011100010010000000100011;
ROM[32393] <= 32'b00000000010000010000000100010011;
ROM[32394] <= 32'b11111111110000010000000100010011;
ROM[32395] <= 32'b00000000000000010010001110000011;
ROM[32396] <= 32'b00000000110100101000010000110011;
ROM[32397] <= 32'b00000000011101000010101000100011;
ROM[32398] <= 32'b00000000010000000000001110010011;
ROM[32399] <= 32'b00000000011100010010000000100011;
ROM[32400] <= 32'b00000000010000010000000100010011;
ROM[32401] <= 32'b11111111110000010000000100010011;
ROM[32402] <= 32'b00000000000000010010001110000011;
ROM[32403] <= 32'b00000000110100101000010000110011;
ROM[32404] <= 32'b00000000011101000010110000100011;
ROM[32405] <= 32'b00000000010000000000001110010011;
ROM[32406] <= 32'b00000000011100010010000000100011;
ROM[32407] <= 32'b00000000010000010000000100010011;
ROM[32408] <= 32'b11111111110000010000000100010011;
ROM[32409] <= 32'b00000000000000010010001110000011;
ROM[32410] <= 32'b00000000110100101000010000110011;
ROM[32411] <= 32'b00000000011101000010111000100011;
ROM[32412] <= 32'b00100000000000000000001110010011;
ROM[32413] <= 32'b00000000011100010010000000100011;
ROM[32414] <= 32'b00000000010000010000000100010011;
ROM[32415] <= 32'b11111111110000010000000100010011;
ROM[32416] <= 32'b00000000000000010010001110000011;
ROM[32417] <= 32'b00000000110100101000010000110011;
ROM[32418] <= 32'b00000010011101000010010000100011;
ROM[32419] <= 32'b00000000110100101000010000110011;
ROM[32420] <= 32'b00000010100001000010001110000011;
ROM[32421] <= 32'b00000000011100010010000000100011;
ROM[32422] <= 32'b00000000010000010000000100010011;
ROM[32423] <= 32'b00000000000000100000001110110111;
ROM[32424] <= 32'b10101110100000111000001110010011;
ROM[32425] <= 32'b00000000111000111000001110110011;
ROM[32426] <= 32'b00000000011100010010000000100011;
ROM[32427] <= 32'b00000000010000010000000100010011;
ROM[32428] <= 32'b00000000001100010010000000100011;
ROM[32429] <= 32'b00000000010000010000000100010011;
ROM[32430] <= 32'b00000000010000010010000000100011;
ROM[32431] <= 32'b00000000010000010000000100010011;
ROM[32432] <= 32'b00000000010100010010000000100011;
ROM[32433] <= 32'b00000000010000010000000100010011;
ROM[32434] <= 32'b00000000011000010010000000100011;
ROM[32435] <= 32'b00000000010000010000000100010011;
ROM[32436] <= 32'b00000001010000000000001110010011;
ROM[32437] <= 32'b00000000010000111000001110010011;
ROM[32438] <= 32'b01000000011100010000001110110011;
ROM[32439] <= 32'b00000000011100000000001000110011;
ROM[32440] <= 32'b00000000001000000000000110110011;
ROM[32441] <= 32'b11011001110011100000000011101111;
ROM[32442] <= 32'b11111111110000010000000100010011;
ROM[32443] <= 32'b00000000000000010010001110000011;
ROM[32444] <= 32'b00000000110100101000010000110011;
ROM[32445] <= 32'b00000010011101000010000000100011;
ROM[32446] <= 32'b00000000110100101000010000110011;
ROM[32447] <= 32'b00000010100001000010001110000011;
ROM[32448] <= 32'b00000000011100010010000000100011;
ROM[32449] <= 32'b00000000010000010000000100010011;
ROM[32450] <= 32'b00000000000000100000001110110111;
ROM[32451] <= 32'b10110101010000111000001110010011;
ROM[32452] <= 32'b00000000111000111000001110110011;
ROM[32453] <= 32'b00000000011100010010000000100011;
ROM[32454] <= 32'b00000000010000010000000100010011;
ROM[32455] <= 32'b00000000001100010010000000100011;
ROM[32456] <= 32'b00000000010000010000000100010011;
ROM[32457] <= 32'b00000000010000010010000000100011;
ROM[32458] <= 32'b00000000010000010000000100010011;
ROM[32459] <= 32'b00000000010100010010000000100011;
ROM[32460] <= 32'b00000000010000010000000100010011;
ROM[32461] <= 32'b00000000011000010010000000100011;
ROM[32462] <= 32'b00000000010000010000000100010011;
ROM[32463] <= 32'b00000001010000000000001110010011;
ROM[32464] <= 32'b00000000010000111000001110010011;
ROM[32465] <= 32'b01000000011100010000001110110011;
ROM[32466] <= 32'b00000000011100000000001000110011;
ROM[32467] <= 32'b00000000001000000000000110110011;
ROM[32468] <= 32'b11010011000011100000000011101111;
ROM[32469] <= 32'b11111111110000010000000100010011;
ROM[32470] <= 32'b00000000000000010010001110000011;
ROM[32471] <= 32'b00000000110100101000010000110011;
ROM[32472] <= 32'b00000010011101000010001000100011;
ROM[32473] <= 32'b00000000000000000000001110010011;
ROM[32474] <= 32'b00000000011100010010000000100011;
ROM[32475] <= 32'b00000000010000010000000100010011;
ROM[32476] <= 32'b11111111110000010000000100010011;
ROM[32477] <= 32'b00000000000000010010001110000011;
ROM[32478] <= 32'b00000000011100011010000000100011;
ROM[32479] <= 32'b00000000000000011010001110000011;
ROM[32480] <= 32'b00000000011100010010000000100011;
ROM[32481] <= 32'b00000000010000010000000100010011;
ROM[32482] <= 32'b00000000110100101000010000110011;
ROM[32483] <= 32'b00000000110001000010001110000011;
ROM[32484] <= 32'b00000000011100010010000000100011;
ROM[32485] <= 32'b00000000010000010000000100010011;
ROM[32486] <= 32'b11111111110000010000000100010011;
ROM[32487] <= 32'b00000000000000010010001110000011;
ROM[32488] <= 32'b11111111110000010000000100010011;
ROM[32489] <= 32'b00000000000000010010010000000011;
ROM[32490] <= 32'b00000000011101000010001110110011;
ROM[32491] <= 32'b00000000011100010010000000100011;
ROM[32492] <= 32'b00000000010000010000000100010011;
ROM[32493] <= 32'b11111111110000010000000100010011;
ROM[32494] <= 32'b00000000000000010010001110000011;
ROM[32495] <= 32'b01000000011100000000001110110011;
ROM[32496] <= 32'b00000000000100111000001110010011;
ROM[32497] <= 32'b00000000011100010010000000100011;
ROM[32498] <= 32'b00000000010000010000000100010011;
ROM[32499] <= 32'b11111111110000010000000100010011;
ROM[32500] <= 32'b00000000000000010010001110000011;
ROM[32501] <= 32'b00000000000000111000101001100011;
ROM[32502] <= 32'b00000000000000100000001110110111;
ROM[32503] <= 32'b11011001100000111000001110010011;
ROM[32504] <= 32'b00000000111000111000001110110011;
ROM[32505] <= 32'b00000000000000111000000011100111;
ROM[32506] <= 32'b00000000110100101000010000110011;
ROM[32507] <= 32'b00000000010001000010001110000011;
ROM[32508] <= 32'b00000000011100010010000000100011;
ROM[32509] <= 32'b00000000010000010000000100010011;
ROM[32510] <= 32'b00000000000100000000001110010011;
ROM[32511] <= 32'b00000000011100010010000000100011;
ROM[32512] <= 32'b00000000010000010000000100010011;
ROM[32513] <= 32'b11111111110000010000000100010011;
ROM[32514] <= 32'b00000000000000010010001110000011;
ROM[32515] <= 32'b11111111110000010000000100010011;
ROM[32516] <= 32'b00000000000000010010010000000011;
ROM[32517] <= 32'b00000000011101000000001110110011;
ROM[32518] <= 32'b00000000011100010010000000100011;
ROM[32519] <= 32'b00000000010000010000000100010011;
ROM[32520] <= 32'b11111111110000010000000100010011;
ROM[32521] <= 32'b00000000000000010010001110000011;
ROM[32522] <= 32'b00000000110100101000010000110011;
ROM[32523] <= 32'b00000000011101000010001000100011;
ROM[32524] <= 32'b00000000010100010010000000100011;
ROM[32525] <= 32'b00000000010000010000000100010011;
ROM[32526] <= 32'b00000000110100101000010000110011;
ROM[32527] <= 32'b00000000000001000010001110000011;
ROM[32528] <= 32'b00000000011100010010000000100011;
ROM[32529] <= 32'b00000000010000010000000100010011;
ROM[32530] <= 32'b00000000000000100000001110110111;
ROM[32531] <= 32'b11001001010000111000001110010011;
ROM[32532] <= 32'b00000000111000111000001110110011;
ROM[32533] <= 32'b00000000011100010010000000100011;
ROM[32534] <= 32'b00000000010000010000000100010011;
ROM[32535] <= 32'b00000000001100010010000000100011;
ROM[32536] <= 32'b00000000010000010000000100010011;
ROM[32537] <= 32'b00000000010000010010000000100011;
ROM[32538] <= 32'b00000000010000010000000100010011;
ROM[32539] <= 32'b00000000010100010010000000100011;
ROM[32540] <= 32'b00000000010000010000000100010011;
ROM[32541] <= 32'b00000000011000010010000000100011;
ROM[32542] <= 32'b00000000010000010000000100010011;
ROM[32543] <= 32'b00000001010000000000001110010011;
ROM[32544] <= 32'b00000000010000111000001110010011;
ROM[32545] <= 32'b01000000011100010000001110110011;
ROM[32546] <= 32'b00000000011100000000001000110011;
ROM[32547] <= 32'b00000000001000000000000110110011;
ROM[32548] <= 32'b01101001010100000011000011101111;
ROM[32549] <= 32'b00000000000000100000001110110111;
ROM[32550] <= 32'b11001110000000111000001110010011;
ROM[32551] <= 32'b00000000111000111000001110110011;
ROM[32552] <= 32'b00000000011100010010000000100011;
ROM[32553] <= 32'b00000000010000010000000100010011;
ROM[32554] <= 32'b00000000001100010010000000100011;
ROM[32555] <= 32'b00000000010000010000000100010011;
ROM[32556] <= 32'b00000000010000010010000000100011;
ROM[32557] <= 32'b00000000010000010000000100010011;
ROM[32558] <= 32'b00000000010100010010000000100011;
ROM[32559] <= 32'b00000000010000010000000100010011;
ROM[32560] <= 32'b00000000011000010010000000100011;
ROM[32561] <= 32'b00000000010000010000000100010011;
ROM[32562] <= 32'b00000001010000000000001110010011;
ROM[32563] <= 32'b00000000100000111000001110010011;
ROM[32564] <= 32'b01000000011100010000001110110011;
ROM[32565] <= 32'b00000000011100000000001000110011;
ROM[32566] <= 32'b00000000001000000000000110110011;
ROM[32567] <= 32'b01011101010000000001000011101111;
ROM[32568] <= 32'b11111111110000010000000100010011;
ROM[32569] <= 32'b00000000000000010010001110000011;
ROM[32570] <= 32'b00000000011101100010000000100011;
ROM[32571] <= 32'b00000000000000011010001110000011;
ROM[32572] <= 32'b00000000011100010010000000100011;
ROM[32573] <= 32'b00000000010000010000000100010011;
ROM[32574] <= 32'b00000000000100000000001110010011;
ROM[32575] <= 32'b00000000011100010010000000100011;
ROM[32576] <= 32'b00000000010000010000000100010011;
ROM[32577] <= 32'b11111111110000010000000100010011;
ROM[32578] <= 32'b00000000000000010010001110000011;
ROM[32579] <= 32'b11111111110000010000000100010011;
ROM[32580] <= 32'b00000000000000010010010000000011;
ROM[32581] <= 32'b00000000011101000000001110110011;
ROM[32582] <= 32'b00000000011100010010000000100011;
ROM[32583] <= 32'b00000000010000010000000100010011;
ROM[32584] <= 32'b11111111110000010000000100010011;
ROM[32585] <= 32'b00000000000000010010001110000011;
ROM[32586] <= 32'b00000000011100011010000000100011;
ROM[32587] <= 32'b00000000110100101000010000110011;
ROM[32588] <= 32'b00000000000001000010001110000011;
ROM[32589] <= 32'b00000000011100010010000000100011;
ROM[32590] <= 32'b00000000010000010000000100010011;
ROM[32591] <= 32'b00000000000000100000001110110111;
ROM[32592] <= 32'b11011000100000111000001110010011;
ROM[32593] <= 32'b00000000111000111000001110110011;
ROM[32594] <= 32'b00000000011100010010000000100011;
ROM[32595] <= 32'b00000000010000010000000100010011;
ROM[32596] <= 32'b00000000001100010010000000100011;
ROM[32597] <= 32'b00000000010000010000000100010011;
ROM[32598] <= 32'b00000000010000010010000000100011;
ROM[32599] <= 32'b00000000010000010000000100010011;
ROM[32600] <= 32'b00000000010100010010000000100011;
ROM[32601] <= 32'b00000000010000010000000100010011;
ROM[32602] <= 32'b00000000011000010010000000100011;
ROM[32603] <= 32'b00000000010000010000000100010011;
ROM[32604] <= 32'b00000001010000000000001110010011;
ROM[32605] <= 32'b00000000010000111000001110010011;
ROM[32606] <= 32'b01000000011100010000001110110011;
ROM[32607] <= 32'b00000000011100000000001000110011;
ROM[32608] <= 32'b00000000001000000000000110110011;
ROM[32609] <= 32'b01000011100100000011000011101111;
ROM[32610] <= 32'b11111111110000010000000100010011;
ROM[32611] <= 32'b00000000000000010010001110000011;
ROM[32612] <= 32'b00000000011101100010000000100011;
ROM[32613] <= 32'b11011110100111111111000011101111;
ROM[32614] <= 32'b00000000010100010010000000100011;
ROM[32615] <= 32'b00000000010000010000000100010011;
ROM[32616] <= 32'b00000001010000000000001110010011;
ROM[32617] <= 32'b01000000011100011000001110110011;
ROM[32618] <= 32'b00000000000000111010000010000011;
ROM[32619] <= 32'b11111111110000010000000100010011;
ROM[32620] <= 32'b00000000000000010010001110000011;
ROM[32621] <= 32'b00000000011100100010000000100011;
ROM[32622] <= 32'b00000000010000100000000100010011;
ROM[32623] <= 32'b00000001010000000000001110010011;
ROM[32624] <= 32'b01000000011100011000001110110011;
ROM[32625] <= 32'b00000000010000111010000110000011;
ROM[32626] <= 32'b00000000100000111010001000000011;
ROM[32627] <= 32'b00000000110000111010001010000011;
ROM[32628] <= 32'b00000001000000111010001100000011;
ROM[32629] <= 32'b00000000000000001000000011100111;
ROM[32630] <= 32'b00000000000000100010001110000011;
ROM[32631] <= 32'b00000000011100010010000000100011;
ROM[32632] <= 32'b00000000010000010000000100010011;
ROM[32633] <= 32'b11111111110000010000000100010011;
ROM[32634] <= 32'b00000000000000010010001110000011;
ROM[32635] <= 32'b00000000000000111000001010010011;
ROM[32636] <= 32'b00000000110100101000010000110011;
ROM[32637] <= 32'b00000010000001000010001110000011;
ROM[32638] <= 32'b00000000011100010010000000100011;
ROM[32639] <= 32'b00000000010000010000000100010011;
ROM[32640] <= 32'b00000000000000100000001110110111;
ROM[32641] <= 32'b11100100110000111000001110010011;
ROM[32642] <= 32'b00000000111000111000001110110011;
ROM[32643] <= 32'b00000000011100010010000000100011;
ROM[32644] <= 32'b00000000010000010000000100010011;
ROM[32645] <= 32'b00000000001100010010000000100011;
ROM[32646] <= 32'b00000000010000010000000100010011;
ROM[32647] <= 32'b00000000010000010010000000100011;
ROM[32648] <= 32'b00000000010000010000000100010011;
ROM[32649] <= 32'b00000000010100010010000000100011;
ROM[32650] <= 32'b00000000010000010000000100010011;
ROM[32651] <= 32'b00000000011000010010000000100011;
ROM[32652] <= 32'b00000000010000010000000100010011;
ROM[32653] <= 32'b00000001010000000000001110010011;
ROM[32654] <= 32'b00000000010000111000001110010011;
ROM[32655] <= 32'b01000000011100010000001110110011;
ROM[32656] <= 32'b00000000011100000000001000110011;
ROM[32657] <= 32'b00000000001000000000000110110011;
ROM[32658] <= 32'b10101100100011100000000011101111;
ROM[32659] <= 32'b11111111110000010000000100010011;
ROM[32660] <= 32'b00000000000000010010001110000011;
ROM[32661] <= 32'b00000000011101100010000000100011;
ROM[32662] <= 32'b00000000110100101000010000110011;
ROM[32663] <= 32'b00000010010001000010001110000011;
ROM[32664] <= 32'b00000000011100010010000000100011;
ROM[32665] <= 32'b00000000010000010000000100010011;
ROM[32666] <= 32'b00000000000000100000001110110111;
ROM[32667] <= 32'b11101011010000111000001110010011;
ROM[32668] <= 32'b00000000111000111000001110110011;
ROM[32669] <= 32'b00000000011100010010000000100011;
ROM[32670] <= 32'b00000000010000010000000100010011;
ROM[32671] <= 32'b00000000001100010010000000100011;
ROM[32672] <= 32'b00000000010000010000000100010011;
ROM[32673] <= 32'b00000000010000010010000000100011;
ROM[32674] <= 32'b00000000010000010000000100010011;
ROM[32675] <= 32'b00000000010100010010000000100011;
ROM[32676] <= 32'b00000000010000010000000100010011;
ROM[32677] <= 32'b00000000011000010010000000100011;
ROM[32678] <= 32'b00000000010000010000000100010011;
ROM[32679] <= 32'b00000001010000000000001110010011;
ROM[32680] <= 32'b00000000010000111000001110010011;
ROM[32681] <= 32'b01000000011100010000001110110011;
ROM[32682] <= 32'b00000000011100000000001000110011;
ROM[32683] <= 32'b00000000001000000000000110110011;
ROM[32684] <= 32'b10100110000011100000000011101111;
ROM[32685] <= 32'b11111111110000010000000100010011;
ROM[32686] <= 32'b00000000000000010010001110000011;
ROM[32687] <= 32'b00000000011101100010000000100011;
ROM[32688] <= 32'b00000000010100010010000000100011;
ROM[32689] <= 32'b00000000010000010000000100010011;
ROM[32690] <= 32'b00000000000000100000001110110111;
ROM[32691] <= 32'b11110001010000111000001110010011;
ROM[32692] <= 32'b00000000111000111000001110110011;
ROM[32693] <= 32'b00000000011100010010000000100011;
ROM[32694] <= 32'b00000000010000010000000100010011;
ROM[32695] <= 32'b00000000001100010010000000100011;
ROM[32696] <= 32'b00000000010000010000000100010011;
ROM[32697] <= 32'b00000000010000010010000000100011;
ROM[32698] <= 32'b00000000010000010000000100010011;
ROM[32699] <= 32'b00000000010100010010000000100011;
ROM[32700] <= 32'b00000000010000010000000100010011;
ROM[32701] <= 32'b00000000011000010010000000100011;
ROM[32702] <= 32'b00000000010000010000000100010011;
ROM[32703] <= 32'b00000001010000000000001110010011;
ROM[32704] <= 32'b00000000010000111000001110010011;
ROM[32705] <= 32'b01000000011100010000001110110011;
ROM[32706] <= 32'b00000000011100000000001000110011;
ROM[32707] <= 32'b00000000001000000000000110110011;
ROM[32708] <= 32'b11000100110111110011000011101111;
ROM[32709] <= 32'b11111111110000010000000100010011;
ROM[32710] <= 32'b00000000000000010010001110000011;
ROM[32711] <= 32'b00000000011101100010000000100011;
ROM[32712] <= 32'b00000000000000000000001110010011;
ROM[32713] <= 32'b00000000011100010010000000100011;
ROM[32714] <= 32'b00000000010000010000000100010011;
ROM[32715] <= 32'b00000001010000000000001110010011;
ROM[32716] <= 32'b01000000011100011000001110110011;
ROM[32717] <= 32'b00000000000000111010000010000011;
ROM[32718] <= 32'b11111111110000010000000100010011;
ROM[32719] <= 32'b00000000000000010010001110000011;
ROM[32720] <= 32'b00000000011100100010000000100011;
ROM[32721] <= 32'b00000000010000100000000100010011;
ROM[32722] <= 32'b00000001010000000000001110010011;
ROM[32723] <= 32'b01000000011100011000001110110011;
ROM[32724] <= 32'b00000000010000111010000110000011;
ROM[32725] <= 32'b00000000100000111010001000000011;
ROM[32726] <= 32'b00000000110000111010001010000011;
ROM[32727] <= 32'b00000001000000111010001100000011;
ROM[32728] <= 32'b00000000000000001000000011100111;
ROM[32729] <= 32'b00000000000000100010001110000011;
ROM[32730] <= 32'b00000000011100010010000000100011;
ROM[32731] <= 32'b00000000010000010000000100010011;
ROM[32732] <= 32'b11111111110000010000000100010011;
ROM[32733] <= 32'b00000000000000010010001110000011;
ROM[32734] <= 32'b00000000000000111000001010010011;
ROM[32735] <= 32'b00000000110100101000010000110011;
ROM[32736] <= 32'b00000000000001000010001110000011;
ROM[32737] <= 32'b00000000011100010010000000100011;
ROM[32738] <= 32'b00000000010000010000000100010011;
ROM[32739] <= 32'b00000000000000100000001110110111;
ROM[32740] <= 32'b11111101100000111000001110010011;
ROM[32741] <= 32'b00000000111000111000001110110011;
ROM[32742] <= 32'b00000000011100010010000000100011;
ROM[32743] <= 32'b00000000010000010000000100010011;
ROM[32744] <= 32'b00000000001100010010000000100011;
ROM[32745] <= 32'b00000000010000010000000100010011;
ROM[32746] <= 32'b00000000010000010010000000100011;
ROM[32747] <= 32'b00000000010000010000000100010011;
ROM[32748] <= 32'b00000000010100010010000000100011;
ROM[32749] <= 32'b00000000010000010000000100010011;
ROM[32750] <= 32'b00000000011000010010000000100011;
ROM[32751] <= 32'b00000000010000010000000100010011;
ROM[32752] <= 32'b00000001010000000000001110010011;
ROM[32753] <= 32'b00000000010000111000001110010011;
ROM[32754] <= 32'b01000000011100010000001110110011;
ROM[32755] <= 32'b00000000011100000000001000110011;
ROM[32756] <= 32'b00000000001000000000000110110011;
ROM[32757] <= 32'b00110101000100000011000011101111;
ROM[32758] <= 32'b00000000110100101000010000110011;
ROM[32759] <= 32'b00000010100001000010001110000011;
ROM[32760] <= 32'b00000000011100010010000000100011;
ROM[32761] <= 32'b00000000010000010000000100010011;
ROM[32762] <= 32'b11111111110000010000000100010011;
ROM[32763] <= 32'b00000000000000010010001110000011;
ROM[32764] <= 32'b11111111110000010000000100010011;
ROM[32765] <= 32'b00000000000000010010010000000011;
ROM[32766] <= 32'b00000000011101000010010010110011;
ROM[32767] <= 32'b00000000100000111010010100110011;
ROM[32768] <= 32'b00000000101001001000001110110011;
ROM[32769] <= 32'b00000000000100111000001110010011;
ROM[32770] <= 32'b00000000000100111111001110010011;
ROM[32771] <= 32'b00000000011100010010000000100011;
ROM[32772] <= 32'b00000000010000010000000100010011;
ROM[32773] <= 32'b11111111110000010000000100010011;
ROM[32774] <= 32'b00000000000000010010001110000011;
ROM[32775] <= 32'b00000000000000111000101001100011;
ROM[32776] <= 32'b00000000000000100000001110110111;
ROM[32777] <= 32'b00000011010000111000001110010011;
ROM[32778] <= 32'b00000000111000111000001110110011;
ROM[32779] <= 32'b00000000000000111000000011100111;
ROM[32780] <= 32'b00001011110000000000000011101111;
ROM[32781] <= 32'b00000000010100010010000000100011;
ROM[32782] <= 32'b00000000010000010000000100010011;
ROM[32783] <= 32'b00000000000000100000001110110111;
ROM[32784] <= 32'b00001000100000111000001110010011;
ROM[32785] <= 32'b00000000111000111000001110110011;
ROM[32786] <= 32'b00000000011100010010000000100011;
ROM[32787] <= 32'b00000000010000010000000100010011;
ROM[32788] <= 32'b00000000001100010010000000100011;
ROM[32789] <= 32'b00000000010000010000000100010011;
ROM[32790] <= 32'b00000000010000010010000000100011;
ROM[32791] <= 32'b00000000010000010000000100010011;
ROM[32792] <= 32'b00000000010100010010000000100011;
ROM[32793] <= 32'b00000000010000010000000100010011;
ROM[32794] <= 32'b00000000011000010010000000100011;
ROM[32795] <= 32'b00000000010000010000000100010011;
ROM[32796] <= 32'b00000001010000000000001110010011;
ROM[32797] <= 32'b00000000010000111000001110010011;
ROM[32798] <= 32'b01000000011100010000001110110011;
ROM[32799] <= 32'b00000000011100000000001000110011;
ROM[32800] <= 32'b00000000001000000000000110110011;
ROM[32801] <= 32'b00001010110000000000000011101111;
ROM[32802] <= 32'b11111111110000010000000100010011;
ROM[32803] <= 32'b00000000000000010010001110000011;
ROM[32804] <= 32'b00000000011101100010000000100011;
ROM[32805] <= 32'b00000000000100000000001110010011;
ROM[32806] <= 32'b00000000011100010010000000100011;
ROM[32807] <= 32'b00000000010000010000000100010011;
ROM[32808] <= 32'b11111111110000010000000100010011;
ROM[32809] <= 32'b00000000000000010010001110000011;
ROM[32810] <= 32'b01000000011100000000001110110011;
ROM[32811] <= 32'b00000000011100010010000000100011;
ROM[32812] <= 32'b00000000010000010000000100010011;
ROM[32813] <= 32'b00000001010000000000001110010011;
ROM[32814] <= 32'b01000000011100011000001110110011;
ROM[32815] <= 32'b00000000000000111010000010000011;
ROM[32816] <= 32'b11111111110000010000000100010011;
ROM[32817] <= 32'b00000000000000010010001110000011;
ROM[32818] <= 32'b00000000011100100010000000100011;
ROM[32819] <= 32'b00000000010000100000000100010011;
ROM[32820] <= 32'b00000001010000000000001110010011;
ROM[32821] <= 32'b01000000011100011000001110110011;
ROM[32822] <= 32'b00000000010000111010000110000011;
ROM[32823] <= 32'b00000000100000111010001000000011;
ROM[32824] <= 32'b00000000110000111010001010000011;
ROM[32825] <= 32'b00000001000000111010001100000011;
ROM[32826] <= 32'b00000000000000001000000011100111;
ROM[32827] <= 32'b00000000000000000000001110010011;
ROM[32828] <= 32'b00000000011100010010000000100011;
ROM[32829] <= 32'b00000000010000010000000100010011;
ROM[32830] <= 32'b00000001010000000000001110010011;
ROM[32831] <= 32'b01000000011100011000001110110011;
ROM[32832] <= 32'b00000000000000111010000010000011;
ROM[32833] <= 32'b11111111110000010000000100010011;
ROM[32834] <= 32'b00000000000000010010001110000011;
ROM[32835] <= 32'b00000000011100100010000000100011;
ROM[32836] <= 32'b00000000010000100000000100010011;
ROM[32837] <= 32'b00000001010000000000001110010011;
ROM[32838] <= 32'b01000000011100011000001110110011;
ROM[32839] <= 32'b00000000010000111010000110000011;
ROM[32840] <= 32'b00000000100000111010001000000011;
ROM[32841] <= 32'b00000000110000111010001010000011;
ROM[32842] <= 32'b00000001000000111010001100000011;
ROM[32843] <= 32'b00000000000000001000000011100111;
ROM[32844] <= 32'b00000000000000010010000000100011;
ROM[32845] <= 32'b00000000010000010000000100010011;
ROM[32846] <= 32'b00000000000000010010000000100011;
ROM[32847] <= 32'b00000000010000010000000100010011;
ROM[32848] <= 32'b00000000000000010010000000100011;
ROM[32849] <= 32'b00000000010000010000000100010011;
ROM[32850] <= 32'b00000000000000100010001110000011;
ROM[32851] <= 32'b00000000011100010010000000100011;
ROM[32852] <= 32'b00000000010000010000000100010011;
ROM[32853] <= 32'b11111111110000010000000100010011;
ROM[32854] <= 32'b00000000000000010010001110000011;
ROM[32855] <= 32'b00000000000000111000001010010011;
ROM[32856] <= 32'b00000000110100101000010000110011;
ROM[32857] <= 32'b00000000110001000010001110000011;
ROM[32858] <= 32'b00000000011100010010000000100011;
ROM[32859] <= 32'b00000000010000010000000100010011;
ROM[32860] <= 32'b11111111110000010000000100010011;
ROM[32861] <= 32'b00000000000000010010001110000011;
ROM[32862] <= 32'b00000000011100011010000000100011;
ROM[32863] <= 32'b00000000000000000000001110010011;
ROM[32864] <= 32'b00000000011100010010000000100011;
ROM[32865] <= 32'b00000000010000010000000100010011;
ROM[32866] <= 32'b11111111110000010000000100010011;
ROM[32867] <= 32'b00000000000000010010001110000011;
ROM[32868] <= 32'b00000000011100011010010000100011;
ROM[32869] <= 32'b00000000110100101000010000110011;
ROM[32870] <= 32'b00000010100001000010001110000011;
ROM[32871] <= 32'b00000000011100010010000000100011;
ROM[32872] <= 32'b00000000010000010000000100010011;
ROM[32873] <= 32'b00000000110100101000010000110011;
ROM[32874] <= 32'b00000000110001000010001110000011;
ROM[32875] <= 32'b00000000011100010010000000100011;
ROM[32876] <= 32'b00000000010000010000000100010011;
ROM[32877] <= 32'b11111111110000010000000100010011;
ROM[32878] <= 32'b00000000000000010010001110000011;
ROM[32879] <= 32'b11111111110000010000000100010011;
ROM[32880] <= 32'b00000000000000010010010000000011;
ROM[32881] <= 32'b01000000011101000000001110110011;
ROM[32882] <= 32'b00000000011100010010000000100011;
ROM[32883] <= 32'b00000000010000010000000100010011;
ROM[32884] <= 32'b11111111110000010000000100010011;
ROM[32885] <= 32'b00000000000000010010001110000011;
ROM[32886] <= 32'b00000000011100011010001000100011;
ROM[32887] <= 32'b00000000000000011010001110000011;
ROM[32888] <= 32'b00000000011100010010000000100011;
ROM[32889] <= 32'b00000000010000010000000100010011;
ROM[32890] <= 32'b00000000000000000000001110010011;
ROM[32891] <= 32'b00000000011100010010000000100011;
ROM[32892] <= 32'b00000000010000010000000100010011;
ROM[32893] <= 32'b11111111110000010000000100010011;
ROM[32894] <= 32'b00000000000000010010001110000011;
ROM[32895] <= 32'b11111111110000010000000100010011;
ROM[32896] <= 32'b00000000000000010010010000000011;
ROM[32897] <= 32'b00000000100000111010001110110011;
ROM[32898] <= 32'b00000000011100010010000000100011;
ROM[32899] <= 32'b00000000010000010000000100010011;
ROM[32900] <= 32'b11111111110000010000000100010011;
ROM[32901] <= 32'b00000000000000010010001110000011;
ROM[32902] <= 32'b01000000011100000000001110110011;
ROM[32903] <= 32'b00000000000100111000001110010011;
ROM[32904] <= 32'b00000000011100010010000000100011;
ROM[32905] <= 32'b00000000010000010000000100010011;
ROM[32906] <= 32'b11111111110000010000000100010011;
ROM[32907] <= 32'b00000000000000010010001110000011;
ROM[32908] <= 32'b00000000000000111000101001100011;
ROM[32909] <= 32'b00000000000000100000001110110111;
ROM[32910] <= 32'b01011011100000111000001110010011;
ROM[32911] <= 32'b00000000111000111000001110110011;
ROM[32912] <= 32'b00000000000000111000000011100111;
ROM[32913] <= 32'b00000000110100101000010000110011;
ROM[32914] <= 32'b00000010000001000010001110000011;
ROM[32915] <= 32'b00000000011100010010000000100011;
ROM[32916] <= 32'b00000000010000010000000100010011;
ROM[32917] <= 32'b00000000010000011010001110000011;
ROM[32918] <= 32'b00000000011100010010000000100011;
ROM[32919] <= 32'b00000000010000010000000100010011;
ROM[32920] <= 32'b00000000010000000000001110010011;
ROM[32921] <= 32'b00000000011100010010000000100011;
ROM[32922] <= 32'b00000000010000010000000100010011;
ROM[32923] <= 32'b00000000000000100000001110110111;
ROM[32924] <= 32'b00101011100000111000001110010011;
ROM[32925] <= 32'b00000000111000111000001110110011;
ROM[32926] <= 32'b00000000011100010010000000100011;
ROM[32927] <= 32'b00000000010000010000000100010011;
ROM[32928] <= 32'b00000000001100010010000000100011;
ROM[32929] <= 32'b00000000010000010000000100010011;
ROM[32930] <= 32'b00000000010000010010000000100011;
ROM[32931] <= 32'b00000000010000010000000100010011;
ROM[32932] <= 32'b00000000010100010010000000100011;
ROM[32933] <= 32'b00000000010000010000000100010011;
ROM[32934] <= 32'b00000000011000010010000000100011;
ROM[32935] <= 32'b00000000010000010000000100010011;
ROM[32936] <= 32'b00000001010000000000001110010011;
ROM[32937] <= 32'b00000000100000111000001110010011;
ROM[32938] <= 32'b01000000011100010000001110110011;
ROM[32939] <= 32'b00000000011100000000001000110011;
ROM[32940] <= 32'b00000000001000000000000110110011;
ROM[32941] <= 32'b11010111100011110001000011101111;
ROM[32942] <= 32'b11111111110000010000000100010011;
ROM[32943] <= 32'b00000000000000010010001110000011;
ROM[32944] <= 32'b11111111110000010000000100010011;
ROM[32945] <= 32'b00000000000000010010010000000011;
ROM[32946] <= 32'b00000000011101000000001110110011;
ROM[32947] <= 32'b00000000011100010010000000100011;
ROM[32948] <= 32'b00000000010000010000000100010011;
ROM[32949] <= 32'b11111111110000010000000100010011;
ROM[32950] <= 32'b00000000000000010010001110000011;
ROM[32951] <= 32'b00000000000000111000001100010011;
ROM[32952] <= 32'b00000000110100110000010000110011;
ROM[32953] <= 32'b00000000000001000010001110000011;
ROM[32954] <= 32'b00000000011100010010000000100011;
ROM[32955] <= 32'b00000000010000010000000100010011;
ROM[32956] <= 32'b00000000110100101000010000110011;
ROM[32957] <= 32'b00000010000001000010001110000011;
ROM[32958] <= 32'b00000000011100010010000000100011;
ROM[32959] <= 32'b00000000010000010000000100010011;
ROM[32960] <= 32'b00000000100000011010001110000011;
ROM[32961] <= 32'b00000000011100010010000000100011;
ROM[32962] <= 32'b00000000010000010000000100010011;
ROM[32963] <= 32'b00000000010000000000001110010011;
ROM[32964] <= 32'b00000000011100010010000000100011;
ROM[32965] <= 32'b00000000010000010000000100010011;
ROM[32966] <= 32'b00000000000000100000001110110111;
ROM[32967] <= 32'b00110110010000111000001110010011;
ROM[32968] <= 32'b00000000111000111000001110110011;
ROM[32969] <= 32'b00000000011100010010000000100011;
ROM[32970] <= 32'b00000000010000010000000100010011;
ROM[32971] <= 32'b00000000001100010010000000100011;
ROM[32972] <= 32'b00000000010000010000000100010011;
ROM[32973] <= 32'b00000000010000010010000000100011;
ROM[32974] <= 32'b00000000010000010000000100010011;
ROM[32975] <= 32'b00000000010100010010000000100011;
ROM[32976] <= 32'b00000000010000010000000100010011;
ROM[32977] <= 32'b00000000011000010010000000100011;
ROM[32978] <= 32'b00000000010000010000000100010011;
ROM[32979] <= 32'b00000001010000000000001110010011;
ROM[32980] <= 32'b00000000100000111000001110010011;
ROM[32981] <= 32'b01000000011100010000001110110011;
ROM[32982] <= 32'b00000000011100000000001000110011;
ROM[32983] <= 32'b00000000001000000000000110110011;
ROM[32984] <= 32'b11001100110011110001000011101111;
ROM[32985] <= 32'b11111111110000010000000100010011;
ROM[32986] <= 32'b00000000000000010010001110000011;
ROM[32987] <= 32'b11111111110000010000000100010011;
ROM[32988] <= 32'b00000000000000010010010000000011;
ROM[32989] <= 32'b00000000011101000000001110110011;
ROM[32990] <= 32'b00000000011100010010000000100011;
ROM[32991] <= 32'b00000000010000010000000100010011;
ROM[32992] <= 32'b11111111110000010000000100010011;
ROM[32993] <= 32'b00000000000000010010001110000011;
ROM[32994] <= 32'b00000000000000111000001100010011;
ROM[32995] <= 32'b11111111110000010000000100010011;
ROM[32996] <= 32'b00000000000000010010001110000011;
ROM[32997] <= 32'b00000000110100110000010000110011;
ROM[32998] <= 32'b00000000011101000010000000100011;
ROM[32999] <= 32'b00000000110100101000010000110011;
ROM[33000] <= 32'b00000010010001000010001110000011;
ROM[33001] <= 32'b00000000011100010010000000100011;
ROM[33002] <= 32'b00000000010000010000000100010011;
ROM[33003] <= 32'b00000000010000011010001110000011;
ROM[33004] <= 32'b00000000011100010010000000100011;
ROM[33005] <= 32'b00000000010000010000000100010011;
ROM[33006] <= 32'b00000000010000000000001110010011;
ROM[33007] <= 32'b00000000011100010010000000100011;
ROM[33008] <= 32'b00000000010000010000000100010011;
ROM[33009] <= 32'b00000000000000100000001110110111;
ROM[33010] <= 32'b01000001000000111000001110010011;
ROM[33011] <= 32'b00000000111000111000001110110011;
ROM[33012] <= 32'b00000000011100010010000000100011;
ROM[33013] <= 32'b00000000010000010000000100010011;
ROM[33014] <= 32'b00000000001100010010000000100011;
ROM[33015] <= 32'b00000000010000010000000100010011;
ROM[33016] <= 32'b00000000010000010010000000100011;
ROM[33017] <= 32'b00000000010000010000000100010011;
ROM[33018] <= 32'b00000000010100010010000000100011;
ROM[33019] <= 32'b00000000010000010000000100010011;
ROM[33020] <= 32'b00000000011000010010000000100011;
ROM[33021] <= 32'b00000000010000010000000100010011;
ROM[33022] <= 32'b00000001010000000000001110010011;
ROM[33023] <= 32'b00000000100000111000001110010011;
ROM[33024] <= 32'b01000000011100010000001110110011;
ROM[33025] <= 32'b00000000011100000000001000110011;
ROM[33026] <= 32'b00000000001000000000000110110011;
ROM[33027] <= 32'b11000010000011110001000011101111;
ROM[33028] <= 32'b11111111110000010000000100010011;
ROM[33029] <= 32'b00000000000000010010001110000011;
ROM[33030] <= 32'b11111111110000010000000100010011;
ROM[33031] <= 32'b00000000000000010010010000000011;
ROM[33032] <= 32'b00000000011101000000001110110011;
ROM[33033] <= 32'b00000000011100010010000000100011;
ROM[33034] <= 32'b00000000010000010000000100010011;
ROM[33035] <= 32'b11111111110000010000000100010011;
ROM[33036] <= 32'b00000000000000010010001110000011;
ROM[33037] <= 32'b00000000000000111000001100010011;
ROM[33038] <= 32'b00000000110100110000010000110011;
ROM[33039] <= 32'b00000000000001000010001110000011;
ROM[33040] <= 32'b00000000011100010010000000100011;
ROM[33041] <= 32'b00000000010000010000000100010011;
ROM[33042] <= 32'b00000000110100101000010000110011;
ROM[33043] <= 32'b00000010010001000010001110000011;
ROM[33044] <= 32'b00000000011100010010000000100011;
ROM[33045] <= 32'b00000000010000010000000100010011;
ROM[33046] <= 32'b00000000100000011010001110000011;
ROM[33047] <= 32'b00000000011100010010000000100011;
ROM[33048] <= 32'b00000000010000010000000100010011;
ROM[33049] <= 32'b00000000010000000000001110010011;
ROM[33050] <= 32'b00000000011100010010000000100011;
ROM[33051] <= 32'b00000000010000010000000100010011;
ROM[33052] <= 32'b00000000000000100000001110110111;
ROM[33053] <= 32'b01001011110000111000001110010011;
ROM[33054] <= 32'b00000000111000111000001110110011;
ROM[33055] <= 32'b00000000011100010010000000100011;
ROM[33056] <= 32'b00000000010000010000000100010011;
ROM[33057] <= 32'b00000000001100010010000000100011;
ROM[33058] <= 32'b00000000010000010000000100010011;
ROM[33059] <= 32'b00000000010000010010000000100011;
ROM[33060] <= 32'b00000000010000010000000100010011;
ROM[33061] <= 32'b00000000010100010010000000100011;
ROM[33062] <= 32'b00000000010000010000000100010011;
ROM[33063] <= 32'b00000000011000010010000000100011;
ROM[33064] <= 32'b00000000010000010000000100010011;
ROM[33065] <= 32'b00000001010000000000001110010011;
ROM[33066] <= 32'b00000000100000111000001110010011;
ROM[33067] <= 32'b01000000011100010000001110110011;
ROM[33068] <= 32'b00000000011100000000001000110011;
ROM[33069] <= 32'b00000000001000000000000110110011;
ROM[33070] <= 32'b10110111010011110001000011101111;
ROM[33071] <= 32'b11111111110000010000000100010011;
ROM[33072] <= 32'b00000000000000010010001110000011;
ROM[33073] <= 32'b11111111110000010000000100010011;
ROM[33074] <= 32'b00000000000000010010010000000011;
ROM[33075] <= 32'b00000000011101000000001110110011;
ROM[33076] <= 32'b00000000011100010010000000100011;
ROM[33077] <= 32'b00000000010000010000000100010011;
ROM[33078] <= 32'b11111111110000010000000100010011;
ROM[33079] <= 32'b00000000000000010010001110000011;
ROM[33080] <= 32'b00000000000000111000001100010011;
ROM[33081] <= 32'b11111111110000010000000100010011;
ROM[33082] <= 32'b00000000000000010010001110000011;
ROM[33083] <= 32'b00000000110100110000010000110011;
ROM[33084] <= 32'b00000000011101000010000000100011;
ROM[33085] <= 32'b00000000010000011010001110000011;
ROM[33086] <= 32'b00000000011100010010000000100011;
ROM[33087] <= 32'b00000000010000010000000100010011;
ROM[33088] <= 32'b00000000000100000000001110010011;
ROM[33089] <= 32'b00000000011100010010000000100011;
ROM[33090] <= 32'b00000000010000010000000100010011;
ROM[33091] <= 32'b11111111110000010000000100010011;
ROM[33092] <= 32'b00000000000000010010001110000011;
ROM[33093] <= 32'b11111111110000010000000100010011;
ROM[33094] <= 32'b00000000000000010010010000000011;
ROM[33095] <= 32'b00000000011101000000001110110011;
ROM[33096] <= 32'b00000000011100010010000000100011;
ROM[33097] <= 32'b00000000010000010000000100010011;
ROM[33098] <= 32'b11111111110000010000000100010011;
ROM[33099] <= 32'b00000000000000010010001110000011;
ROM[33100] <= 32'b00000000011100011010001000100011;
ROM[33101] <= 32'b00000000100000011010001110000011;
ROM[33102] <= 32'b00000000011100010010000000100011;
ROM[33103] <= 32'b00000000010000010000000100010011;
ROM[33104] <= 32'b00000000000100000000001110010011;
ROM[33105] <= 32'b00000000011100010010000000100011;
ROM[33106] <= 32'b00000000010000010000000100010011;
ROM[33107] <= 32'b11111111110000010000000100010011;
ROM[33108] <= 32'b00000000000000010010001110000011;
ROM[33109] <= 32'b11111111110000010000000100010011;
ROM[33110] <= 32'b00000000000000010010010000000011;
ROM[33111] <= 32'b00000000011101000000001110110011;
ROM[33112] <= 32'b00000000011100010010000000100011;
ROM[33113] <= 32'b00000000010000010000000100010011;
ROM[33114] <= 32'b11111111110000010000000100010011;
ROM[33115] <= 32'b00000000000000010010001110000011;
ROM[33116] <= 32'b00000000011100011010010000100011;
ROM[33117] <= 32'b00000000000000011010001110000011;
ROM[33118] <= 32'b00000000011100010010000000100011;
ROM[33119] <= 32'b00000000010000010000000100010011;
ROM[33120] <= 32'b00000000000100000000001110010011;
ROM[33121] <= 32'b00000000011100010010000000100011;
ROM[33122] <= 32'b00000000010000010000000100010011;
ROM[33123] <= 32'b11111111110000010000000100010011;
ROM[33124] <= 32'b00000000000000010010001110000011;
ROM[33125] <= 32'b11111111110000010000000100010011;
ROM[33126] <= 32'b00000000000000010010010000000011;
ROM[33127] <= 32'b01000000011101000000001110110011;
ROM[33128] <= 32'b00000000011100010010000000100011;
ROM[33129] <= 32'b00000000010000010000000100010011;
ROM[33130] <= 32'b11111111110000010000000100010011;
ROM[33131] <= 32'b00000000000000010010001110000011;
ROM[33132] <= 32'b00000000011100011010000000100011;
ROM[33133] <= 32'b11000010100111111111000011101111;
ROM[33134] <= 32'b00000000000000000000001110010011;
ROM[33135] <= 32'b00000000011100010010000000100011;
ROM[33136] <= 32'b00000000010000010000000100010011;
ROM[33137] <= 32'b00000001010000000000001110010011;
ROM[33138] <= 32'b01000000011100011000001110110011;
ROM[33139] <= 32'b00000000000000111010000010000011;
ROM[33140] <= 32'b11111111110000010000000100010011;
ROM[33141] <= 32'b00000000000000010010001110000011;
ROM[33142] <= 32'b00000000011100100010000000100011;
ROM[33143] <= 32'b00000000010000100000000100010011;
ROM[33144] <= 32'b00000001010000000000001110010011;
ROM[33145] <= 32'b01000000011100011000001110110011;
ROM[33146] <= 32'b00000000010000111010000110000011;
ROM[33147] <= 32'b00000000100000111010001000000011;
ROM[33148] <= 32'b00000000110000111010001010000011;
ROM[33149] <= 32'b00000001000000111010001100000011;
ROM[33150] <= 32'b00000000000000001000000011100111;
ROM[33151] <= 32'b00000000000000100010001110000011;
ROM[33152] <= 32'b00000000011100010010000000100011;
ROM[33153] <= 32'b00000000010000010000000100010011;
ROM[33154] <= 32'b11111111110000010000000100010011;
ROM[33155] <= 32'b00000000000000010010001110000011;
ROM[33156] <= 32'b00000000000000111000001010010011;
ROM[33157] <= 32'b00000000110100101000010000110011;
ROM[33158] <= 32'b00000000010001000010001110000011;
ROM[33159] <= 32'b00000000011100010010000000100011;
ROM[33160] <= 32'b00000000010000010000000100010011;
ROM[33161] <= 32'b00000001010000000000001110010011;
ROM[33162] <= 32'b01000000011100011000001110110011;
ROM[33163] <= 32'b00000000000000111010000010000011;
ROM[33164] <= 32'b11111111110000010000000100010011;
ROM[33165] <= 32'b00000000000000010010001110000011;
ROM[33166] <= 32'b00000000011100100010000000100011;
ROM[33167] <= 32'b00000000010000100000000100010011;
ROM[33168] <= 32'b00000001010000000000001110010011;
ROM[33169] <= 32'b01000000011100011000001110110011;
ROM[33170] <= 32'b00000000010000111010000110000011;
ROM[33171] <= 32'b00000000100000111010001000000011;
ROM[33172] <= 32'b00000000110000111010001010000011;
ROM[33173] <= 32'b00000001000000111010001100000011;
ROM[33174] <= 32'b00000000000000001000000011100111;
ROM[33175] <= 32'b00000000000000100010001110000011;
ROM[33176] <= 32'b00000000011100010010000000100011;
ROM[33177] <= 32'b00000000010000010000000100010011;
ROM[33178] <= 32'b11111111110000010000000100010011;
ROM[33179] <= 32'b00000000000000010010001110000011;
ROM[33180] <= 32'b00000000000000111000001010010011;
ROM[33181] <= 32'b00000000110100101000010000110011;
ROM[33182] <= 32'b00000000100001000010001110000011;
ROM[33183] <= 32'b00000000011100010010000000100011;
ROM[33184] <= 32'b00000000010000010000000100010011;
ROM[33185] <= 32'b00000001010000000000001110010011;
ROM[33186] <= 32'b01000000011100011000001110110011;
ROM[33187] <= 32'b00000000000000111010000010000011;
ROM[33188] <= 32'b11111111110000010000000100010011;
ROM[33189] <= 32'b00000000000000010010001110000011;
ROM[33190] <= 32'b00000000011100100010000000100011;
ROM[33191] <= 32'b00000000010000100000000100010011;
ROM[33192] <= 32'b00000001010000000000001110010011;
ROM[33193] <= 32'b01000000011100011000001110110011;
ROM[33194] <= 32'b00000000010000111010000110000011;
ROM[33195] <= 32'b00000000100000111010001000000011;
ROM[33196] <= 32'b00000000110000111010001010000011;
ROM[33197] <= 32'b00000001000000111010001100000011;
ROM[33198] <= 32'b00000000000000001000000011100111;
ROM[33199] <= 32'b00000000000000100010001110000011;
ROM[33200] <= 32'b00000000011100010010000000100011;
ROM[33201] <= 32'b00000000010000010000000100010011;
ROM[33202] <= 32'b11111111110000010000000100010011;
ROM[33203] <= 32'b00000000000000010010001110000011;
ROM[33204] <= 32'b00000000000000111000001010010011;
ROM[33205] <= 32'b00000000110100101000010000110011;
ROM[33206] <= 32'b00000000110001000010001110000011;
ROM[33207] <= 32'b00000000011100010010000000100011;
ROM[33208] <= 32'b00000000010000010000000100010011;
ROM[33209] <= 32'b00000001010000000000001110010011;
ROM[33210] <= 32'b01000000011100011000001110110011;
ROM[33211] <= 32'b00000000000000111010000010000011;
ROM[33212] <= 32'b11111111110000010000000100010011;
ROM[33213] <= 32'b00000000000000010010001110000011;
ROM[33214] <= 32'b00000000011100100010000000100011;
ROM[33215] <= 32'b00000000010000100000000100010011;
ROM[33216] <= 32'b00000001010000000000001110010011;
ROM[33217] <= 32'b01000000011100011000001110110011;
ROM[33218] <= 32'b00000000010000111010000110000011;
ROM[33219] <= 32'b00000000100000111010001000000011;
ROM[33220] <= 32'b00000000110000111010001010000011;
ROM[33221] <= 32'b00000001000000111010001100000011;
ROM[33222] <= 32'b00000000000000001000000011100111;
ROM[33223] <= 32'b00000000000000100010001110000011;
ROM[33224] <= 32'b00000000011100010010000000100011;
ROM[33225] <= 32'b00000000010000010000000100010011;
ROM[33226] <= 32'b11111111110000010000000100010011;
ROM[33227] <= 32'b00000000000000010010001110000011;
ROM[33228] <= 32'b00000000000000111000001010010011;
ROM[33229] <= 32'b00000000110100101000010000110011;
ROM[33230] <= 32'b00000001100001000010001110000011;
ROM[33231] <= 32'b00000000011100010010000000100011;
ROM[33232] <= 32'b00000000010000010000000100010011;
ROM[33233] <= 32'b00000001010000000000001110010011;
ROM[33234] <= 32'b01000000011100011000001110110011;
ROM[33235] <= 32'b00000000000000111010000010000011;
ROM[33236] <= 32'b11111111110000010000000100010011;
ROM[33237] <= 32'b00000000000000010010001110000011;
ROM[33238] <= 32'b00000000011100100010000000100011;
ROM[33239] <= 32'b00000000010000100000000100010011;
ROM[33240] <= 32'b00000001010000000000001110010011;
ROM[33241] <= 32'b01000000011100011000001110110011;
ROM[33242] <= 32'b00000000010000111010000110000011;
ROM[33243] <= 32'b00000000100000111010001000000011;
ROM[33244] <= 32'b00000000110000111010001010000011;
ROM[33245] <= 32'b00000001000000111010001100000011;
ROM[33246] <= 32'b00000000000000001000000011100111;
ROM[33247] <= 32'b00000000000000100010001110000011;
ROM[33248] <= 32'b00000000011100010010000000100011;
ROM[33249] <= 32'b00000000010000010000000100010011;
ROM[33250] <= 32'b11111111110000010000000100010011;
ROM[33251] <= 32'b00000000000000010010001110000011;
ROM[33252] <= 32'b00000000000000111000001010010011;
ROM[33253] <= 32'b00000000110100101000010000110011;
ROM[33254] <= 32'b00000001110001000010001110000011;
ROM[33255] <= 32'b00000000011100010010000000100011;
ROM[33256] <= 32'b00000000010000010000000100010011;
ROM[33257] <= 32'b00000001010000000000001110010011;
ROM[33258] <= 32'b01000000011100011000001110110011;
ROM[33259] <= 32'b00000000000000111010000010000011;
ROM[33260] <= 32'b11111111110000010000000100010011;
ROM[33261] <= 32'b00000000000000010010001110000011;
ROM[33262] <= 32'b00000000011100100010000000100011;
ROM[33263] <= 32'b00000000010000100000000100010011;
ROM[33264] <= 32'b00000001010000000000001110010011;
ROM[33265] <= 32'b01000000011100011000001110110011;
ROM[33266] <= 32'b00000000010000111010000110000011;
ROM[33267] <= 32'b00000000100000111010001000000011;
ROM[33268] <= 32'b00000000110000111010001010000011;
ROM[33269] <= 32'b00000001000000111010001100000011;
ROM[33270] <= 32'b00000000000000001000000011100111;
ROM[33271] <= 32'b00000000000000100010001110000011;
ROM[33272] <= 32'b00000000011100010010000000100011;
ROM[33273] <= 32'b00000000010000010000000100010011;
ROM[33274] <= 32'b11111111110000010000000100010011;
ROM[33275] <= 32'b00000000000000010010001110000011;
ROM[33276] <= 32'b00000000000000111000001010010011;
ROM[33277] <= 32'b00000000010000100010001110000011;
ROM[33278] <= 32'b00000000011100010010000000100011;
ROM[33279] <= 32'b00000000010000010000000100010011;
ROM[33280] <= 32'b11111111110000010000000100010011;
ROM[33281] <= 32'b00000000000000010010001110000011;
ROM[33282] <= 32'b00000000110100101000010000110011;
ROM[33283] <= 32'b00000000011101000010110000100011;
ROM[33284] <= 32'b00000000000000000000001110010011;
ROM[33285] <= 32'b00000000011100010010000000100011;
ROM[33286] <= 32'b00000000010000010000000100010011;
ROM[33287] <= 32'b00000001010000000000001110010011;
ROM[33288] <= 32'b01000000011100011000001110110011;
ROM[33289] <= 32'b00000000000000111010000010000011;
ROM[33290] <= 32'b11111111110000010000000100010011;
ROM[33291] <= 32'b00000000000000010010001110000011;
ROM[33292] <= 32'b00000000011100100010000000100011;
ROM[33293] <= 32'b00000000010000100000000100010011;
ROM[33294] <= 32'b00000001010000000000001110010011;
ROM[33295] <= 32'b01000000011100011000001110110011;
ROM[33296] <= 32'b00000000010000111010000110000011;
ROM[33297] <= 32'b00000000100000111010001000000011;
ROM[33298] <= 32'b00000000110000111010001010000011;
ROM[33299] <= 32'b00000001000000111010001100000011;
ROM[33300] <= 32'b00000000000000001000000011100111;
ROM[33301] <= 32'b00000000000000100010001110000011;
ROM[33302] <= 32'b00000000011100010010000000100011;
ROM[33303] <= 32'b00000000010000010000000100010011;
ROM[33304] <= 32'b11111111110000010000000100010011;
ROM[33305] <= 32'b00000000000000010010001110000011;
ROM[33306] <= 32'b00000000000000111000001010010011;
ROM[33307] <= 32'b00000000110100101000010000110011;
ROM[33308] <= 32'b00000001100001000010001110000011;
ROM[33309] <= 32'b00000000011100010010000000100011;
ROM[33310] <= 32'b00000000010000010000000100010011;
ROM[33311] <= 32'b11111111110000010000000100010011;
ROM[33312] <= 32'b00000000000000010010001110000011;
ROM[33313] <= 32'b00000000110100101000010000110011;
ROM[33314] <= 32'b00000000011101000010111000100011;
ROM[33315] <= 32'b00000000000000000000001110010011;
ROM[33316] <= 32'b00000000011100010010000000100011;
ROM[33317] <= 32'b00000000010000010000000100010011;
ROM[33318] <= 32'b00000001010000000000001110010011;
ROM[33319] <= 32'b01000000011100011000001110110011;
ROM[33320] <= 32'b00000000000000111010000010000011;
ROM[33321] <= 32'b11111111110000010000000100010011;
ROM[33322] <= 32'b00000000000000010010001110000011;
ROM[33323] <= 32'b00000000011100100010000000100011;
ROM[33324] <= 32'b00000000010000100000000100010011;
ROM[33325] <= 32'b00000001010000000000001110010011;
ROM[33326] <= 32'b01000000011100011000001110110011;
ROM[33327] <= 32'b00000000010000111010000110000011;
ROM[33328] <= 32'b00000000100000111010001000000011;
ROM[33329] <= 32'b00000000110000111010001010000011;
ROM[33330] <= 32'b00000001000000111010001100000011;
ROM[33331] <= 32'b00000000000000001000000011100111;
ROM[33332] <= 32'b00000000000000010010000000100011;
ROM[33333] <= 32'b00000000010000010000000100010011;
ROM[33334] <= 32'b00000000000000100010001110000011;
ROM[33335] <= 32'b00000000011100010010000000100011;
ROM[33336] <= 32'b00000000010000010000000100010011;
ROM[33337] <= 32'b11111111110000010000000100010011;
ROM[33338] <= 32'b00000000000000010010001110000011;
ROM[33339] <= 32'b00000000000000111000001010010011;
ROM[33340] <= 32'b00000000110100101000010000110011;
ROM[33341] <= 32'b00000000000001000010001110000011;
ROM[33342] <= 32'b00000000011100010010000000100011;
ROM[33343] <= 32'b00000000010000010000000100010011;
ROM[33344] <= 32'b00000000000000100001001110110111;
ROM[33345] <= 32'b10010100110000111000001110010011;
ROM[33346] <= 32'b00000000111000111000001110110011;
ROM[33347] <= 32'b00000000011100010010000000100011;
ROM[33348] <= 32'b00000000010000010000000100010011;
ROM[33349] <= 32'b00000000001100010010000000100011;
ROM[33350] <= 32'b00000000010000010000000100010011;
ROM[33351] <= 32'b00000000010000010010000000100011;
ROM[33352] <= 32'b00000000010000010000000100010011;
ROM[33353] <= 32'b00000000010100010010000000100011;
ROM[33354] <= 32'b00000000010000010000000100010011;
ROM[33355] <= 32'b00000000011000010010000000100011;
ROM[33356] <= 32'b00000000010000010000000100010011;
ROM[33357] <= 32'b00000001010000000000001110010011;
ROM[33358] <= 32'b00000000010000111000001110010011;
ROM[33359] <= 32'b01000000011100010000001110110011;
ROM[33360] <= 32'b00000000011100000000001000110011;
ROM[33361] <= 32'b00000000001000000000000110110011;
ROM[33362] <= 32'b00010001110000000011000011101111;
ROM[33363] <= 32'b11111111110000010000000100010011;
ROM[33364] <= 32'b00000000000000010010001110000011;
ROM[33365] <= 32'b00000000011100011010000000100011;
ROM[33366] <= 32'b00000000110100101000010000110011;
ROM[33367] <= 32'b00000001100001000010001110000011;
ROM[33368] <= 32'b00000000011100010010000000100011;
ROM[33369] <= 32'b00000000010000010000000100010011;
ROM[33370] <= 32'b00000000000100000000001110010011;
ROM[33371] <= 32'b00000000011100010010000000100011;
ROM[33372] <= 32'b00000000010000010000000100010011;
ROM[33373] <= 32'b11111111110000010000000100010011;
ROM[33374] <= 32'b00000000000000010010001110000011;
ROM[33375] <= 32'b11111111110000010000000100010011;
ROM[33376] <= 32'b00000000000000010010010000000011;
ROM[33377] <= 32'b00000000011101000010010010110011;
ROM[33378] <= 32'b00000000100000111010010100110011;
ROM[33379] <= 32'b00000000101001001000001110110011;
ROM[33380] <= 32'b00000000000100111000001110010011;
ROM[33381] <= 32'b00000000000100111111001110010011;
ROM[33382] <= 32'b00000000011100010010000000100011;
ROM[33383] <= 32'b00000000010000010000000100010011;
ROM[33384] <= 32'b11111111110000010000000100010011;
ROM[33385] <= 32'b00000000000000010010001110000011;
ROM[33386] <= 32'b00000000000000111000101001100011;
ROM[33387] <= 32'b00000000000000100001001110110111;
ROM[33388] <= 32'b10011100000000111000001110010011;
ROM[33389] <= 32'b00000000111000111000001110110011;
ROM[33390] <= 32'b00000000000000111000000011100111;
ROM[33391] <= 32'b00001111100000000000000011101111;
ROM[33392] <= 32'b00000000110100101000010000110011;
ROM[33393] <= 32'b00000000100001000010001110000011;
ROM[33394] <= 32'b00000000011100010010000000100011;
ROM[33395] <= 32'b00000000010000010000000100010011;
ROM[33396] <= 32'b00000000000000000000001110010011;
ROM[33397] <= 32'b00000000011100010010000000100011;
ROM[33398] <= 32'b00000000010000010000000100010011;
ROM[33399] <= 32'b11111111110000010000000100010011;
ROM[33400] <= 32'b00000000000000010010001110000011;
ROM[33401] <= 32'b11111111110000010000000100010011;
ROM[33402] <= 32'b00000000000000010010010000000011;
ROM[33403] <= 32'b00000000011101000010010010110011;
ROM[33404] <= 32'b00000000100000111010010100110011;
ROM[33405] <= 32'b00000000101001001000001110110011;
ROM[33406] <= 32'b00000000000100111000001110010011;
ROM[33407] <= 32'b00000000000100111111001110010011;
ROM[33408] <= 32'b00000000011100010010000000100011;
ROM[33409] <= 32'b00000000010000010000000100010011;
ROM[33410] <= 32'b11111111110000010000000100010011;
ROM[33411] <= 32'b00000000000000010010001110000011;
ROM[33412] <= 32'b00000000000000111000101001100011;
ROM[33413] <= 32'b00000000000000100001001110110111;
ROM[33414] <= 32'b10100111000000111000001110010011;
ROM[33415] <= 32'b00000000111000111000001110110011;
ROM[33416] <= 32'b00000000000000111000000011100111;
ROM[33417] <= 32'b00000000110100101000010000110011;
ROM[33418] <= 32'b00000000100001000010001110000011;
ROM[33419] <= 32'b00000000011100010010000000100011;
ROM[33420] <= 32'b00000000010000010000000100010011;
ROM[33421] <= 32'b00000000000100000000001110010011;
ROM[33422] <= 32'b00000000011100010010000000100011;
ROM[33423] <= 32'b00000000010000010000000100010011;
ROM[33424] <= 32'b11111111110000010000000100010011;
ROM[33425] <= 32'b00000000000000010010001110000011;
ROM[33426] <= 32'b11111111110000010000000100010011;
ROM[33427] <= 32'b00000000000000010010010000000011;
ROM[33428] <= 32'b01000000011101000000001110110011;
ROM[33429] <= 32'b00000000011100010010000000100011;
ROM[33430] <= 32'b00000000010000010000000100010011;
ROM[33431] <= 32'b11111111110000010000000100010011;
ROM[33432] <= 32'b00000000000000010010001110000011;
ROM[33433] <= 32'b00000000110100101000010000110011;
ROM[33434] <= 32'b00000000011101000010010000100011;
ROM[33435] <= 32'b00000100100000000000000011101111;
ROM[33436] <= 32'b00000000000000000000001110010011;
ROM[33437] <= 32'b00000000011100010010000000100011;
ROM[33438] <= 32'b00000000010000010000000100010011;
ROM[33439] <= 32'b00000001010000000000001110010011;
ROM[33440] <= 32'b01000000011100011000001110110011;
ROM[33441] <= 32'b00000000000000111010000010000011;
ROM[33442] <= 32'b11111111110000010000000100010011;
ROM[33443] <= 32'b00000000000000010010001110000011;
ROM[33444] <= 32'b00000000011100100010000000100011;
ROM[33445] <= 32'b00000000010000100000000100010011;
ROM[33446] <= 32'b00000001010000000000001110010011;
ROM[33447] <= 32'b01000000011100011000001110110011;
ROM[33448] <= 32'b00000000010000111010000110000011;
ROM[33449] <= 32'b00000000100000111010001000000011;
ROM[33450] <= 32'b00000000110000111010001010000011;
ROM[33451] <= 32'b00000001000000111010001100000011;
ROM[33452] <= 32'b00000000000000001000000011100111;
ROM[33453] <= 32'b00000000110100101000010000110011;
ROM[33454] <= 32'b00000001100001000010001110000011;
ROM[33455] <= 32'b00000000011100010010000000100011;
ROM[33456] <= 32'b00000000010000010000000100010011;
ROM[33457] <= 32'b00000000001000000000001110010011;
ROM[33458] <= 32'b00000000011100010010000000100011;
ROM[33459] <= 32'b00000000010000010000000100010011;
ROM[33460] <= 32'b11111111110000010000000100010011;
ROM[33461] <= 32'b00000000000000010010001110000011;
ROM[33462] <= 32'b11111111110000010000000100010011;
ROM[33463] <= 32'b00000000000000010010010000000011;
ROM[33464] <= 32'b00000000011101000010010010110011;
ROM[33465] <= 32'b00000000100000111010010100110011;
ROM[33466] <= 32'b00000000101001001000001110110011;
ROM[33467] <= 32'b00000000000100111000001110010011;
ROM[33468] <= 32'b00000000000100111111001110010011;
ROM[33469] <= 32'b00000000011100010010000000100011;
ROM[33470] <= 32'b00000000010000010000000100010011;
ROM[33471] <= 32'b11111111110000010000000100010011;
ROM[33472] <= 32'b00000000000000010010001110000011;
ROM[33473] <= 32'b00000000000000111000101001100011;
ROM[33474] <= 32'b00000000000000100001001110110111;
ROM[33475] <= 32'b10110001110000111000001110010011;
ROM[33476] <= 32'b00000000111000111000001110110011;
ROM[33477] <= 32'b00000000000000111000000011100111;
ROM[33478] <= 32'b00010100010000000000000011101111;
ROM[33479] <= 32'b00000000110100101000010000110011;
ROM[33480] <= 32'b00000000100001000010001110000011;
ROM[33481] <= 32'b00000000011100010010000000100011;
ROM[33482] <= 32'b00000000010000010000000100010011;
ROM[33483] <= 32'b00000000000000011010001110000011;
ROM[33484] <= 32'b00000000011100010010000000100011;
ROM[33485] <= 32'b00000000010000010000000100010011;
ROM[33486] <= 32'b00000000000000100001001110110111;
ROM[33487] <= 32'b10111000010000111000001110010011;
ROM[33488] <= 32'b00000000111000111000001110110011;
ROM[33489] <= 32'b00000000011100010010000000100011;
ROM[33490] <= 32'b00000000010000010000000100010011;
ROM[33491] <= 32'b00000000001100010010000000100011;
ROM[33492] <= 32'b00000000010000010000000100010011;
ROM[33493] <= 32'b00000000010000010010000000100011;
ROM[33494] <= 32'b00000000010000010000000100010011;
ROM[33495] <= 32'b00000000010100010010000000100011;
ROM[33496] <= 32'b00000000010000010000000100010011;
ROM[33497] <= 32'b00000000011000010010000000100011;
ROM[33498] <= 32'b00000000010000010000000100010011;
ROM[33499] <= 32'b00000001010000000000001110010011;
ROM[33500] <= 32'b00000000010000111000001110010011;
ROM[33501] <= 32'b01000000011100010000001110110011;
ROM[33502] <= 32'b00000000011100000000001000110011;
ROM[33503] <= 32'b00000000001000000000000110110011;
ROM[33504] <= 32'b01000111100000000101000011101111;
ROM[33505] <= 32'b11111111110000010000000100010011;
ROM[33506] <= 32'b00000000000000010010001110000011;
ROM[33507] <= 32'b11111111110000010000000100010011;
ROM[33508] <= 32'b00000000000000010010010000000011;
ROM[33509] <= 32'b00000000011101000010010010110011;
ROM[33510] <= 32'b00000000100000111010010100110011;
ROM[33511] <= 32'b00000000101001001000001110110011;
ROM[33512] <= 32'b00000000000100111000001110010011;
ROM[33513] <= 32'b00000000000100111111001110010011;
ROM[33514] <= 32'b00000000011100010010000000100011;
ROM[33515] <= 32'b00000000010000010000000100010011;
ROM[33516] <= 32'b11111111110000010000000100010011;
ROM[33517] <= 32'b00000000000000010010001110000011;
ROM[33518] <= 32'b00000000000000111000101001100011;
ROM[33519] <= 32'b00000000000000100001001110110111;
ROM[33520] <= 32'b11000001100000111000001110010011;
ROM[33521] <= 32'b00000000111000111000001110110011;
ROM[33522] <= 32'b00000000000000111000000011100111;
ROM[33523] <= 32'b00000000110100101000010000110011;
ROM[33524] <= 32'b00000000100001000010001110000011;
ROM[33525] <= 32'b00000000011100010010000000100011;
ROM[33526] <= 32'b00000000010000010000000100010011;
ROM[33527] <= 32'b00000000000100000000001110010011;
ROM[33528] <= 32'b00000000011100010010000000100011;
ROM[33529] <= 32'b00000000010000010000000100010011;
ROM[33530] <= 32'b11111111110000010000000100010011;
ROM[33531] <= 32'b00000000000000010010001110000011;
ROM[33532] <= 32'b11111111110000010000000100010011;
ROM[33533] <= 32'b00000000000000010010010000000011;
ROM[33534] <= 32'b00000000011101000000001110110011;
ROM[33535] <= 32'b00000000011100010010000000100011;
ROM[33536] <= 32'b00000000010000010000000100010011;
ROM[33537] <= 32'b11111111110000010000000100010011;
ROM[33538] <= 32'b00000000000000010010001110000011;
ROM[33539] <= 32'b00000000110100101000010000110011;
ROM[33540] <= 32'b00000000011101000010010000100011;
ROM[33541] <= 32'b00000100100000000000000011101111;
ROM[33542] <= 32'b00000000000000000000001110010011;
ROM[33543] <= 32'b00000000011100010010000000100011;
ROM[33544] <= 32'b00000000010000010000000100010011;
ROM[33545] <= 32'b00000001010000000000001110010011;
ROM[33546] <= 32'b01000000011100011000001110110011;
ROM[33547] <= 32'b00000000000000111010000010000011;
ROM[33548] <= 32'b11111111110000010000000100010011;
ROM[33549] <= 32'b00000000000000010010001110000011;
ROM[33550] <= 32'b00000000011100100010000000100011;
ROM[33551] <= 32'b00000000010000100000000100010011;
ROM[33552] <= 32'b00000001010000000000001110010011;
ROM[33553] <= 32'b01000000011100011000001110110011;
ROM[33554] <= 32'b00000000010000111010000110000011;
ROM[33555] <= 32'b00000000100000111010001000000011;
ROM[33556] <= 32'b00000000110000111010001010000011;
ROM[33557] <= 32'b00000001000000111010001100000011;
ROM[33558] <= 32'b00000000000000001000000011100111;
ROM[33559] <= 32'b00000000110100101000010000110011;
ROM[33560] <= 32'b00000001100001000010001110000011;
ROM[33561] <= 32'b00000000011100010010000000100011;
ROM[33562] <= 32'b00000000010000010000000100010011;
ROM[33563] <= 32'b00000000001100000000001110010011;
ROM[33564] <= 32'b00000000011100010010000000100011;
ROM[33565] <= 32'b00000000010000010000000100010011;
ROM[33566] <= 32'b11111111110000010000000100010011;
ROM[33567] <= 32'b00000000000000010010001110000011;
ROM[33568] <= 32'b11111111110000010000000100010011;
ROM[33569] <= 32'b00000000000000010010010000000011;
ROM[33570] <= 32'b00000000011101000010010010110011;
ROM[33571] <= 32'b00000000100000111010010100110011;
ROM[33572] <= 32'b00000000101001001000001110110011;
ROM[33573] <= 32'b00000000000100111000001110010011;
ROM[33574] <= 32'b00000000000100111111001110010011;
ROM[33575] <= 32'b00000000011100010010000000100011;
ROM[33576] <= 32'b00000000010000010000000100010011;
ROM[33577] <= 32'b11111111110000010000000100010011;
ROM[33578] <= 32'b00000000000000010010001110000011;
ROM[33579] <= 32'b00000000000000111000101001100011;
ROM[33580] <= 32'b00000000000000100001001110110111;
ROM[33581] <= 32'b11001100010000111000001110010011;
ROM[33582] <= 32'b00000000111000111000001110110011;
ROM[33583] <= 32'b00000000000000111000000011100111;
ROM[33584] <= 32'b00001111100000000000000011101111;
ROM[33585] <= 32'b00000000110100101000010000110011;
ROM[33586] <= 32'b00000000010001000010001110000011;
ROM[33587] <= 32'b00000000011100010010000000100011;
ROM[33588] <= 32'b00000000010000010000000100010011;
ROM[33589] <= 32'b00000000000000000000001110010011;
ROM[33590] <= 32'b00000000011100010010000000100011;
ROM[33591] <= 32'b00000000010000010000000100010011;
ROM[33592] <= 32'b11111111110000010000000100010011;
ROM[33593] <= 32'b00000000000000010010001110000011;
ROM[33594] <= 32'b11111111110000010000000100010011;
ROM[33595] <= 32'b00000000000000010010010000000011;
ROM[33596] <= 32'b00000000011101000010010010110011;
ROM[33597] <= 32'b00000000100000111010010100110011;
ROM[33598] <= 32'b00000000101001001000001110110011;
ROM[33599] <= 32'b00000000000100111000001110010011;
ROM[33600] <= 32'b00000000000100111111001110010011;
ROM[33601] <= 32'b00000000011100010010000000100011;
ROM[33602] <= 32'b00000000010000010000000100010011;
ROM[33603] <= 32'b11111111110000010000000100010011;
ROM[33604] <= 32'b00000000000000010010001110000011;
ROM[33605] <= 32'b00000000000000111000101001100011;
ROM[33606] <= 32'b00000000000000100001001110110111;
ROM[33607] <= 32'b11010111010000111000001110010011;
ROM[33608] <= 32'b00000000111000111000001110110011;
ROM[33609] <= 32'b00000000000000111000000011100111;
ROM[33610] <= 32'b00000000110100101000010000110011;
ROM[33611] <= 32'b00000000010001000010001110000011;
ROM[33612] <= 32'b00000000011100010010000000100011;
ROM[33613] <= 32'b00000000010000010000000100010011;
ROM[33614] <= 32'b00000000000100000000001110010011;
ROM[33615] <= 32'b00000000011100010010000000100011;
ROM[33616] <= 32'b00000000010000010000000100010011;
ROM[33617] <= 32'b11111111110000010000000100010011;
ROM[33618] <= 32'b00000000000000010010001110000011;
ROM[33619] <= 32'b11111111110000010000000100010011;
ROM[33620] <= 32'b00000000000000010010010000000011;
ROM[33621] <= 32'b01000000011101000000001110110011;
ROM[33622] <= 32'b00000000011100010010000000100011;
ROM[33623] <= 32'b00000000010000010000000100010011;
ROM[33624] <= 32'b11111111110000010000000100010011;
ROM[33625] <= 32'b00000000000000010010001110000011;
ROM[33626] <= 32'b00000000110100101000010000110011;
ROM[33627] <= 32'b00000000011101000010001000100011;
ROM[33628] <= 32'b00000100100000000000000011101111;
ROM[33629] <= 32'b00000000000000000000001110010011;
ROM[33630] <= 32'b00000000011100010010000000100011;
ROM[33631] <= 32'b00000000010000010000000100010011;
ROM[33632] <= 32'b00000001010000000000001110010011;
ROM[33633] <= 32'b01000000011100011000001110110011;
ROM[33634] <= 32'b00000000000000111010000010000011;
ROM[33635] <= 32'b11111111110000010000000100010011;
ROM[33636] <= 32'b00000000000000010010001110000011;
ROM[33637] <= 32'b00000000011100100010000000100011;
ROM[33638] <= 32'b00000000010000100000000100010011;
ROM[33639] <= 32'b00000001010000000000001110010011;
ROM[33640] <= 32'b01000000011100011000001110110011;
ROM[33641] <= 32'b00000000010000111010000110000011;
ROM[33642] <= 32'b00000000100000111010001000000011;
ROM[33643] <= 32'b00000000110000111010001010000011;
ROM[33644] <= 32'b00000001000000111010001100000011;
ROM[33645] <= 32'b00000000000000001000000011100111;
ROM[33646] <= 32'b00000000110100101000010000110011;
ROM[33647] <= 32'b00000001100001000010001110000011;
ROM[33648] <= 32'b00000000011100010010000000100011;
ROM[33649] <= 32'b00000000010000010000000100010011;
ROM[33650] <= 32'b00000000010000000000001110010011;
ROM[33651] <= 32'b00000000011100010010000000100011;
ROM[33652] <= 32'b00000000010000010000000100010011;
ROM[33653] <= 32'b11111111110000010000000100010011;
ROM[33654] <= 32'b00000000000000010010001110000011;
ROM[33655] <= 32'b11111111110000010000000100010011;
ROM[33656] <= 32'b00000000000000010010010000000011;
ROM[33657] <= 32'b00000000011101000010010010110011;
ROM[33658] <= 32'b00000000100000111010010100110011;
ROM[33659] <= 32'b00000000101001001000001110110011;
ROM[33660] <= 32'b00000000000100111000001110010011;
ROM[33661] <= 32'b00000000000100111111001110010011;
ROM[33662] <= 32'b00000000011100010010000000100011;
ROM[33663] <= 32'b00000000010000010000000100010011;
ROM[33664] <= 32'b11111111110000010000000100010011;
ROM[33665] <= 32'b00000000000000010010001110000011;
ROM[33666] <= 32'b00000000000000111000101001100011;
ROM[33667] <= 32'b00000000000000100001001110110111;
ROM[33668] <= 32'b11100010000000111000001110010011;
ROM[33669] <= 32'b00000000111000111000001110110011;
ROM[33670] <= 32'b00000000000000111000000011100111;
ROM[33671] <= 32'b00010100010000000000000011101111;
ROM[33672] <= 32'b00000000110100101000010000110011;
ROM[33673] <= 32'b00000000010001000010001110000011;
ROM[33674] <= 32'b00000000011100010010000000100011;
ROM[33675] <= 32'b00000000010000010000000100010011;
ROM[33676] <= 32'b00000000000000011010001110000011;
ROM[33677] <= 32'b00000000011100010010000000100011;
ROM[33678] <= 32'b00000000010000010000000100010011;
ROM[33679] <= 32'b00000000000000100001001110110111;
ROM[33680] <= 32'b11101000100000111000001110010011;
ROM[33681] <= 32'b00000000111000111000001110110011;
ROM[33682] <= 32'b00000000011100010010000000100011;
ROM[33683] <= 32'b00000000010000010000000100010011;
ROM[33684] <= 32'b00000000001100010010000000100011;
ROM[33685] <= 32'b00000000010000010000000100010011;
ROM[33686] <= 32'b00000000010000010010000000100011;
ROM[33687] <= 32'b00000000010000010000000100010011;
ROM[33688] <= 32'b00000000010100010010000000100011;
ROM[33689] <= 32'b00000000010000010000000100010011;
ROM[33690] <= 32'b00000000011000010010000000100011;
ROM[33691] <= 32'b00000000010000010000000100010011;
ROM[33692] <= 32'b00000001010000000000001110010011;
ROM[33693] <= 32'b00000000010000111000001110010011;
ROM[33694] <= 32'b01000000011100010000001110110011;
ROM[33695] <= 32'b00000000011100000000001000110011;
ROM[33696] <= 32'b00000000001000000000000110110011;
ROM[33697] <= 32'b00010001010000000101000011101111;
ROM[33698] <= 32'b11111111110000010000000100010011;
ROM[33699] <= 32'b00000000000000010010001110000011;
ROM[33700] <= 32'b11111111110000010000000100010011;
ROM[33701] <= 32'b00000000000000010010010000000011;
ROM[33702] <= 32'b00000000011101000010010010110011;
ROM[33703] <= 32'b00000000100000111010010100110011;
ROM[33704] <= 32'b00000000101001001000001110110011;
ROM[33705] <= 32'b00000000000100111000001110010011;
ROM[33706] <= 32'b00000000000100111111001110010011;
ROM[33707] <= 32'b00000000011100010010000000100011;
ROM[33708] <= 32'b00000000010000010000000100010011;
ROM[33709] <= 32'b11111111110000010000000100010011;
ROM[33710] <= 32'b00000000000000010010001110000011;
ROM[33711] <= 32'b00000000000000111000101001100011;
ROM[33712] <= 32'b00000000000000100001001110110111;
ROM[33713] <= 32'b11110001110000111000001110010011;
ROM[33714] <= 32'b00000000111000111000001110110011;
ROM[33715] <= 32'b00000000000000111000000011100111;
ROM[33716] <= 32'b00000000110100101000010000110011;
ROM[33717] <= 32'b00000000010001000010001110000011;
ROM[33718] <= 32'b00000000011100010010000000100011;
ROM[33719] <= 32'b00000000010000010000000100010011;
ROM[33720] <= 32'b00000000000100000000001110010011;
ROM[33721] <= 32'b00000000011100010010000000100011;
ROM[33722] <= 32'b00000000010000010000000100010011;
ROM[33723] <= 32'b11111111110000010000000100010011;
ROM[33724] <= 32'b00000000000000010010001110000011;
ROM[33725] <= 32'b11111111110000010000000100010011;
ROM[33726] <= 32'b00000000000000010010010000000011;
ROM[33727] <= 32'b00000000011101000000001110110011;
ROM[33728] <= 32'b00000000011100010010000000100011;
ROM[33729] <= 32'b00000000010000010000000100010011;
ROM[33730] <= 32'b11111111110000010000000100010011;
ROM[33731] <= 32'b00000000000000010010001110000011;
ROM[33732] <= 32'b00000000110100101000010000110011;
ROM[33733] <= 32'b00000000011101000010001000100011;
ROM[33734] <= 32'b00000100100000000000000011101111;
ROM[33735] <= 32'b00000000000000000000001110010011;
ROM[33736] <= 32'b00000000011100010010000000100011;
ROM[33737] <= 32'b00000000010000010000000100010011;
ROM[33738] <= 32'b00000001010000000000001110010011;
ROM[33739] <= 32'b01000000011100011000001110110011;
ROM[33740] <= 32'b00000000000000111010000010000011;
ROM[33741] <= 32'b11111111110000010000000100010011;
ROM[33742] <= 32'b00000000000000010010001110000011;
ROM[33743] <= 32'b00000000011100100010000000100011;
ROM[33744] <= 32'b00000000010000100000000100010011;
ROM[33745] <= 32'b00000001010000000000001110010011;
ROM[33746] <= 32'b01000000011100011000001110110011;
ROM[33747] <= 32'b00000000010000111010000110000011;
ROM[33748] <= 32'b00000000100000111010001000000011;
ROM[33749] <= 32'b00000000110000111010001010000011;
ROM[33750] <= 32'b00000001000000111010001100000011;
ROM[33751] <= 32'b00000000000000001000000011100111;
ROM[33752] <= 32'b00000000000000011010001110000011;
ROM[33753] <= 32'b00000000011100010010000000100011;
ROM[33754] <= 32'b00000000010000010000000100010011;
ROM[33755] <= 32'b00000000110100101000010000110011;
ROM[33756] <= 32'b00000000010001000010001110000011;
ROM[33757] <= 32'b00000000011100010010000000100011;
ROM[33758] <= 32'b00000000010000010000000100010011;
ROM[33759] <= 32'b00000000110100101000010000110011;
ROM[33760] <= 32'b00000000100001000010001110000011;
ROM[33761] <= 32'b00000000011100010010000000100011;
ROM[33762] <= 32'b00000000010000010000000100010011;
ROM[33763] <= 32'b00000000000000100001001110110111;
ROM[33764] <= 32'b11111101100000111000001110010011;
ROM[33765] <= 32'b00000000111000111000001110110011;
ROM[33766] <= 32'b00000000011100010010000000100011;
ROM[33767] <= 32'b00000000010000010000000100010011;
ROM[33768] <= 32'b00000000001100010010000000100011;
ROM[33769] <= 32'b00000000010000010000000100010011;
ROM[33770] <= 32'b00000000010000010010000000100011;
ROM[33771] <= 32'b00000000010000010000000100010011;
ROM[33772] <= 32'b00000000010100010010000000100011;
ROM[33773] <= 32'b00000000010000010000000100010011;
ROM[33774] <= 32'b00000000011000010010000000100011;
ROM[33775] <= 32'b00000000010000010000000100010011;
ROM[33776] <= 32'b00000001010000000000001110010011;
ROM[33777] <= 32'b00000000110000111000001110010011;
ROM[33778] <= 32'b01000000011100010000001110110011;
ROM[33779] <= 32'b00000000011100000000001000110011;
ROM[33780] <= 32'b00000000001000000000000110110011;
ROM[33781] <= 32'b00110001010000000101000011101111;
ROM[33782] <= 32'b11111111110000010000000100010011;
ROM[33783] <= 32'b00000000000000010010001110000011;
ROM[33784] <= 32'b00000000000000111000101001100011;
ROM[33785] <= 32'b00000000000000100001001110110111;
ROM[33786] <= 32'b11111111100000111000001110010011;
ROM[33787] <= 32'b00000000111000111000001110110011;
ROM[33788] <= 32'b00000000000000111000000011100111;
ROM[33789] <= 32'b00000100100000000000000011101111;
ROM[33790] <= 32'b00000000000000000000001110010011;
ROM[33791] <= 32'b00000000011100010010000000100011;
ROM[33792] <= 32'b00000000010000010000000100010011;
ROM[33793] <= 32'b00000001010000000000001110010011;
ROM[33794] <= 32'b01000000011100011000001110110011;
ROM[33795] <= 32'b00000000000000111010000010000011;
ROM[33796] <= 32'b11111111110000010000000100010011;
ROM[33797] <= 32'b00000000000000010010001110000011;
ROM[33798] <= 32'b00000000011100100010000000100011;
ROM[33799] <= 32'b00000000010000100000000100010011;
ROM[33800] <= 32'b00000001010000000000001110010011;
ROM[33801] <= 32'b01000000011100011000001110110011;
ROM[33802] <= 32'b00000000010000111010000110000011;
ROM[33803] <= 32'b00000000100000111010001000000011;
ROM[33804] <= 32'b00000000110000111010001010000011;
ROM[33805] <= 32'b00000001000000111010001100000011;
ROM[33806] <= 32'b00000000000000001000000011100111;
ROM[33807] <= 32'b00000000000100000000001110010011;
ROM[33808] <= 32'b00000000011100010010000000100011;
ROM[33809] <= 32'b00000000010000010000000100010011;
ROM[33810] <= 32'b11111111110000010000000100010011;
ROM[33811] <= 32'b00000000000000010010001110000011;
ROM[33812] <= 32'b01000000011100000000001110110011;
ROM[33813] <= 32'b00000000011100010010000000100011;
ROM[33814] <= 32'b00000000010000010000000100010011;
ROM[33815] <= 32'b00000001010000000000001110010011;
ROM[33816] <= 32'b01000000011100011000001110110011;
ROM[33817] <= 32'b00000000000000111010000010000011;
ROM[33818] <= 32'b11111111110000010000000100010011;
ROM[33819] <= 32'b00000000000000010010001110000011;
ROM[33820] <= 32'b00000000011100100010000000100011;
ROM[33821] <= 32'b00000000010000100000000100010011;
ROM[33822] <= 32'b00000001010000000000001110010011;
ROM[33823] <= 32'b01000000011100011000001110110011;
ROM[33824] <= 32'b00000000010000111010000110000011;
ROM[33825] <= 32'b00000000100000111010001000000011;
ROM[33826] <= 32'b00000000110000111010001010000011;
ROM[33827] <= 32'b00000001000000111010001100000011;
ROM[33828] <= 32'b00000000000000001000000011100111;
ROM[33829] <= 32'b00000000000000100010001110000011;
ROM[33830] <= 32'b00000000011100010010000000100011;
ROM[33831] <= 32'b00000000010000010000000100010011;
ROM[33832] <= 32'b11111111110000010000000100010011;
ROM[33833] <= 32'b00000000000000010010001110000011;
ROM[33834] <= 32'b00000000000000111000001010010011;
ROM[33835] <= 32'b00000000010100010010000000100011;
ROM[33836] <= 32'b00000000010000010000000100010011;
ROM[33837] <= 32'b00000000010000100010001110000011;
ROM[33838] <= 32'b00000000011100010010000000100011;
ROM[33839] <= 32'b00000000010000010000000100010011;
ROM[33840] <= 32'b00000000000000100001001110110111;
ROM[33841] <= 32'b00010000110000111000001110010011;
ROM[33842] <= 32'b00000000111000111000001110110011;
ROM[33843] <= 32'b00000000011100010010000000100011;
ROM[33844] <= 32'b00000000010000010000000100010011;
ROM[33845] <= 32'b00000000001100010010000000100011;
ROM[33846] <= 32'b00000000010000010000000100010011;
ROM[33847] <= 32'b00000000010000010010000000100011;
ROM[33848] <= 32'b00000000010000010000000100010011;
ROM[33849] <= 32'b00000000010100010010000000100011;
ROM[33850] <= 32'b00000000010000010000000100010011;
ROM[33851] <= 32'b00000000011000010010000000100011;
ROM[33852] <= 32'b00000000010000010000000100010011;
ROM[33853] <= 32'b00000001010000000000001110010011;
ROM[33854] <= 32'b00000000100000111000001110010011;
ROM[33855] <= 32'b01000000011100010000001110110011;
ROM[33856] <= 32'b00000000011100000000001000110011;
ROM[33857] <= 32'b00000000001000000000000110110011;
ROM[33858] <= 32'b00011010100000000000000011101111;
ROM[33859] <= 32'b11111111110000010000000100010011;
ROM[33860] <= 32'b00000000000000010010001110000011;
ROM[33861] <= 32'b00000000011101100010000000100011;
ROM[33862] <= 32'b00000000110100101000010000110011;
ROM[33863] <= 32'b00000001010001000010001110000011;
ROM[33864] <= 32'b00000000011100010010000000100011;
ROM[33865] <= 32'b00000000010000010000000100010011;
ROM[33866] <= 32'b00000000000000000000001110010011;
ROM[33867] <= 32'b00000000011100010010000000100011;
ROM[33868] <= 32'b00000000010000010000000100010011;
ROM[33869] <= 32'b11111111110000010000000100010011;
ROM[33870] <= 32'b00000000000000010010001110000011;
ROM[33871] <= 32'b11111111110000010000000100010011;
ROM[33872] <= 32'b00000000000000010010010000000011;
ROM[33873] <= 32'b00000000100000111010001110110011;
ROM[33874] <= 32'b00000000011100010010000000100011;
ROM[33875] <= 32'b00000000010000010000000100010011;
ROM[33876] <= 32'b11111111110000010000000100010011;
ROM[33877] <= 32'b00000000000000010010001110000011;
ROM[33878] <= 32'b00000000000000111000101001100011;
ROM[33879] <= 32'b00000000000000100001001110110111;
ROM[33880] <= 32'b00011101110000111000001110010011;
ROM[33881] <= 32'b00000000111000111000001110110011;
ROM[33882] <= 32'b00000000000000111000000011100111;
ROM[33883] <= 32'b00000000010100010010000000100011;
ROM[33884] <= 32'b00000000010000010000000100010011;
ROM[33885] <= 32'b00000000010000100010001110000011;
ROM[33886] <= 32'b00000000011100010010000000100011;
ROM[33887] <= 32'b00000000010000010000000100010011;
ROM[33888] <= 32'b00000000000000100001001110110111;
ROM[33889] <= 32'b00011100110000111000001110010011;
ROM[33890] <= 32'b00000000111000111000001110110011;
ROM[33891] <= 32'b00000000011100010010000000100011;
ROM[33892] <= 32'b00000000010000010000000100010011;
ROM[33893] <= 32'b00000000001100010010000000100011;
ROM[33894] <= 32'b00000000010000010000000100010011;
ROM[33895] <= 32'b00000000010000010010000000100011;
ROM[33896] <= 32'b00000000010000010000000100010011;
ROM[33897] <= 32'b00000000010100010010000000100011;
ROM[33898] <= 32'b00000000010000010000000100010011;
ROM[33899] <= 32'b00000000011000010010000000100011;
ROM[33900] <= 32'b00000000010000010000000100010011;
ROM[33901] <= 32'b00000001010000000000001110010011;
ROM[33902] <= 32'b00000000100000111000001110010011;
ROM[33903] <= 32'b01000000011100010000001110110011;
ROM[33904] <= 32'b00000000011100000000001000110011;
ROM[33905] <= 32'b00000000001000000000000110110011;
ROM[33906] <= 32'b00111011000000000000000011101111;
ROM[33907] <= 32'b11111111110000010000000100010011;
ROM[33908] <= 32'b00000000000000010010001110000011;
ROM[33909] <= 32'b00000000011101100010000000100011;
ROM[33910] <= 32'b00001001010000000000000011101111;
ROM[33911] <= 32'b00000000110100101000010000110011;
ROM[33912] <= 32'b00000001010001000010001110000011;
ROM[33913] <= 32'b00000000011100010010000000100011;
ROM[33914] <= 32'b00000000010000010000000100010011;
ROM[33915] <= 32'b00000000000100000000001110010011;
ROM[33916] <= 32'b00000000011100010010000000100011;
ROM[33917] <= 32'b00000000010000010000000100010011;
ROM[33918] <= 32'b11111111110000010000000100010011;
ROM[33919] <= 32'b00000000000000010010001110000011;
ROM[33920] <= 32'b11111111110000010000000100010011;
ROM[33921] <= 32'b00000000000000010010010000000011;
ROM[33922] <= 32'b01000000011101000000001110110011;
ROM[33923] <= 32'b00000000011100010010000000100011;
ROM[33924] <= 32'b00000000010000010000000100010011;
ROM[33925] <= 32'b11111111110000010000000100010011;
ROM[33926] <= 32'b00000000000000010010001110000011;
ROM[33927] <= 32'b00000000110100101000010000110011;
ROM[33928] <= 32'b00000000011101000010101000100011;
ROM[33929] <= 32'b00000000110100101000010000110011;
ROM[33930] <= 32'b00000000110001000010001110000011;
ROM[33931] <= 32'b00000000011100010010000000100011;
ROM[33932] <= 32'b00000000010000010000000100010011;
ROM[33933] <= 32'b00000000000100000000001110010011;
ROM[33934] <= 32'b00000000011100010010000000100011;
ROM[33935] <= 32'b00000000010000010000000100010011;
ROM[33936] <= 32'b11111111110000010000000100010011;
ROM[33937] <= 32'b00000000000000010010001110000011;
ROM[33938] <= 32'b11111111110000010000000100010011;
ROM[33939] <= 32'b00000000000000010010010000000011;
ROM[33940] <= 32'b00000000011101000000001110110011;
ROM[33941] <= 32'b00000000011100010010000000100011;
ROM[33942] <= 32'b00000000010000010000000100010011;
ROM[33943] <= 32'b11111111110000010000000100010011;
ROM[33944] <= 32'b00000000000000010010001110000011;
ROM[33945] <= 32'b00000000110100101000010000110011;
ROM[33946] <= 32'b00000000011101000010011000100011;
ROM[33947] <= 32'b00000000000000000000001110010011;
ROM[33948] <= 32'b00000000011100010010000000100011;
ROM[33949] <= 32'b00000000010000010000000100010011;
ROM[33950] <= 32'b00000001010000000000001110010011;
ROM[33951] <= 32'b01000000011100011000001110110011;
ROM[33952] <= 32'b00000000000000111010000010000011;
ROM[33953] <= 32'b11111111110000010000000100010011;
ROM[33954] <= 32'b00000000000000010010001110000011;
ROM[33955] <= 32'b00000000011100100010000000100011;
ROM[33956] <= 32'b00000000010000100000000100010011;
ROM[33957] <= 32'b00000001010000000000001110010011;
ROM[33958] <= 32'b01000000011100011000001110110011;
ROM[33959] <= 32'b00000000010000111010000110000011;
ROM[33960] <= 32'b00000000100000111010001000000011;
ROM[33961] <= 32'b00000000110000111010001010000011;
ROM[33962] <= 32'b00000001000000111010001100000011;
ROM[33963] <= 32'b00000000000000001000000011100111;
ROM[33964] <= 32'b00000000000000010010000000100011;
ROM[33965] <= 32'b00000000010000010000000100010011;
ROM[33966] <= 32'b00000000000000100010001110000011;
ROM[33967] <= 32'b00000000011100010010000000100011;
ROM[33968] <= 32'b00000000010000010000000100010011;
ROM[33969] <= 32'b11111111110000010000000100010011;
ROM[33970] <= 32'b00000000000000010010001110000011;
ROM[33971] <= 32'b00000000000000111000001010010011;
ROM[33972] <= 32'b00000000110100101000010000110011;
ROM[33973] <= 32'b00000000000001000010001110000011;
ROM[33974] <= 32'b00000000011100010010000000100011;
ROM[33975] <= 32'b00000000010000010000000100010011;
ROM[33976] <= 32'b00000000000000100001001110110111;
ROM[33977] <= 32'b00110010110000111000001110010011;
ROM[33978] <= 32'b00000000111000111000001110110011;
ROM[33979] <= 32'b00000000011100010010000000100011;
ROM[33980] <= 32'b00000000010000010000000100010011;
ROM[33981] <= 32'b00000000001100010010000000100011;
ROM[33982] <= 32'b00000000010000010000000100010011;
ROM[33983] <= 32'b00000000010000010010000000100011;
ROM[33984] <= 32'b00000000010000010000000100010011;
ROM[33985] <= 32'b00000000010100010010000000100011;
ROM[33986] <= 32'b00000000010000010000000100010011;
ROM[33987] <= 32'b00000000011000010010000000100011;
ROM[33988] <= 32'b00000000010000010000000100010011;
ROM[33989] <= 32'b00000001010000000000001110010011;
ROM[33990] <= 32'b00000000010000111000001110010011;
ROM[33991] <= 32'b01000000011100010000001110110011;
ROM[33992] <= 32'b00000000011100000000001000110011;
ROM[33993] <= 32'b00000000001000000000000110110011;
ROM[33994] <= 32'b01110011110000000010000011101111;
ROM[33995] <= 32'b11111111110000010000000100010011;
ROM[33996] <= 32'b00000000000000010010001110000011;
ROM[33997] <= 32'b00000000011100011010000000100011;
ROM[33998] <= 32'b00000000000000011010001110000011;
ROM[33999] <= 32'b00000000011100010010000000100011;
ROM[34000] <= 32'b00000000010000010000000100010011;
ROM[34001] <= 32'b00000000110100101000010000110011;
ROM[34002] <= 32'b00000000010001000010001110000011;
ROM[34003] <= 32'b00000000011100010010000000100011;
ROM[34004] <= 32'b00000000010000010000000100010011;
ROM[34005] <= 32'b00000000110100101000010000110011;
ROM[34006] <= 32'b00000000100001000010001110000011;
ROM[34007] <= 32'b00000000011100010010000000100011;
ROM[34008] <= 32'b00000000010000010000000100010011;
ROM[34009] <= 32'b00000000000000100001001110110111;
ROM[34010] <= 32'b00111011000000111000001110010011;
ROM[34011] <= 32'b00000000111000111000001110110011;
ROM[34012] <= 32'b00000000011100010010000000100011;
ROM[34013] <= 32'b00000000010000010000000100010011;
ROM[34014] <= 32'b00000000001100010010000000100011;
ROM[34015] <= 32'b00000000010000010000000100010011;
ROM[34016] <= 32'b00000000010000010010000000100011;
ROM[34017] <= 32'b00000000010000010000000100010011;
ROM[34018] <= 32'b00000000010100010010000000100011;
ROM[34019] <= 32'b00000000010000010000000100010011;
ROM[34020] <= 32'b00000000011000010010000000100011;
ROM[34021] <= 32'b00000000010000010000000100010011;
ROM[34022] <= 32'b00000001010000000000001110010011;
ROM[34023] <= 32'b00000000110000111000001110010011;
ROM[34024] <= 32'b01000000011100010000001110110011;
ROM[34025] <= 32'b00000000011100000000001000110011;
ROM[34026] <= 32'b00000000001000000000000110110011;
ROM[34027] <= 32'b01100010010000000101000011101111;
ROM[34028] <= 32'b11111111110000010000000100010011;
ROM[34029] <= 32'b00000000000000010010001110000011;
ROM[34030] <= 32'b00000000011101100010000000100011;
ROM[34031] <= 32'b00000000110100101000010000110011;
ROM[34032] <= 32'b00000000010001000010001110000011;
ROM[34033] <= 32'b00000000011100010010000000100011;
ROM[34034] <= 32'b00000000010000010000000100010011;
ROM[34035] <= 32'b00000000110100101000010000110011;
ROM[34036] <= 32'b00000010000001000010001110000011;
ROM[34037] <= 32'b00000000011100010010000000100011;
ROM[34038] <= 32'b00000000010000010000000100010011;
ROM[34039] <= 32'b00000000010000100010001110000011;
ROM[34040] <= 32'b00000000011100010010000000100011;
ROM[34041] <= 32'b00000000010000010000000100010011;
ROM[34042] <= 32'b00000000010000000000001110010011;
ROM[34043] <= 32'b00000000011100010010000000100011;
ROM[34044] <= 32'b00000000010000010000000100010011;
ROM[34045] <= 32'b00000000000000100001001110110111;
ROM[34046] <= 32'b01000100000000111000001110010011;
ROM[34047] <= 32'b00000000111000111000001110110011;
ROM[34048] <= 32'b00000000011100010010000000100011;
ROM[34049] <= 32'b00000000010000010000000100010011;
ROM[34050] <= 32'b00000000001100010010000000100011;
ROM[34051] <= 32'b00000000010000010000000100010011;
ROM[34052] <= 32'b00000000010000010010000000100011;
ROM[34053] <= 32'b00000000010000010000000100010011;
ROM[34054] <= 32'b00000000010100010010000000100011;
ROM[34055] <= 32'b00000000010000010000000100010011;
ROM[34056] <= 32'b00000000011000010010000000100011;
ROM[34057] <= 32'b00000000010000010000000100010011;
ROM[34058] <= 32'b00000001010000000000001110010011;
ROM[34059] <= 32'b00000000100000111000001110010011;
ROM[34060] <= 32'b01000000011100010000001110110011;
ROM[34061] <= 32'b00000000011100000000001000110011;
ROM[34062] <= 32'b00000000001000000000000110110011;
ROM[34063] <= 32'b10111111000011110000000011101111;
ROM[34064] <= 32'b11111111110000010000000100010011;
ROM[34065] <= 32'b00000000000000010010001110000011;
ROM[34066] <= 32'b11111111110000010000000100010011;
ROM[34067] <= 32'b00000000000000010010010000000011;
ROM[34068] <= 32'b00000000011101000000001110110011;
ROM[34069] <= 32'b00000000011100010010000000100011;
ROM[34070] <= 32'b00000000010000010000000100010011;
ROM[34071] <= 32'b11111111110000010000000100010011;
ROM[34072] <= 32'b00000000000000010010001110000011;
ROM[34073] <= 32'b00000000000000111000001100010011;
ROM[34074] <= 32'b11111111110000010000000100010011;
ROM[34075] <= 32'b00000000000000010010001110000011;
ROM[34076] <= 32'b00000000110100110000010000110011;
ROM[34077] <= 32'b00000000011101000010000000100011;
ROM[34078] <= 32'b00000000110100101000010000110011;
ROM[34079] <= 32'b00000000100001000010001110000011;
ROM[34080] <= 32'b00000000011100010010000000100011;
ROM[34081] <= 32'b00000000010000010000000100010011;
ROM[34082] <= 32'b00000000110100101000010000110011;
ROM[34083] <= 32'b00000010010001000010001110000011;
ROM[34084] <= 32'b00000000011100010010000000100011;
ROM[34085] <= 32'b00000000010000010000000100010011;
ROM[34086] <= 32'b00000000010000100010001110000011;
ROM[34087] <= 32'b00000000011100010010000000100011;
ROM[34088] <= 32'b00000000010000010000000100010011;
ROM[34089] <= 32'b00000000010000000000001110010011;
ROM[34090] <= 32'b00000000011100010010000000100011;
ROM[34091] <= 32'b00000000010000010000000100010011;
ROM[34092] <= 32'b00000000000000100001001110110111;
ROM[34093] <= 32'b01001111110000111000001110010011;
ROM[34094] <= 32'b00000000111000111000001110110011;
ROM[34095] <= 32'b00000000011100010010000000100011;
ROM[34096] <= 32'b00000000010000010000000100010011;
ROM[34097] <= 32'b00000000001100010010000000100011;
ROM[34098] <= 32'b00000000010000010000000100010011;
ROM[34099] <= 32'b00000000010000010010000000100011;
ROM[34100] <= 32'b00000000010000010000000100010011;
ROM[34101] <= 32'b00000000010100010010000000100011;
ROM[34102] <= 32'b00000000010000010000000100010011;
ROM[34103] <= 32'b00000000011000010010000000100011;
ROM[34104] <= 32'b00000000010000010000000100010011;
ROM[34105] <= 32'b00000001010000000000001110010011;
ROM[34106] <= 32'b00000000100000111000001110010011;
ROM[34107] <= 32'b01000000011100010000001110110011;
ROM[34108] <= 32'b00000000011100000000001000110011;
ROM[34109] <= 32'b00000000001000000000000110110011;
ROM[34110] <= 32'b10110011010011110000000011101111;
ROM[34111] <= 32'b11111111110000010000000100010011;
ROM[34112] <= 32'b00000000000000010010001110000011;
ROM[34113] <= 32'b11111111110000010000000100010011;
ROM[34114] <= 32'b00000000000000010010010000000011;
ROM[34115] <= 32'b00000000011101000000001110110011;
ROM[34116] <= 32'b00000000011100010010000000100011;
ROM[34117] <= 32'b00000000010000010000000100010011;
ROM[34118] <= 32'b11111111110000010000000100010011;
ROM[34119] <= 32'b00000000000000010010001110000011;
ROM[34120] <= 32'b00000000000000111000001100010011;
ROM[34121] <= 32'b11111111110000010000000100010011;
ROM[34122] <= 32'b00000000000000010010001110000011;
ROM[34123] <= 32'b00000000110100110000010000110011;
ROM[34124] <= 32'b00000000011101000010000000100011;
ROM[34125] <= 32'b00000000000000000000001110010011;
ROM[34126] <= 32'b00000000011100010010000000100011;
ROM[34127] <= 32'b00000000010000010000000100010011;
ROM[34128] <= 32'b00000001010000000000001110010011;
ROM[34129] <= 32'b01000000011100011000001110110011;
ROM[34130] <= 32'b00000000000000111010000010000011;
ROM[34131] <= 32'b11111111110000010000000100010011;
ROM[34132] <= 32'b00000000000000010010001110000011;
ROM[34133] <= 32'b00000000011100100010000000100011;
ROM[34134] <= 32'b00000000010000100000000100010011;
ROM[34135] <= 32'b00000001010000000000001110010011;
ROM[34136] <= 32'b01000000011100011000001110110011;
ROM[34137] <= 32'b00000000010000111010000110000011;
ROM[34138] <= 32'b00000000100000111010001000000011;
ROM[34139] <= 32'b00000000110000111010001010000011;
ROM[34140] <= 32'b00000001000000111010001100000011;
ROM[34141] <= 32'b00000000000000001000000011100111;
ROM[34142] <= 32'b00000000000000010010000000100011;
ROM[34143] <= 32'b00000000010000010000000100010011;
ROM[34144] <= 32'b00000000000000010010000000100011;
ROM[34145] <= 32'b00000000010000010000000100010011;
ROM[34146] <= 32'b00000000000000010010000000100011;
ROM[34147] <= 32'b00000000010000010000000100010011;
ROM[34148] <= 32'b00000000000000010010000000100011;
ROM[34149] <= 32'b00000000010000010000000100010011;
ROM[34150] <= 32'b00000000000000100010001110000011;
ROM[34151] <= 32'b00000000011100010010000000100011;
ROM[34152] <= 32'b00000000010000010000000100010011;
ROM[34153] <= 32'b11111111110000010000000100010011;
ROM[34154] <= 32'b00000000000000010010001110000011;
ROM[34155] <= 32'b00000000000000111000001010010011;
ROM[34156] <= 32'b00000000010000100010001110000011;
ROM[34157] <= 32'b00000000011100010010000000100011;
ROM[34158] <= 32'b00000000010000010000000100010011;
ROM[34159] <= 32'b00000000110100101000010000110011;
ROM[34160] <= 32'b00000000110001000010001110000011;
ROM[34161] <= 32'b00000000011100010010000000100011;
ROM[34162] <= 32'b00000000010000010000000100010011;
ROM[34163] <= 32'b11111111110000010000000100010011;
ROM[34164] <= 32'b00000000000000010010001110000011;
ROM[34165] <= 32'b11111111110000010000000100010011;
ROM[34166] <= 32'b00000000000000010010010000000011;
ROM[34167] <= 32'b01000000011101000000001110110011;
ROM[34168] <= 32'b00000000011100010010000000100011;
ROM[34169] <= 32'b00000000010000010000000100010011;
ROM[34170] <= 32'b11111111110000010000000100010011;
ROM[34171] <= 32'b00000000000000010010001110000011;
ROM[34172] <= 32'b00000000011100011010001000100011;
ROM[34173] <= 32'b00000000110100101000010000110011;
ROM[34174] <= 32'b00000010000001000010001110000011;
ROM[34175] <= 32'b00000000011100010010000000100011;
ROM[34176] <= 32'b00000000010000010000000100010011;
ROM[34177] <= 32'b00000000010000011010001110000011;
ROM[34178] <= 32'b00000000011100010010000000100011;
ROM[34179] <= 32'b00000000010000010000000100010011;
ROM[34180] <= 32'b00000000010000000000001110010011;
ROM[34181] <= 32'b00000000011100010010000000100011;
ROM[34182] <= 32'b00000000010000010000000100010011;
ROM[34183] <= 32'b00000000000000100001001110110111;
ROM[34184] <= 32'b01100110100000111000001110010011;
ROM[34185] <= 32'b00000000111000111000001110110011;
ROM[34186] <= 32'b00000000011100010010000000100011;
ROM[34187] <= 32'b00000000010000010000000100010011;
ROM[34188] <= 32'b00000000001100010010000000100011;
ROM[34189] <= 32'b00000000010000010000000100010011;
ROM[34190] <= 32'b00000000010000010010000000100011;
ROM[34191] <= 32'b00000000010000010000000100010011;
ROM[34192] <= 32'b00000000010100010010000000100011;
ROM[34193] <= 32'b00000000010000010000000100010011;
ROM[34194] <= 32'b00000000011000010010000000100011;
ROM[34195] <= 32'b00000000010000010000000100010011;
ROM[34196] <= 32'b00000001010000000000001110010011;
ROM[34197] <= 32'b00000000100000111000001110010011;
ROM[34198] <= 32'b01000000011100010000001110110011;
ROM[34199] <= 32'b00000000011100000000001000110011;
ROM[34200] <= 32'b00000000001000000000000110110011;
ROM[34201] <= 32'b10011100100011110000000011101111;
ROM[34202] <= 32'b11111111110000010000000100010011;
ROM[34203] <= 32'b00000000000000010010001110000011;
ROM[34204] <= 32'b11111111110000010000000100010011;
ROM[34205] <= 32'b00000000000000010010010000000011;
ROM[34206] <= 32'b00000000011101000000001110110011;
ROM[34207] <= 32'b00000000011100010010000000100011;
ROM[34208] <= 32'b00000000010000010000000100010011;
ROM[34209] <= 32'b11111111110000010000000100010011;
ROM[34210] <= 32'b00000000000000010010001110000011;
ROM[34211] <= 32'b00000000000000111000001100010011;
ROM[34212] <= 32'b00000000110100110000010000110011;
ROM[34213] <= 32'b00000000000001000010001110000011;
ROM[34214] <= 32'b00000000011100010010000000100011;
ROM[34215] <= 32'b00000000010000010000000100010011;
ROM[34216] <= 32'b11111111110000010000000100010011;
ROM[34217] <= 32'b00000000000000010010001110000011;
ROM[34218] <= 32'b00000000011100011010010000100011;
ROM[34219] <= 32'b00000000110100101000010000110011;
ROM[34220] <= 32'b00000010010001000010001110000011;
ROM[34221] <= 32'b00000000011100010010000000100011;
ROM[34222] <= 32'b00000000010000010000000100010011;
ROM[34223] <= 32'b00000000010000011010001110000011;
ROM[34224] <= 32'b00000000011100010010000000100011;
ROM[34225] <= 32'b00000000010000010000000100010011;
ROM[34226] <= 32'b00000000010000000000001110010011;
ROM[34227] <= 32'b00000000011100010010000000100011;
ROM[34228] <= 32'b00000000010000010000000100010011;
ROM[34229] <= 32'b00000000000000100001001110110111;
ROM[34230] <= 32'b01110010000000111000001110010011;
ROM[34231] <= 32'b00000000111000111000001110110011;
ROM[34232] <= 32'b00000000011100010010000000100011;
ROM[34233] <= 32'b00000000010000010000000100010011;
ROM[34234] <= 32'b00000000001100010010000000100011;
ROM[34235] <= 32'b00000000010000010000000100010011;
ROM[34236] <= 32'b00000000010000010010000000100011;
ROM[34237] <= 32'b00000000010000010000000100010011;
ROM[34238] <= 32'b00000000010100010010000000100011;
ROM[34239] <= 32'b00000000010000010000000100010011;
ROM[34240] <= 32'b00000000011000010010000000100011;
ROM[34241] <= 32'b00000000010000010000000100010011;
ROM[34242] <= 32'b00000001010000000000001110010011;
ROM[34243] <= 32'b00000000100000111000001110010011;
ROM[34244] <= 32'b01000000011100010000001110110011;
ROM[34245] <= 32'b00000000011100000000001000110011;
ROM[34246] <= 32'b00000000001000000000000110110011;
ROM[34247] <= 32'b10010001000011110000000011101111;
ROM[34248] <= 32'b11111111110000010000000100010011;
ROM[34249] <= 32'b00000000000000010010001110000011;
ROM[34250] <= 32'b11111111110000010000000100010011;
ROM[34251] <= 32'b00000000000000010010010000000011;
ROM[34252] <= 32'b00000000011101000000001110110011;
ROM[34253] <= 32'b00000000011100010010000000100011;
ROM[34254] <= 32'b00000000010000010000000100010011;
ROM[34255] <= 32'b11111111110000010000000100010011;
ROM[34256] <= 32'b00000000000000010010001110000011;
ROM[34257] <= 32'b00000000000000111000001100010011;
ROM[34258] <= 32'b00000000110100110000010000110011;
ROM[34259] <= 32'b00000000000001000010001110000011;
ROM[34260] <= 32'b00000000011100010010000000100011;
ROM[34261] <= 32'b00000000010000010000000100010011;
ROM[34262] <= 32'b11111111110000010000000100010011;
ROM[34263] <= 32'b00000000000000010010001110000011;
ROM[34264] <= 32'b00000000011100011010011000100011;
ROM[34265] <= 32'b00000000110100101000010000110011;
ROM[34266] <= 32'b00000000000001000010001110000011;
ROM[34267] <= 32'b00000000011100010010000000100011;
ROM[34268] <= 32'b00000000010000010000000100010011;
ROM[34269] <= 32'b00000000000000100001001110110111;
ROM[34270] <= 32'b01111100000000111000001110010011;
ROM[34271] <= 32'b00000000111000111000001110110011;
ROM[34272] <= 32'b00000000011100010010000000100011;
ROM[34273] <= 32'b00000000010000010000000100010011;
ROM[34274] <= 32'b00000000001100010010000000100011;
ROM[34275] <= 32'b00000000010000010000000100010011;
ROM[34276] <= 32'b00000000010000010010000000100011;
ROM[34277] <= 32'b00000000010000010000000100010011;
ROM[34278] <= 32'b00000000010100010010000000100011;
ROM[34279] <= 32'b00000000010000010000000100010011;
ROM[34280] <= 32'b00000000011000010010000000100011;
ROM[34281] <= 32'b00000000010000010000000100010011;
ROM[34282] <= 32'b00000001010000000000001110010011;
ROM[34283] <= 32'b00000000010000111000001110010011;
ROM[34284] <= 32'b01000000011100010000001110110011;
ROM[34285] <= 32'b00000000011100000000001000110011;
ROM[34286] <= 32'b00000000001000000000000110110011;
ROM[34287] <= 32'b00101010100000000010000011101111;
ROM[34288] <= 32'b11111111110000010000000100010011;
ROM[34289] <= 32'b00000000000000010010001110000011;
ROM[34290] <= 32'b00000000011100011010000000100011;
ROM[34291] <= 32'b00000000000000011010001110000011;
ROM[34292] <= 32'b00000000011100010010000000100011;
ROM[34293] <= 32'b00000000010000010000000100010011;
ROM[34294] <= 32'b00000000100000011010001110000011;
ROM[34295] <= 32'b00000000011100010010000000100011;
ROM[34296] <= 32'b00000000010000010000000100010011;
ROM[34297] <= 32'b00000000110000011010001110000011;
ROM[34298] <= 32'b00000000011100010010000000100011;
ROM[34299] <= 32'b00000000010000010000000100010011;
ROM[34300] <= 32'b00000000000000100010001110110111;
ROM[34301] <= 32'b10000011110000111000001110010011;
ROM[34302] <= 32'b00000000111000111000001110110011;
ROM[34303] <= 32'b00000000011100010010000000100011;
ROM[34304] <= 32'b00000000010000010000000100010011;
ROM[34305] <= 32'b00000000001100010010000000100011;
ROM[34306] <= 32'b00000000010000010000000100010011;
ROM[34307] <= 32'b00000000010000010010000000100011;
ROM[34308] <= 32'b00000000010000010000000100010011;
ROM[34309] <= 32'b00000000010100010010000000100011;
ROM[34310] <= 32'b00000000010000010000000100010011;
ROM[34311] <= 32'b00000000011000010010000000100011;
ROM[34312] <= 32'b00000000010000010000000100010011;
ROM[34313] <= 32'b00000001010000000000001110010011;
ROM[34314] <= 32'b00000000110000111000001110010011;
ROM[34315] <= 32'b01000000011100010000001110110011;
ROM[34316] <= 32'b00000000011100000000001000110011;
ROM[34317] <= 32'b00000000001000000000000110110011;
ROM[34318] <= 32'b01010011110000000101000011101111;
ROM[34319] <= 32'b11111111110000010000000100010011;
ROM[34320] <= 32'b00000000000000010010001110000011;
ROM[34321] <= 32'b00000000011101100010000000100011;
ROM[34322] <= 32'b00000000000000000000001110010011;
ROM[34323] <= 32'b00000000011100010010000000100011;
ROM[34324] <= 32'b00000000010000010000000100010011;
ROM[34325] <= 32'b00000001010000000000001110010011;
ROM[34326] <= 32'b01000000011100011000001110110011;
ROM[34327] <= 32'b00000000000000111010000010000011;
ROM[34328] <= 32'b11111111110000010000000100010011;
ROM[34329] <= 32'b00000000000000010010001110000011;
ROM[34330] <= 32'b00000000011100100010000000100011;
ROM[34331] <= 32'b00000000010000100000000100010011;
ROM[34332] <= 32'b00000001010000000000001110010011;
ROM[34333] <= 32'b01000000011100011000001110110011;
ROM[34334] <= 32'b00000000010000111010000110000011;
ROM[34335] <= 32'b00000000100000111010001000000011;
ROM[34336] <= 32'b00000000110000111010001010000011;
ROM[34337] <= 32'b00000001000000111010001100000011;
ROM[34338] <= 32'b00000000000000001000000011100111;
ROM[34339] <= 32'b00000000000000100010001110000011;
ROM[34340] <= 32'b00000000011100010010000000100011;
ROM[34341] <= 32'b00000000010000010000000100010011;
ROM[34342] <= 32'b11111111110000010000000100010011;
ROM[34343] <= 32'b00000000000000010010001110000011;
ROM[34344] <= 32'b00000000000000111000001010010011;
ROM[34345] <= 32'b00000000110100101000010000110011;
ROM[34346] <= 32'b00000001010001000010001110000011;
ROM[34347] <= 32'b00000000011100010010000000100011;
ROM[34348] <= 32'b00000000010000010000000100010011;
ROM[34349] <= 32'b00000000110100101000010000110011;
ROM[34350] <= 32'b00000001000001000010001110000011;
ROM[34351] <= 32'b00000000011100010010000000100011;
ROM[34352] <= 32'b00000000010000010000000100010011;
ROM[34353] <= 32'b11111111110000010000000100010011;
ROM[34354] <= 32'b00000000000000010010001110000011;
ROM[34355] <= 32'b11111111110000010000000100010011;
ROM[34356] <= 32'b00000000000000010010010000000011;
ROM[34357] <= 32'b00000000011101000000001110110011;
ROM[34358] <= 32'b00000000011100010010000000100011;
ROM[34359] <= 32'b00000000010000010000000100010011;
ROM[34360] <= 32'b11111111110000010000000100010011;
ROM[34361] <= 32'b00000000000000010010001110000011;
ROM[34362] <= 32'b00000000110100101000010000110011;
ROM[34363] <= 32'b00000000011101000010101000100011;
ROM[34364] <= 32'b00000000000000000000001110010011;
ROM[34365] <= 32'b00000000011100010010000000100011;
ROM[34366] <= 32'b00000000010000010000000100010011;
ROM[34367] <= 32'b00000001010000000000001110010011;
ROM[34368] <= 32'b01000000011100011000001110110011;
ROM[34369] <= 32'b00000000000000111010000010000011;
ROM[34370] <= 32'b11111111110000010000000100010011;
ROM[34371] <= 32'b00000000000000010010001110000011;
ROM[34372] <= 32'b00000000011100100010000000100011;
ROM[34373] <= 32'b00000000010000100000000100010011;
ROM[34374] <= 32'b00000001010000000000001110010011;
ROM[34375] <= 32'b01000000011100011000001110110011;
ROM[34376] <= 32'b00000000010000111010000110000011;
ROM[34377] <= 32'b00000000100000111010001000000011;
ROM[34378] <= 32'b00000000110000111010001010000011;
ROM[34379] <= 32'b00000001000000111010001100000011;
ROM[34380] <= 32'b00000000000000001000000011100111;
ROM[34381] <= 32'b00000000011100000000001110010011;
ROM[34382] <= 32'b00000000011100010010000000100011;
ROM[34383] <= 32'b00000000010000010000000100010011;
ROM[34384] <= 32'b00000000000000100010001110110111;
ROM[34385] <= 32'b10011000110000111000001110010011;
ROM[34386] <= 32'b00000000111000111000001110110011;
ROM[34387] <= 32'b00000000011100010010000000100011;
ROM[34388] <= 32'b00000000010000010000000100010011;
ROM[34389] <= 32'b00000000001100010010000000100011;
ROM[34390] <= 32'b00000000010000010000000100010011;
ROM[34391] <= 32'b00000000010000010010000000100011;
ROM[34392] <= 32'b00000000010000010000000100010011;
ROM[34393] <= 32'b00000000010100010010000000100011;
ROM[34394] <= 32'b00000000010000010000000100010011;
ROM[34395] <= 32'b00000000011000010010000000100011;
ROM[34396] <= 32'b00000000010000010000000100010011;
ROM[34397] <= 32'b00000001010000000000001110010011;
ROM[34398] <= 32'b00000000010000111000001110010011;
ROM[34399] <= 32'b01000000011100010000001110110011;
ROM[34400] <= 32'b00000000011100000000001000110011;
ROM[34401] <= 32'b00000000001000000000000110110011;
ROM[34402] <= 32'b11010100110111110010000011101111;
ROM[34403] <= 32'b11111111110000010000000100010011;
ROM[34404] <= 32'b00000000000000010010001110000011;
ROM[34405] <= 32'b00000000000000111000001010010011;
ROM[34406] <= 32'b00000000000000000000001110010011;
ROM[34407] <= 32'b00000000011100010010000000100011;
ROM[34408] <= 32'b00000000010000010000000100010011;
ROM[34409] <= 32'b11111111110000010000000100010011;
ROM[34410] <= 32'b00000000000000010010001110000011;
ROM[34411] <= 32'b00000000110100101000010000110011;
ROM[34412] <= 32'b00000000011101000010010000100011;
ROM[34413] <= 32'b00000000000100000000001110010011;
ROM[34414] <= 32'b00000000011100010010000000100011;
ROM[34415] <= 32'b00000000010000010000000100010011;
ROM[34416] <= 32'b11111111110000010000000100010011;
ROM[34417] <= 32'b00000000000000010010001110000011;
ROM[34418] <= 32'b00000000110100101000010000110011;
ROM[34419] <= 32'b00000000011101000010011000100011;
ROM[34420] <= 32'b00000000000000000000001110010011;
ROM[34421] <= 32'b00000000011100010010000000100011;
ROM[34422] <= 32'b00000000010000010000000100010011;
ROM[34423] <= 32'b11111111110000010000000100010011;
ROM[34424] <= 32'b00000000000000010010001110000011;
ROM[34425] <= 32'b00000000110100101000010000110011;
ROM[34426] <= 32'b00000000011101000010100000100011;
ROM[34427] <= 32'b00000000000000000000001110010011;
ROM[34428] <= 32'b00000000011100010010000000100011;
ROM[34429] <= 32'b00000000010000010000000100010011;
ROM[34430] <= 32'b11111111110000010000000100010011;
ROM[34431] <= 32'b00000000000000010010001110000011;
ROM[34432] <= 32'b00000000110100101000010000110011;
ROM[34433] <= 32'b00000000011101000010101000100011;
ROM[34434] <= 32'b00000110010000000000001110010011;
ROM[34435] <= 32'b00000000011100010010000000100011;
ROM[34436] <= 32'b00000000010000010000000100010011;
ROM[34437] <= 32'b11111111110000010000000100010011;
ROM[34438] <= 32'b00000000000000010010001110000011;
ROM[34439] <= 32'b00000000110100101000010000110011;
ROM[34440] <= 32'b00000000011101000010110000100011;
ROM[34441] <= 32'b00000000010100010010000000100011;
ROM[34442] <= 32'b00000000010000010000000100010011;
ROM[34443] <= 32'b00100000000000000000001110010011;
ROM[34444] <= 32'b00000000011100010010000000100011;
ROM[34445] <= 32'b00000000010000010000000100010011;
ROM[34446] <= 32'b00010000000000000000001110010011;
ROM[34447] <= 32'b00000000011100010010000000100011;
ROM[34448] <= 32'b00000000010000010000000100010011;
ROM[34449] <= 32'b00000000000000100010001110110111;
ROM[34450] <= 32'b10101001000000111000001110010011;
ROM[34451] <= 32'b00000000111000111000001110110011;
ROM[34452] <= 32'b00000000011100010010000000100011;
ROM[34453] <= 32'b00000000010000010000000100010011;
ROM[34454] <= 32'b00000000001100010010000000100011;
ROM[34455] <= 32'b00000000010000010000000100010011;
ROM[34456] <= 32'b00000000010000010010000000100011;
ROM[34457] <= 32'b00000000010000010000000100010011;
ROM[34458] <= 32'b00000000010100010010000000100011;
ROM[34459] <= 32'b00000000010000010000000100010011;
ROM[34460] <= 32'b00000000011000010010000000100011;
ROM[34461] <= 32'b00000000010000010000000100010011;
ROM[34462] <= 32'b00000001010000000000001110010011;
ROM[34463] <= 32'b00000000110000111000001110010011;
ROM[34464] <= 32'b01000000011100010000001110110011;
ROM[34465] <= 32'b00000000011100000000001000110011;
ROM[34466] <= 32'b00000000001000000000000110110011;
ROM[34467] <= 32'b00111000010000000010000011101111;
ROM[34468] <= 32'b11111111110000010000000100010011;
ROM[34469] <= 32'b00000000000000010010001110000011;
ROM[34470] <= 32'b00000000110100101000010000110011;
ROM[34471] <= 32'b00000000011101000010001000100011;
ROM[34472] <= 32'b00000000010100010010000000100011;
ROM[34473] <= 32'b00000000010000010000000100010011;
ROM[34474] <= 32'b00000000110100101000010000110011;
ROM[34475] <= 32'b00000000010001000010001110000011;
ROM[34476] <= 32'b00000000011100010010000000100011;
ROM[34477] <= 32'b00000000010000010000000100010011;
ROM[34478] <= 32'b00000000000000100010001110110111;
ROM[34479] <= 32'b10110000010000111000001110010011;
ROM[34480] <= 32'b00000000111000111000001110110011;
ROM[34481] <= 32'b00000000011100010010000000100011;
ROM[34482] <= 32'b00000000010000010000000100010011;
ROM[34483] <= 32'b00000000001100010010000000100011;
ROM[34484] <= 32'b00000000010000010000000100010011;
ROM[34485] <= 32'b00000000010000010010000000100011;
ROM[34486] <= 32'b00000000010000010000000100010011;
ROM[34487] <= 32'b00000000010100010010000000100011;
ROM[34488] <= 32'b00000000010000010000000100010011;
ROM[34489] <= 32'b00000000011000010010000000100011;
ROM[34490] <= 32'b00000000010000010000000100010011;
ROM[34491] <= 32'b00000001010000000000001110010011;
ROM[34492] <= 32'b00000000010000111000001110010011;
ROM[34493] <= 32'b01000000011100010000001110110011;
ROM[34494] <= 32'b00000000011100000000001000110011;
ROM[34495] <= 32'b00000000001000000000000110110011;
ROM[34496] <= 32'b01001001100000000100000011101111;
ROM[34497] <= 32'b00000000001000000000001110010011;
ROM[34498] <= 32'b00000000011100010010000000100011;
ROM[34499] <= 32'b00000000010000010000000100010011;
ROM[34500] <= 32'b00000000000000100010001110110111;
ROM[34501] <= 32'b10110101110000111000001110010011;
ROM[34502] <= 32'b00000000111000111000001110110011;
ROM[34503] <= 32'b00000000011100010010000000100011;
ROM[34504] <= 32'b00000000010000010000000100010011;
ROM[34505] <= 32'b00000000001100010010000000100011;
ROM[34506] <= 32'b00000000010000010000000100010011;
ROM[34507] <= 32'b00000000010000010010000000100011;
ROM[34508] <= 32'b00000000010000010000000100010011;
ROM[34509] <= 32'b00000000010100010010000000100011;
ROM[34510] <= 32'b00000000010000010000000100010011;
ROM[34511] <= 32'b00000000011000010010000000100011;
ROM[34512] <= 32'b00000000010000010000000100010011;
ROM[34513] <= 32'b00000001010000000000001110010011;
ROM[34514] <= 32'b00000000100000111000001110010011;
ROM[34515] <= 32'b01000000011100010000001110110011;
ROM[34516] <= 32'b00000000011100000000001000110011;
ROM[34517] <= 32'b00000000001000000000000110110011;
ROM[34518] <= 32'b10000101000011110000000011101111;
ROM[34519] <= 32'b00000000110100101000010000110011;
ROM[34520] <= 32'b00000000010001000010001110000011;
ROM[34521] <= 32'b00000000011100010010000000100011;
ROM[34522] <= 32'b00000000010000010000000100010011;
ROM[34523] <= 32'b00000000000000100010001110110111;
ROM[34524] <= 32'b10111011100000111000001110010011;
ROM[34525] <= 32'b00000000111000111000001110110011;
ROM[34526] <= 32'b00000000011100010010000000100011;
ROM[34527] <= 32'b00000000010000010000000100010011;
ROM[34528] <= 32'b00000000001100010010000000100011;
ROM[34529] <= 32'b00000000010000010000000100010011;
ROM[34530] <= 32'b00000000010000010010000000100011;
ROM[34531] <= 32'b00000000010000010000000100010011;
ROM[34532] <= 32'b00000000010100010010000000100011;
ROM[34533] <= 32'b00000000010000010000000100010011;
ROM[34534] <= 32'b00000000011000010010000000100011;
ROM[34535] <= 32'b00000000010000010000000100010011;
ROM[34536] <= 32'b00000001010000000000001110010011;
ROM[34537] <= 32'b00000000010000111000001110010011;
ROM[34538] <= 32'b01000000011100010000001110110011;
ROM[34539] <= 32'b00000000011100000000001000110011;
ROM[34540] <= 32'b00000000001000000000000110110011;
ROM[34541] <= 32'b01000100010000000100000011101111;
ROM[34542] <= 32'b00000000001000000000001110010011;
ROM[34543] <= 32'b00000000011100010010000000100011;
ROM[34544] <= 32'b00000000010000010000000100010011;
ROM[34545] <= 32'b00000000000000100010001110110111;
ROM[34546] <= 32'b11000001000000111000001110010011;
ROM[34547] <= 32'b00000000111000111000001110110011;
ROM[34548] <= 32'b00000000011100010010000000100011;
ROM[34549] <= 32'b00000000010000010000000100010011;
ROM[34550] <= 32'b00000000001100010010000000100011;
ROM[34551] <= 32'b00000000010000010000000100010011;
ROM[34552] <= 32'b00000000010000010010000000100011;
ROM[34553] <= 32'b00000000010000010000000100010011;
ROM[34554] <= 32'b00000000010100010010000000100011;
ROM[34555] <= 32'b00000000010000010000000100010011;
ROM[34556] <= 32'b00000000011000010010000000100011;
ROM[34557] <= 32'b00000000010000010000000100010011;
ROM[34558] <= 32'b00000001010000000000001110010011;
ROM[34559] <= 32'b00000000100000111000001110010011;
ROM[34560] <= 32'b01000000011100010000001110110011;
ROM[34561] <= 32'b00000000011100000000001000110011;
ROM[34562] <= 32'b00000000001000000000000110110011;
ROM[34563] <= 32'b11111001110111101111000011101111;
ROM[34564] <= 32'b00000000101000000000001110010011;
ROM[34565] <= 32'b00000000011100010010000000100011;
ROM[34566] <= 32'b00000000010000010000000100010011;
ROM[34567] <= 32'b00000000001100000000001110010011;
ROM[34568] <= 32'b00000000011100010010000000100011;
ROM[34569] <= 32'b00000000010000010000000100010011;
ROM[34570] <= 32'b00000000000000100010001110110111;
ROM[34571] <= 32'b11000111010000111000001110010011;
ROM[34572] <= 32'b00000000111000111000001110110011;
ROM[34573] <= 32'b00000000011100010010000000100011;
ROM[34574] <= 32'b00000000010000010000000100010011;
ROM[34575] <= 32'b00000000001100010010000000100011;
ROM[34576] <= 32'b00000000010000010000000100010011;
ROM[34577] <= 32'b00000000010000010010000000100011;
ROM[34578] <= 32'b00000000010000010000000100010011;
ROM[34579] <= 32'b00000000010100010010000000100011;
ROM[34580] <= 32'b00000000010000010000000100010011;
ROM[34581] <= 32'b00000000011000010010000000100011;
ROM[34582] <= 32'b00000000010000010000000100010011;
ROM[34583] <= 32'b00000001010000000000001110010011;
ROM[34584] <= 32'b00000001010000111000001110010011;
ROM[34585] <= 32'b01000000011100010000001110110011;
ROM[34586] <= 32'b00000000011100000000001000110011;
ROM[34587] <= 32'b00000000001000000000000110110011;
ROM[34588] <= 32'b11001000110111111101000011101111;
ROM[34589] <= 32'b11111111110000010000000100010011;
ROM[34590] <= 32'b00000000000000010010001110000011;
ROM[34591] <= 32'b00000000110100101000010000110011;
ROM[34592] <= 32'b00000000011101000010000000100011;
ROM[34593] <= 32'b00000000110100101000010000110011;
ROM[34594] <= 32'b00000000010001000010001110000011;
ROM[34595] <= 32'b00000000011100010010000000100011;
ROM[34596] <= 32'b00000000010000010000000100010011;
ROM[34597] <= 32'b00000000000000100010001110110111;
ROM[34598] <= 32'b11001110000000111000001110010011;
ROM[34599] <= 32'b00000000111000111000001110110011;
ROM[34600] <= 32'b00000000011100010010000000100011;
ROM[34601] <= 32'b00000000010000010000000100010011;
ROM[34602] <= 32'b00000000001100010010000000100011;
ROM[34603] <= 32'b00000000010000010000000100010011;
ROM[34604] <= 32'b00000000010000010010000000100011;
ROM[34605] <= 32'b00000000010000010000000100010011;
ROM[34606] <= 32'b00000000010100010010000000100011;
ROM[34607] <= 32'b00000000010000010000000100010011;
ROM[34608] <= 32'b00000000011000010010000000100011;
ROM[34609] <= 32'b00000000010000010000000100010011;
ROM[34610] <= 32'b00000001010000000000001110010011;
ROM[34611] <= 32'b00000000010000111000001110010011;
ROM[34612] <= 32'b01000000011100010000001110110011;
ROM[34613] <= 32'b00000000011100000000001000110011;
ROM[34614] <= 32'b00000000001000000000000110110011;
ROM[34615] <= 32'b01010110000000000011000011101111;
ROM[34616] <= 32'b11111111110000010000000100010011;
ROM[34617] <= 32'b00000000000000010010001110000011;
ROM[34618] <= 32'b00000000011101100010000000100011;
ROM[34619] <= 32'b00000000110100101000010000110011;
ROM[34620] <= 32'b00000000010001000010001110000011;
ROM[34621] <= 32'b00000000011100010010000000100011;
ROM[34622] <= 32'b00000000010000010000000100010011;
ROM[34623] <= 32'b00000000000000100010001110110111;
ROM[34624] <= 32'b11010100100000111000001110010011;
ROM[34625] <= 32'b00000000111000111000001110110011;
ROM[34626] <= 32'b00000000011100010010000000100011;
ROM[34627] <= 32'b00000000010000010000000100010011;
ROM[34628] <= 32'b00000000001100010010000000100011;
ROM[34629] <= 32'b00000000010000010000000100010011;
ROM[34630] <= 32'b00000000010000010010000000100011;
ROM[34631] <= 32'b00000000010000010000000100010011;
ROM[34632] <= 32'b00000000010100010010000000100011;
ROM[34633] <= 32'b00000000010000010000000100010011;
ROM[34634] <= 32'b00000000011000010010000000100011;
ROM[34635] <= 32'b00000000010000010000000100010011;
ROM[34636] <= 32'b00000001010000000000001110010011;
ROM[34637] <= 32'b00000000010000111000001110010011;
ROM[34638] <= 32'b01000000011100010000001110110011;
ROM[34639] <= 32'b00000000011100000000001000110011;
ROM[34640] <= 32'b00000000001000000000000110110011;
ROM[34641] <= 32'b00111010110000000101000011101111;
ROM[34642] <= 32'b11111111110000010000000100010011;
ROM[34643] <= 32'b00000000000000010010001110000011;
ROM[34644] <= 32'b00000000011101100010000000100011;
ROM[34645] <= 32'b00000000010100010010000000100011;
ROM[34646] <= 32'b00000000010000010000000100010011;
ROM[34647] <= 32'b00000001010000000000001110010011;
ROM[34648] <= 32'b01000000011100011000001110110011;
ROM[34649] <= 32'b00000000000000111010000010000011;
ROM[34650] <= 32'b11111111110000010000000100010011;
ROM[34651] <= 32'b00000000000000010010001110000011;
ROM[34652] <= 32'b00000000011100100010000000100011;
ROM[34653] <= 32'b00000000010000100000000100010011;
ROM[34654] <= 32'b00000001010000000000001110010011;
ROM[34655] <= 32'b01000000011100011000001110110011;
ROM[34656] <= 32'b00000000010000111010000110000011;
ROM[34657] <= 32'b00000000100000111010001000000011;
ROM[34658] <= 32'b00000000110000111010001010000011;
ROM[34659] <= 32'b00000001000000111010001100000011;
ROM[34660] <= 32'b00000000000000001000000011100111;
ROM[34661] <= 32'b00000000000000100010001110000011;
ROM[34662] <= 32'b00000000011100010010000000100011;
ROM[34663] <= 32'b00000000010000010000000100010011;
ROM[34664] <= 32'b11111111110000010000000100010011;
ROM[34665] <= 32'b00000000000000010010001110000011;
ROM[34666] <= 32'b00000000000000111000001010010011;
ROM[34667] <= 32'b00000000110100101000010000110011;
ROM[34668] <= 32'b00000000000001000010001110000011;
ROM[34669] <= 32'b00000000011100010010000000100011;
ROM[34670] <= 32'b00000000010000010000000100010011;
ROM[34671] <= 32'b00000000000000100010001110110111;
ROM[34672] <= 32'b11100000100000111000001110010011;
ROM[34673] <= 32'b00000000111000111000001110110011;
ROM[34674] <= 32'b00000000011100010010000000100011;
ROM[34675] <= 32'b00000000010000010000000100010011;
ROM[34676] <= 32'b00000000001100010010000000100011;
ROM[34677] <= 32'b00000000010000010000000100010011;
ROM[34678] <= 32'b00000000010000010010000000100011;
ROM[34679] <= 32'b00000000010000010000000100010011;
ROM[34680] <= 32'b00000000010100010010000000100011;
ROM[34681] <= 32'b00000000010000010000000100010011;
ROM[34682] <= 32'b00000000011000010010000000100011;
ROM[34683] <= 32'b00000000010000010000000100010011;
ROM[34684] <= 32'b00000001010000000000001110010011;
ROM[34685] <= 32'b00000000010000111000001110010011;
ROM[34686] <= 32'b01000000011100010000001110110011;
ROM[34687] <= 32'b00000000011100000000001000110011;
ROM[34688] <= 32'b00000000001000000000000110110011;
ROM[34689] <= 32'b11111101010111111101000011101111;
ROM[34690] <= 32'b11111111110000010000000100010011;
ROM[34691] <= 32'b00000000000000010010001110000011;
ROM[34692] <= 32'b00000000011101100010000000100011;
ROM[34693] <= 32'b00000000110100101000010000110011;
ROM[34694] <= 32'b00000000010001000010001110000011;
ROM[34695] <= 32'b00000000011100010010000000100011;
ROM[34696] <= 32'b00000000010000010000000100010011;
ROM[34697] <= 32'b00000000000000100010001110110111;
ROM[34698] <= 32'b11100111000000111000001110010011;
ROM[34699] <= 32'b00000000111000111000001110110011;
ROM[34700] <= 32'b00000000011100010010000000100011;
ROM[34701] <= 32'b00000000010000010000000100010011;
ROM[34702] <= 32'b00000000001100010010000000100011;
ROM[34703] <= 32'b00000000010000010000000100010011;
ROM[34704] <= 32'b00000000010000010010000000100011;
ROM[34705] <= 32'b00000000010000010000000100010011;
ROM[34706] <= 32'b00000000010100010010000000100011;
ROM[34707] <= 32'b00000000010000010000000100010011;
ROM[34708] <= 32'b00000000011000010010000000100011;
ROM[34709] <= 32'b00000000010000010000000100010011;
ROM[34710] <= 32'b00000001010000000000001110010011;
ROM[34711] <= 32'b00000000010000111000001110010011;
ROM[34712] <= 32'b01000000011100010000001110110011;
ROM[34713] <= 32'b00000000011100000000001000110011;
ROM[34714] <= 32'b00000000001000000000000110110011;
ROM[34715] <= 32'b00010010000000000011000011101111;
ROM[34716] <= 32'b11111111110000010000000100010011;
ROM[34717] <= 32'b00000000000000010010001110000011;
ROM[34718] <= 32'b00000000011101100010000000100011;
ROM[34719] <= 32'b00000000010100010010000000100011;
ROM[34720] <= 32'b00000000010000010000000100010011;
ROM[34721] <= 32'b00000000000000100010001110110111;
ROM[34722] <= 32'b11101101000000111000001110010011;
ROM[34723] <= 32'b00000000111000111000001110110011;
ROM[34724] <= 32'b00000000011100010010000000100011;
ROM[34725] <= 32'b00000000010000010000000100010011;
ROM[34726] <= 32'b00000000001100010010000000100011;
ROM[34727] <= 32'b00000000010000010000000100010011;
ROM[34728] <= 32'b00000000010000010010000000100011;
ROM[34729] <= 32'b00000000010000010000000100010011;
ROM[34730] <= 32'b00000000010100010010000000100011;
ROM[34731] <= 32'b00000000010000010000000100010011;
ROM[34732] <= 32'b00000000011000010010000000100011;
ROM[34733] <= 32'b00000000010000010000000100010011;
ROM[34734] <= 32'b00000001010000000000001110010011;
ROM[34735] <= 32'b00000000010000111000001110010011;
ROM[34736] <= 32'b01000000011100010000001110110011;
ROM[34737] <= 32'b00000000011100000000001000110011;
ROM[34738] <= 32'b00000000001000000000000110110011;
ROM[34739] <= 32'b11001001000111110001000011101111;
ROM[34740] <= 32'b11111111110000010000000100010011;
ROM[34741] <= 32'b00000000000000010010001110000011;
ROM[34742] <= 32'b00000000011101100010000000100011;
ROM[34743] <= 32'b00000000000000000000001110010011;
ROM[34744] <= 32'b00000000011100010010000000100011;
ROM[34745] <= 32'b00000000010000010000000100010011;
ROM[34746] <= 32'b00000001010000000000001110010011;
ROM[34747] <= 32'b01000000011100011000001110110011;
ROM[34748] <= 32'b00000000000000111010000010000011;
ROM[34749] <= 32'b11111111110000010000000100010011;
ROM[34750] <= 32'b00000000000000010010001110000011;
ROM[34751] <= 32'b00000000011100100010000000100011;
ROM[34752] <= 32'b00000000010000100000000100010011;
ROM[34753] <= 32'b00000001010000000000001110010011;
ROM[34754] <= 32'b01000000011100011000001110110011;
ROM[34755] <= 32'b00000000010000111010000110000011;
ROM[34756] <= 32'b00000000100000111010001000000011;
ROM[34757] <= 32'b00000000110000111010001010000011;
ROM[34758] <= 32'b00000001000000111010001100000011;
ROM[34759] <= 32'b00000000000000001000000011100111;
ROM[34760] <= 32'b00000000000000010010000000100011;
ROM[34761] <= 32'b00000000010000010000000100010011;
ROM[34762] <= 32'b00000000000000010010000000100011;
ROM[34763] <= 32'b00000000010000010000000100010011;
ROM[34764] <= 32'b00000000000000010010000000100011;
ROM[34765] <= 32'b00000000010000010000000100010011;
ROM[34766] <= 32'b00000000000000100010001110000011;
ROM[34767] <= 32'b00000000011100010010000000100011;
ROM[34768] <= 32'b00000000010000010000000100010011;
ROM[34769] <= 32'b11111111110000010000000100010011;
ROM[34770] <= 32'b00000000000000010010001110000011;
ROM[34771] <= 32'b00000000000000111000001010010011;
ROM[34772] <= 32'b00000000000000000000001110010011;
ROM[34773] <= 32'b00000000011100010010000000100011;
ROM[34774] <= 32'b00000000010000010000000100010011;
ROM[34775] <= 32'b11111111110000010000000100010011;
ROM[34776] <= 32'b00000000000000010010001110000011;
ROM[34777] <= 32'b00000000011100011010001000100011;
ROM[34778] <= 32'b00000000010000011010001110000011;
ROM[34779] <= 32'b00000000011100010010000000100011;
ROM[34780] <= 32'b00000000010000010000000100010011;
ROM[34781] <= 32'b11111111110000010000000100010011;
ROM[34782] <= 32'b00000000000000010010001110000011;
ROM[34783] <= 32'b01000000011100000000001110110011;
ROM[34784] <= 32'b00000000000100111000001110010011;
ROM[34785] <= 32'b00000000011100010010000000100011;
ROM[34786] <= 32'b00000000010000010000000100010011;
ROM[34787] <= 32'b11111111110000010000000100010011;
ROM[34788] <= 32'b00000000000000010010001110000011;
ROM[34789] <= 32'b01000000011100000000001110110011;
ROM[34790] <= 32'b00000000000100111000001110010011;
ROM[34791] <= 32'b00000000011100010010000000100011;
ROM[34792] <= 32'b00000000010000010000000100010011;
ROM[34793] <= 32'b11111111110000010000000100010011;
ROM[34794] <= 32'b00000000000000010010001110000011;
ROM[34795] <= 32'b00000000000000111000101001100011;
ROM[34796] <= 32'b00000000000000100011001110110111;
ROM[34797] <= 32'b01101101000000111000001110010011;
ROM[34798] <= 32'b00000000111000111000001110110011;
ROM[34799] <= 32'b00000000000000111000000011100111;
ROM[34800] <= 32'b00000000110100101000010000110011;
ROM[34801] <= 32'b00000000000001000010001110000011;
ROM[34802] <= 32'b00000000011100010010000000100011;
ROM[34803] <= 32'b00000000010000010000000100010011;
ROM[34804] <= 32'b00000000000000100010001110110111;
ROM[34805] <= 32'b00000001110000111000001110010011;
ROM[34806] <= 32'b00000000111000111000001110110011;
ROM[34807] <= 32'b00000000011100010010000000100011;
ROM[34808] <= 32'b00000000010000010000000100010011;
ROM[34809] <= 32'b00000000001100010010000000100011;
ROM[34810] <= 32'b00000000010000010000000100010011;
ROM[34811] <= 32'b00000000010000010010000000100011;
ROM[34812] <= 32'b00000000010000010000000100010011;
ROM[34813] <= 32'b00000000010100010010000000100011;
ROM[34814] <= 32'b00000000010000010000000100010011;
ROM[34815] <= 32'b00000000011000010010000000100011;
ROM[34816] <= 32'b00000000010000010000000100010011;
ROM[34817] <= 32'b00000001010000000000001110010011;
ROM[34818] <= 32'b00000000010000111000001110010011;
ROM[34819] <= 32'b01000000011100010000001110110011;
ROM[34820] <= 32'b00000000011100000000001000110011;
ROM[34821] <= 32'b00000000001000000000000110110011;
ROM[34822] <= 32'b10000011110111111110000011101111;
ROM[34823] <= 32'b11111111110000010000000100010011;
ROM[34824] <= 32'b00000000000000010010001110000011;
ROM[34825] <= 32'b00000000011101100010000000100011;
ROM[34826] <= 32'b00000000110100101000010000110011;
ROM[34827] <= 32'b00000001000001000010001110000011;
ROM[34828] <= 32'b00000000011100010010000000100011;
ROM[34829] <= 32'b00000000010000010000000100010011;
ROM[34830] <= 32'b11111111110000010000000100010011;
ROM[34831] <= 32'b00000000000000010010001110000011;
ROM[34832] <= 32'b00000000000000111000101001100011;
ROM[34833] <= 32'b00000000000000100010001110110111;
ROM[34834] <= 32'b00000101100000111000001110010011;
ROM[34835] <= 32'b00000000111000111000001110110011;
ROM[34836] <= 32'b00000000000000111000000011100111;
ROM[34837] <= 32'b00110111110000000000000011101111;
ROM[34838] <= 32'b00000000000000000000001110010011;
ROM[34839] <= 32'b00000000011100010010000000100011;
ROM[34840] <= 32'b00000000010000010000000100010011;
ROM[34841] <= 32'b11111111110000010000000100010011;
ROM[34842] <= 32'b00000000000000010010001110000011;
ROM[34843] <= 32'b00000000011100011010000000100011;
ROM[34844] <= 32'b00000000000000011010001110000011;
ROM[34845] <= 32'b00000000011100010010000000100011;
ROM[34846] <= 32'b00000000010000010000000100010011;
ROM[34847] <= 32'b11111111110000010000000100010011;
ROM[34848] <= 32'b00000000000000010010001110000011;
ROM[34849] <= 32'b01000000011100000000001110110011;
ROM[34850] <= 32'b00000000000100111000001110010011;
ROM[34851] <= 32'b00000000011100010010000000100011;
ROM[34852] <= 32'b00000000010000010000000100010011;
ROM[34853] <= 32'b11111111110000010000000100010011;
ROM[34854] <= 32'b00000000000000010010001110000011;
ROM[34855] <= 32'b01000000011100000000001110110011;
ROM[34856] <= 32'b00000000000100111000001110010011;
ROM[34857] <= 32'b00000000011100010010000000100011;
ROM[34858] <= 32'b00000000010000010000000100010011;
ROM[34859] <= 32'b11111111110000010000000100010011;
ROM[34860] <= 32'b00000000000000010010001110000011;
ROM[34861] <= 32'b00000000000000111000101001100011;
ROM[34862] <= 32'b00000000000000100010001110110111;
ROM[34863] <= 32'b00111101000000111000001110010011;
ROM[34864] <= 32'b00000000111000111000001110110011;
ROM[34865] <= 32'b00000000000000111000000011100111;
ROM[34866] <= 32'b00000000000000000000001110010011;
ROM[34867] <= 32'b00000000011100010010000000100011;
ROM[34868] <= 32'b00000000010000010000000100010011;
ROM[34869] <= 32'b11111111110000010000000100010011;
ROM[34870] <= 32'b00000000000000010010001110000011;
ROM[34871] <= 32'b00000000011100011010010000100011;
ROM[34872] <= 32'b00000000100000011010001110000011;
ROM[34873] <= 32'b00000000011100010010000000100011;
ROM[34874] <= 32'b00000000010000010000000100010011;
ROM[34875] <= 32'b11111111110000010000000100010011;
ROM[34876] <= 32'b00000000000000010010001110000011;
ROM[34877] <= 32'b01000000011100000000001110110011;
ROM[34878] <= 32'b00000000000100111000001110010011;
ROM[34879] <= 32'b00000000011100010010000000100011;
ROM[34880] <= 32'b00000000010000010000000100010011;
ROM[34881] <= 32'b11111111110000010000000100010011;
ROM[34882] <= 32'b00000000000000010010001110000011;
ROM[34883] <= 32'b01000000011100000000001110110011;
ROM[34884] <= 32'b00000000000100111000001110010011;
ROM[34885] <= 32'b00000000011100010010000000100011;
ROM[34886] <= 32'b00000000010000010000000100010011;
ROM[34887] <= 32'b11111111110000010000000100010011;
ROM[34888] <= 32'b00000000000000010010001110000011;
ROM[34889] <= 32'b00000000000000111000101001100011;
ROM[34890] <= 32'b00000000000000100010001110110111;
ROM[34891] <= 32'b00011001010000111000001110010011;
ROM[34892] <= 32'b00000000111000111000001110110011;
ROM[34893] <= 32'b00000000000000111000000011100111;
ROM[34894] <= 32'b00000000000000100010001110110111;
ROM[34895] <= 32'b00011000010000111000001110010011;
ROM[34896] <= 32'b00000000111000111000001110110011;
ROM[34897] <= 32'b00000000011100010010000000100011;
ROM[34898] <= 32'b00000000010000010000000100010011;
ROM[34899] <= 32'b00000000001100010010000000100011;
ROM[34900] <= 32'b00000000010000010000000100010011;
ROM[34901] <= 32'b00000000010000010010000000100011;
ROM[34902] <= 32'b00000000010000010000000100010011;
ROM[34903] <= 32'b00000000010100010010000000100011;
ROM[34904] <= 32'b00000000010000010000000100010011;
ROM[34905] <= 32'b00000000011000010010000000100011;
ROM[34906] <= 32'b00000000010000010000000100010011;
ROM[34907] <= 32'b00000001010000000000001110010011;
ROM[34908] <= 32'b00000000000000111000001110010011;
ROM[34909] <= 32'b01000000011100010000001110110011;
ROM[34910] <= 32'b00000000011100000000001000110011;
ROM[34911] <= 32'b00000000001000000000000110110011;
ROM[34912] <= 32'b11101101100011101011000011101111;
ROM[34913] <= 32'b11111111110000010000000100010011;
ROM[34914] <= 32'b00000000000000010010001110000011;
ROM[34915] <= 32'b00000000011100011010010000100011;
ROM[34916] <= 32'b11110101000111111111000011101111;
ROM[34917] <= 32'b00000000100000011010001110000011;
ROM[34918] <= 32'b00000000011100010010000000100011;
ROM[34919] <= 32'b00000000010000010000000100010011;
ROM[34920] <= 32'b00000101000000000000001110010011;
ROM[34921] <= 32'b00000000011100010010000000100011;
ROM[34922] <= 32'b00000000010000010000000100010011;
ROM[34923] <= 32'b11111111110000010000000100010011;
ROM[34924] <= 32'b00000000000000010010001110000011;
ROM[34925] <= 32'b11111111110000010000000100010011;
ROM[34926] <= 32'b00000000000000010010010000000011;
ROM[34927] <= 32'b00000000011101000010010010110011;
ROM[34928] <= 32'b00000000100000111010010100110011;
ROM[34929] <= 32'b00000000101001001000001110110011;
ROM[34930] <= 32'b00000000000100111000001110010011;
ROM[34931] <= 32'b00000000000100111111001110010011;
ROM[34932] <= 32'b00000000011100010010000000100011;
ROM[34933] <= 32'b00000000010000010000000100010011;
ROM[34934] <= 32'b11111111110000010000000100010011;
ROM[34935] <= 32'b00000000000000010010001110000011;
ROM[34936] <= 32'b00000000000000111000101001100011;
ROM[34937] <= 32'b00000000000000100010001110110111;
ROM[34938] <= 32'b00011111100000111000001110010011;
ROM[34939] <= 32'b00000000111000111000001110110011;
ROM[34940] <= 32'b00000000000000111000000011100111;
ROM[34941] <= 32'b00000100110000000000000011101111;
ROM[34942] <= 32'b00000000000100000000001110010011;
ROM[34943] <= 32'b00000000011100010010000000100011;
ROM[34944] <= 32'b00000000010000010000000100010011;
ROM[34945] <= 32'b11111111110000010000000100010011;
ROM[34946] <= 32'b00000000000000010010001110000011;
ROM[34947] <= 32'b01000000011100000000001110110011;
ROM[34948] <= 32'b00000000011100010010000000100011;
ROM[34949] <= 32'b00000000010000010000000100010011;
ROM[34950] <= 32'b11111111110000010000000100010011;
ROM[34951] <= 32'b00000000000000010010001110000011;
ROM[34952] <= 32'b00000000011100011010000000100011;
ROM[34953] <= 32'b00000000000000000000001110010011;
ROM[34954] <= 32'b00000000011100010010000000100011;
ROM[34955] <= 32'b00000000010000010000000100010011;
ROM[34956] <= 32'b11111111110000010000000100010011;
ROM[34957] <= 32'b00000000000000010010001110000011;
ROM[34958] <= 32'b00000000110100101000010000110011;
ROM[34959] <= 32'b00000000011101000010100000100011;
ROM[34960] <= 32'b00000000100000011010001110000011;
ROM[34961] <= 32'b00000000011100010010000000100011;
ROM[34962] <= 32'b00000000010000010000000100010011;
ROM[34963] <= 32'b00000101000100000000001110010011;
ROM[34964] <= 32'b00000000011100010010000000100011;
ROM[34965] <= 32'b00000000010000010000000100010011;
ROM[34966] <= 32'b11111111110000010000000100010011;
ROM[34967] <= 32'b00000000000000010010001110000011;
ROM[34968] <= 32'b11111111110000010000000100010011;
ROM[34969] <= 32'b00000000000000010010010000000011;
ROM[34970] <= 32'b00000000011101000010010010110011;
ROM[34971] <= 32'b00000000100000111010010100110011;
ROM[34972] <= 32'b00000000101001001000001110110011;
ROM[34973] <= 32'b00000000000100111000001110010011;
ROM[34974] <= 32'b00000000000100111111001110010011;
ROM[34975] <= 32'b00000000011100010010000000100011;
ROM[34976] <= 32'b00000000010000010000000100010011;
ROM[34977] <= 32'b11111111110000010000000100010011;
ROM[34978] <= 32'b00000000000000010010001110000011;
ROM[34979] <= 32'b00000000000000111000101001100011;
ROM[34980] <= 32'b00000000000000100010001110110111;
ROM[34981] <= 32'b00101010010000111000001110010011;
ROM[34982] <= 32'b00000000111000111000001110110011;
ROM[34983] <= 32'b00000000000000111000000011100111;
ROM[34984] <= 32'b00000101110000000000000011101111;
ROM[34985] <= 32'b00000000000100000000001110010011;
ROM[34986] <= 32'b00000000011100010010000000100011;
ROM[34987] <= 32'b00000000010000010000000100010011;
ROM[34988] <= 32'b11111111110000010000000100010011;
ROM[34989] <= 32'b00000000000000010010001110000011;
ROM[34990] <= 32'b01000000011100000000001110110011;
ROM[34991] <= 32'b00000000011100010010000000100011;
ROM[34992] <= 32'b00000000010000010000000100010011;
ROM[34993] <= 32'b11111111110000010000000100010011;
ROM[34994] <= 32'b00000000000000010010001110000011;
ROM[34995] <= 32'b00000000011100011010000000100011;
ROM[34996] <= 32'b00000000000100000000001110010011;
ROM[34997] <= 32'b00000000011100010010000000100011;
ROM[34998] <= 32'b00000000010000010000000100010011;
ROM[34999] <= 32'b11111111110000010000000100010011;
ROM[35000] <= 32'b00000000000000010010001110000011;
ROM[35001] <= 32'b01000000011100000000001110110011;
ROM[35002] <= 32'b00000000011100010010000000100011;
ROM[35003] <= 32'b00000000010000010000000100010011;
ROM[35004] <= 32'b11111111110000010000000100010011;
ROM[35005] <= 32'b00000000000000010010001110000011;
ROM[35006] <= 32'b00000000011100011010001000100011;
ROM[35007] <= 32'b00000000110100101000010000110011;
ROM[35008] <= 32'b00000000010001000010001110000011;
ROM[35009] <= 32'b00000000011100010010000000100011;
ROM[35010] <= 32'b00000000010000010000000100010011;
ROM[35011] <= 32'b00000000000000100010001110110111;
ROM[35012] <= 32'b00110101100000111000001110010011;
ROM[35013] <= 32'b00000000111000111000001110110011;
ROM[35014] <= 32'b00000000011100010010000000100011;
ROM[35015] <= 32'b00000000010000010000000100010011;
ROM[35016] <= 32'b00000000001100010010000000100011;
ROM[35017] <= 32'b00000000010000010000000100010011;
ROM[35018] <= 32'b00000000010000010010000000100011;
ROM[35019] <= 32'b00000000010000010000000100010011;
ROM[35020] <= 32'b00000000010100010010000000100011;
ROM[35021] <= 32'b00000000010000010000000100010011;
ROM[35022] <= 32'b00000000011000010010000000100011;
ROM[35023] <= 32'b00000000010000010000000100010011;
ROM[35024] <= 32'b00000001010000000000001110010011;
ROM[35025] <= 32'b00000000010000111000001110010011;
ROM[35026] <= 32'b01000000011100010000001110110011;
ROM[35027] <= 32'b00000000011100000000001000110011;
ROM[35028] <= 32'b00000000001000000000000110110011;
ROM[35029] <= 32'b01011001110100000100000011101111;
ROM[35030] <= 32'b11111111110000010000000100010011;
ROM[35031] <= 32'b00000000000000010010001110000011;
ROM[35032] <= 32'b00000000011101100010000000100011;
ROM[35033] <= 32'b00000000110100101000010000110011;
ROM[35034] <= 32'b00000001100001000010001110000011;
ROM[35035] <= 32'b00000000011100010010000000100011;
ROM[35036] <= 32'b00000000010000010000000100010011;
ROM[35037] <= 32'b00000000000000100010001110110111;
ROM[35038] <= 32'b00111100000000111000001110010011;
ROM[35039] <= 32'b00000000111000111000001110110011;
ROM[35040] <= 32'b00000000011100010010000000100011;
ROM[35041] <= 32'b00000000010000010000000100010011;
ROM[35042] <= 32'b00000000001100010010000000100011;
ROM[35043] <= 32'b00000000010000010000000100010011;
ROM[35044] <= 32'b00000000010000010010000000100011;
ROM[35045] <= 32'b00000000010000010000000100010011;
ROM[35046] <= 32'b00000000010100010010000000100011;
ROM[35047] <= 32'b00000000010000010000000100010011;
ROM[35048] <= 32'b00000000011000010010000000100011;
ROM[35049] <= 32'b00000000010000010000000100010011;
ROM[35050] <= 32'b00000001010000000000001110010011;
ROM[35051] <= 32'b00000000010000111000001110010011;
ROM[35052] <= 32'b01000000011100010000001110110011;
ROM[35053] <= 32'b00000000011100000000001000110011;
ROM[35054] <= 32'b00000000001000000000000110110011;
ROM[35055] <= 32'b01010000100100001000000011101111;
ROM[35056] <= 32'b11111111110000010000000100010011;
ROM[35057] <= 32'b00000000000000010010001110000011;
ROM[35058] <= 32'b00000000011101100010000000100011;
ROM[35059] <= 32'b11001010010111111111000011101111;
ROM[35060] <= 32'b00000000000000100010001110110111;
ROM[35061] <= 32'b01000001110000111000001110010011;
ROM[35062] <= 32'b00000000111000111000001110110011;
ROM[35063] <= 32'b00000000011100010010000000100011;
ROM[35064] <= 32'b00000000010000010000000100010011;
ROM[35065] <= 32'b00000000001100010010000000100011;
ROM[35066] <= 32'b00000000010000010000000100010011;
ROM[35067] <= 32'b00000000010000010010000000100011;
ROM[35068] <= 32'b00000000010000010000000100010011;
ROM[35069] <= 32'b00000000010100010010000000100011;
ROM[35070] <= 32'b00000000010000010000000100010011;
ROM[35071] <= 32'b00000000011000010010000000100011;
ROM[35072] <= 32'b00000000010000010000000100010011;
ROM[35073] <= 32'b00000001010000000000001110010011;
ROM[35074] <= 32'b00000000000000111000001110010011;
ROM[35075] <= 32'b01000000011100010000001110110011;
ROM[35076] <= 32'b00000000011100000000001000110011;
ROM[35077] <= 32'b00000000001000000000000110110011;
ROM[35078] <= 32'b11000100000011101011000011101111;
ROM[35079] <= 32'b11111111110000010000000100010011;
ROM[35080] <= 32'b00000000000000010010001110000011;
ROM[35081] <= 32'b00000000011100011010010000100011;
ROM[35082] <= 32'b00000000100000011010001110000011;
ROM[35083] <= 32'b00000000011100010010000000100011;
ROM[35084] <= 32'b00000000010000010000000100010011;
ROM[35085] <= 32'b00000101000000000000001110010011;
ROM[35086] <= 32'b00000000011100010010000000100011;
ROM[35087] <= 32'b00000000010000010000000100010011;
ROM[35088] <= 32'b11111111110000010000000100010011;
ROM[35089] <= 32'b00000000000000010010001110000011;
ROM[35090] <= 32'b11111111110000010000000100010011;
ROM[35091] <= 32'b00000000000000010010010000000011;
ROM[35092] <= 32'b00000000011101000010010010110011;
ROM[35093] <= 32'b00000000100000111010010100110011;
ROM[35094] <= 32'b00000000101001001000001110110011;
ROM[35095] <= 32'b00000000000100111000001110010011;
ROM[35096] <= 32'b00000000000100111111001110010011;
ROM[35097] <= 32'b00000000011100010010000000100011;
ROM[35098] <= 32'b00000000010000010000000100010011;
ROM[35099] <= 32'b11111111110000010000000100010011;
ROM[35100] <= 32'b00000000000000010010001110000011;
ROM[35101] <= 32'b00000000000000111000101001100011;
ROM[35102] <= 32'b00000000000000100010001110110111;
ROM[35103] <= 32'b01001000110000111000001110010011;
ROM[35104] <= 32'b00000000111000111000001110110011;
ROM[35105] <= 32'b00000000000000111000000011100111;
ROM[35106] <= 32'b00000011010000000000000011101111;
ROM[35107] <= 32'b00000000000100000000001110010011;
ROM[35108] <= 32'b00000000011100010010000000100011;
ROM[35109] <= 32'b00000000010000010000000100010011;
ROM[35110] <= 32'b11111111110000010000000100010011;
ROM[35111] <= 32'b00000000000000010010001110000011;
ROM[35112] <= 32'b01000000011100000000001110110011;
ROM[35113] <= 32'b00000000011100010010000000100011;
ROM[35114] <= 32'b00000000010000010000000100010011;
ROM[35115] <= 32'b11111111110000010000000100010011;
ROM[35116] <= 32'b00000000000000010010001110000011;
ROM[35117] <= 32'b00000000110100101000010000110011;
ROM[35118] <= 32'b00000000011101000010100000100011;
ROM[35119] <= 32'b00000000100000011010001110000011;
ROM[35120] <= 32'b00000000011100010010000000100011;
ROM[35121] <= 32'b00000000010000010000000100010011;
ROM[35122] <= 32'b00000101000100000000001110010011;
ROM[35123] <= 32'b00000000011100010010000000100011;
ROM[35124] <= 32'b00000000010000010000000100010011;
ROM[35125] <= 32'b11111111110000010000000100010011;
ROM[35126] <= 32'b00000000000000010010001110000011;
ROM[35127] <= 32'b11111111110000010000000100010011;
ROM[35128] <= 32'b00000000000000010010010000000011;
ROM[35129] <= 32'b00000000011101000010010010110011;
ROM[35130] <= 32'b00000000100000111010010100110011;
ROM[35131] <= 32'b00000000101001001000001110110011;
ROM[35132] <= 32'b00000000000100111000001110010011;
ROM[35133] <= 32'b00000000000100111111001110010011;
ROM[35134] <= 32'b00000000011100010010000000100011;
ROM[35135] <= 32'b00000000010000010000000100010011;
ROM[35136] <= 32'b11111111110000010000000100010011;
ROM[35137] <= 32'b00000000000000010010001110000011;
ROM[35138] <= 32'b00000000000000111000101001100011;
ROM[35139] <= 32'b00000000000000100010001110110111;
ROM[35140] <= 32'b01010010000000111000001110010011;
ROM[35141] <= 32'b00000000111000111000001110110011;
ROM[35142] <= 32'b00000000000000111000000011100111;
ROM[35143] <= 32'b00000011000000000000000011101111;
ROM[35144] <= 32'b00000000000100000000001110010011;
ROM[35145] <= 32'b00000000011100010010000000100011;
ROM[35146] <= 32'b00000000010000010000000100010011;
ROM[35147] <= 32'b11111111110000010000000100010011;
ROM[35148] <= 32'b00000000000000010010001110000011;
ROM[35149] <= 32'b01000000011100000000001110110011;
ROM[35150] <= 32'b00000000011100010010000000100011;
ROM[35151] <= 32'b00000000010000010000000100010011;
ROM[35152] <= 32'b11111111110000010000000100010011;
ROM[35153] <= 32'b00000000000000010010001110000011;
ROM[35154] <= 32'b00000000011100011010001000100011;
ROM[35155] <= 32'b00000000100000011010001110000011;
ROM[35156] <= 32'b00000000011100010010000000100011;
ROM[35157] <= 32'b00000000010000010000000100010011;
ROM[35158] <= 32'b00001000001000000000001110010011;
ROM[35159] <= 32'b00000000011100010010000000100011;
ROM[35160] <= 32'b00000000010000010000000100010011;
ROM[35161] <= 32'b11111111110000010000000100010011;
ROM[35162] <= 32'b00000000000000010010001110000011;
ROM[35163] <= 32'b11111111110000010000000100010011;
ROM[35164] <= 32'b00000000000000010010010000000011;
ROM[35165] <= 32'b00000000011101000010010010110011;
ROM[35166] <= 32'b00000000100000111010010100110011;
ROM[35167] <= 32'b00000000101001001000001110110011;
ROM[35168] <= 32'b00000000000100111000001110010011;
ROM[35169] <= 32'b00000000000100111111001110010011;
ROM[35170] <= 32'b00000000011100010010000000100011;
ROM[35171] <= 32'b00000000010000010000000100010011;
ROM[35172] <= 32'b11111111110000010000000100010011;
ROM[35173] <= 32'b00000000000000010010001110000011;
ROM[35174] <= 32'b00000000000000111000101001100011;
ROM[35175] <= 32'b00000000000000100010001110110111;
ROM[35176] <= 32'b01011011000000111000001110010011;
ROM[35177] <= 32'b00000000111000111000001110110011;
ROM[35178] <= 32'b00000000000000111000000011100111;
ROM[35179] <= 32'b00100101010000000000000011101111;
ROM[35180] <= 32'b00000000110100101000010000110011;
ROM[35181] <= 32'b00000000000001000010001110000011;
ROM[35182] <= 32'b00000000011100010010000000100011;
ROM[35183] <= 32'b00000000010000010000000100010011;
ROM[35184] <= 32'b00000000000000100010001110110111;
ROM[35185] <= 32'b01100000110000111000001110010011;
ROM[35186] <= 32'b00000000111000111000001110110011;
ROM[35187] <= 32'b00000000011100010010000000100011;
ROM[35188] <= 32'b00000000010000010000000100010011;
ROM[35189] <= 32'b00000000001100010010000000100011;
ROM[35190] <= 32'b00000000010000010000000100010011;
ROM[35191] <= 32'b00000000010000010010000000100011;
ROM[35192] <= 32'b00000000010000010000000100010011;
ROM[35193] <= 32'b00000000010100010010000000100011;
ROM[35194] <= 32'b00000000010000010000000100010011;
ROM[35195] <= 32'b00000000011000010010000000100011;
ROM[35196] <= 32'b00000000010000010000000100010011;
ROM[35197] <= 32'b00000001010000000000001110010011;
ROM[35198] <= 32'b00000000010000111000001110010011;
ROM[35199] <= 32'b01000000011100010000001110110011;
ROM[35200] <= 32'b00000000011100000000001000110011;
ROM[35201] <= 32'b00000000001000000000000110110011;
ROM[35202] <= 32'b10010111010011111110000011101111;
ROM[35203] <= 32'b00000000000100000000001110010011;
ROM[35204] <= 32'b00000000011100010010000000100011;
ROM[35205] <= 32'b00000000010000010000000100010011;
ROM[35206] <= 32'b11111111110000010000000100010011;
ROM[35207] <= 32'b00000000000000010010001110000011;
ROM[35208] <= 32'b11111111110000010000000100010011;
ROM[35209] <= 32'b00000000000000010010010000000011;
ROM[35210] <= 32'b00000000011101000010010010110011;
ROM[35211] <= 32'b00000000100000111010010100110011;
ROM[35212] <= 32'b00000000101001001000001110110011;
ROM[35213] <= 32'b00000000000100111000001110010011;
ROM[35214] <= 32'b00000000000100111111001110010011;
ROM[35215] <= 32'b00000000011100010010000000100011;
ROM[35216] <= 32'b00000000010000010000000100010011;
ROM[35217] <= 32'b11111111110000010000000100010011;
ROM[35218] <= 32'b00000000000000010010001110000011;
ROM[35219] <= 32'b00000000000000111000101001100011;
ROM[35220] <= 32'b00000000000000100010001110110111;
ROM[35221] <= 32'b01100110010000111000001110010011;
ROM[35222] <= 32'b00000000111000111000001110110011;
ROM[35223] <= 32'b00000000000000111000000011100111;
ROM[35224] <= 32'b00000111100000000000000011101111;
ROM[35225] <= 32'b00000000110100101000010000110011;
ROM[35226] <= 32'b00000000000001000010001110000011;
ROM[35227] <= 32'b00000000011100010010000000100011;
ROM[35228] <= 32'b00000000010000010000000100010011;
ROM[35229] <= 32'b00000000001100000000001110010011;
ROM[35230] <= 32'b00000000011100010010000000100011;
ROM[35231] <= 32'b00000000010000010000000100010011;
ROM[35232] <= 32'b00000000000000100010001110110111;
ROM[35233] <= 32'b01101100110000111000001110010011;
ROM[35234] <= 32'b00000000111000111000001110110011;
ROM[35235] <= 32'b00000000011100010010000000100011;
ROM[35236] <= 32'b00000000010000010000000100010011;
ROM[35237] <= 32'b00000000001100010010000000100011;
ROM[35238] <= 32'b00000000010000010000000100010011;
ROM[35239] <= 32'b00000000010000010010000000100011;
ROM[35240] <= 32'b00000000010000010000000100010011;
ROM[35241] <= 32'b00000000010100010010000000100011;
ROM[35242] <= 32'b00000000010000010000000100010011;
ROM[35243] <= 32'b00000000011000010010000000100011;
ROM[35244] <= 32'b00000000010000010000000100010011;
ROM[35245] <= 32'b00000001010000000000001110010011;
ROM[35246] <= 32'b00000000100000111000001110010011;
ROM[35247] <= 32'b01000000011100010000001110110011;
ROM[35248] <= 32'b00000000011100000000001000110011;
ROM[35249] <= 32'b00000000001000000000000110110011;
ROM[35250] <= 32'b10010001010011111110000011101111;
ROM[35251] <= 32'b11111111110000010000000100010011;
ROM[35252] <= 32'b00000000000000010010001110000011;
ROM[35253] <= 32'b00000000011101100010000000100011;
ROM[35254] <= 32'b00000000110100101000010000110011;
ROM[35255] <= 32'b00000000000001000010001110000011;
ROM[35256] <= 32'b00000000011100010010000000100011;
ROM[35257] <= 32'b00000000010000010000000100010011;
ROM[35258] <= 32'b00000000000000100010001110110111;
ROM[35259] <= 32'b01110011010000111000001110010011;
ROM[35260] <= 32'b00000000111000111000001110110011;
ROM[35261] <= 32'b00000000011100010010000000100011;
ROM[35262] <= 32'b00000000010000010000000100010011;
ROM[35263] <= 32'b00000000001100010010000000100011;
ROM[35264] <= 32'b00000000010000010000000100010011;
ROM[35265] <= 32'b00000000010000010010000000100011;
ROM[35266] <= 32'b00000000010000010000000100010011;
ROM[35267] <= 32'b00000000010100010010000000100011;
ROM[35268] <= 32'b00000000010000010000000100010011;
ROM[35269] <= 32'b00000000011000010010000000100011;
ROM[35270] <= 32'b00000000010000010000000100010011;
ROM[35271] <= 32'b00000001010000000000001110010011;
ROM[35272] <= 32'b00000000010000111000001110010011;
ROM[35273] <= 32'b01000000011100010000001110110011;
ROM[35274] <= 32'b00000000011100000000001000110011;
ROM[35275] <= 32'b00000000001000000000000110110011;
ROM[35276] <= 32'b10000100110011111110000011101111;
ROM[35277] <= 32'b00000000001000000000001110010011;
ROM[35278] <= 32'b00000000011100010010000000100011;
ROM[35279] <= 32'b00000000010000010000000100010011;
ROM[35280] <= 32'b11111111110000010000000100010011;
ROM[35281] <= 32'b00000000000000010010001110000011;
ROM[35282] <= 32'b11111111110000010000000100010011;
ROM[35283] <= 32'b00000000000000010010010000000011;
ROM[35284] <= 32'b00000000011101000010010010110011;
ROM[35285] <= 32'b00000000100000111010010100110011;
ROM[35286] <= 32'b00000000101001001000001110110011;
ROM[35287] <= 32'b00000000000100111000001110010011;
ROM[35288] <= 32'b00000000000100111111001110010011;
ROM[35289] <= 32'b00000000011100010010000000100011;
ROM[35290] <= 32'b00000000010000010000000100010011;
ROM[35291] <= 32'b11111111110000010000000100010011;
ROM[35292] <= 32'b00000000000000010010001110000011;
ROM[35293] <= 32'b00000000000000111000101001100011;
ROM[35294] <= 32'b00000000000000100010001110110111;
ROM[35295] <= 32'b01111000110000111000001110010011;
ROM[35296] <= 32'b00000000111000111000001110110011;
ROM[35297] <= 32'b00000000000000111000000011100111;
ROM[35298] <= 32'b00000111100000000000000011101111;
ROM[35299] <= 32'b00000000110100101000010000110011;
ROM[35300] <= 32'b00000000000001000010001110000011;
ROM[35301] <= 32'b00000000011100010010000000100011;
ROM[35302] <= 32'b00000000010000010000000100010011;
ROM[35303] <= 32'b00000000001100000000001110010011;
ROM[35304] <= 32'b00000000011100010010000000100011;
ROM[35305] <= 32'b00000000010000010000000100010011;
ROM[35306] <= 32'b00000000000000100010001110110111;
ROM[35307] <= 32'b01111111010000111000001110010011;
ROM[35308] <= 32'b00000000111000111000001110110011;
ROM[35309] <= 32'b00000000011100010010000000100011;
ROM[35310] <= 32'b00000000010000010000000100010011;
ROM[35311] <= 32'b00000000001100010010000000100011;
ROM[35312] <= 32'b00000000010000010000000100010011;
ROM[35313] <= 32'b00000000010000010010000000100011;
ROM[35314] <= 32'b00000000010000010000000100010011;
ROM[35315] <= 32'b00000000010100010010000000100011;
ROM[35316] <= 32'b00000000010000010000000100010011;
ROM[35317] <= 32'b00000000011000010010000000100011;
ROM[35318] <= 32'b00000000010000010000000100010011;
ROM[35319] <= 32'b00000001010000000000001110010011;
ROM[35320] <= 32'b00000000100000111000001110010011;
ROM[35321] <= 32'b01000000011100010000001110110011;
ROM[35322] <= 32'b00000000011100000000001000110011;
ROM[35323] <= 32'b00000000001000000000000110110011;
ROM[35324] <= 32'b11111110110111111101000011101111;
ROM[35325] <= 32'b11111111110000010000000100010011;
ROM[35326] <= 32'b00000000000000010010001110000011;
ROM[35327] <= 32'b00000000011101100010000000100011;
ROM[35328] <= 32'b00000000100000011010001110000011;
ROM[35329] <= 32'b00000000011100010010000000100011;
ROM[35330] <= 32'b00000000010000010000000100010011;
ROM[35331] <= 32'b00001000001100000000001110010011;
ROM[35332] <= 32'b00000000011100010010000000100011;
ROM[35333] <= 32'b00000000010000010000000100010011;
ROM[35334] <= 32'b11111111110000010000000100010011;
ROM[35335] <= 32'b00000000000000010010001110000011;
ROM[35336] <= 32'b11111111110000010000000100010011;
ROM[35337] <= 32'b00000000000000010010010000000011;
ROM[35338] <= 32'b00000000011101000010010010110011;
ROM[35339] <= 32'b00000000100000111010010100110011;
ROM[35340] <= 32'b00000000101001001000001110110011;
ROM[35341] <= 32'b00000000000100111000001110010011;
ROM[35342] <= 32'b00000000000100111111001110010011;
ROM[35343] <= 32'b00000000011100010010000000100011;
ROM[35344] <= 32'b00000000010000010000000100010011;
ROM[35345] <= 32'b11111111110000010000000100010011;
ROM[35346] <= 32'b00000000000000010010001110000011;
ROM[35347] <= 32'b00000000000000111000101001100011;
ROM[35348] <= 32'b00000000000000100011001110110111;
ROM[35349] <= 32'b10000110010000111000001110010011;
ROM[35350] <= 32'b00000000111000111000001110110011;
ROM[35351] <= 32'b00000000000000111000000011100111;
ROM[35352] <= 32'b00100101010000000000000011101111;
ROM[35353] <= 32'b00000000110100101000010000110011;
ROM[35354] <= 32'b00000000000001000010001110000011;
ROM[35355] <= 32'b00000000011100010010000000100011;
ROM[35356] <= 32'b00000000010000010000000100010011;
ROM[35357] <= 32'b00000000000000100011001110110111;
ROM[35358] <= 32'b10001100000000111000001110010011;
ROM[35359] <= 32'b00000000111000111000001110110011;
ROM[35360] <= 32'b00000000011100010010000000100011;
ROM[35361] <= 32'b00000000010000010000000100010011;
ROM[35362] <= 32'b00000000001100010010000000100011;
ROM[35363] <= 32'b00000000010000010000000100010011;
ROM[35364] <= 32'b00000000010000010010000000100011;
ROM[35365] <= 32'b00000000010000010000000100010011;
ROM[35366] <= 32'b00000000010100010010000000100011;
ROM[35367] <= 32'b00000000010000010000000100010011;
ROM[35368] <= 32'b00000000011000010010000000100011;
ROM[35369] <= 32'b00000000010000010000000100010011;
ROM[35370] <= 32'b00000001010000000000001110010011;
ROM[35371] <= 32'b00000000010000111000001110010011;
ROM[35372] <= 32'b01000000011100010000001110110011;
ROM[35373] <= 32'b00000000011100000000001000110011;
ROM[35374] <= 32'b00000000001000000000000110110011;
ROM[35375] <= 32'b11101100000111111101000011101111;
ROM[35376] <= 32'b00000000001100000000001110010011;
ROM[35377] <= 32'b00000000011100010010000000100011;
ROM[35378] <= 32'b00000000010000010000000100010011;
ROM[35379] <= 32'b11111111110000010000000100010011;
ROM[35380] <= 32'b00000000000000010010001110000011;
ROM[35381] <= 32'b11111111110000010000000100010011;
ROM[35382] <= 32'b00000000000000010010010000000011;
ROM[35383] <= 32'b00000000011101000010010010110011;
ROM[35384] <= 32'b00000000100000111010010100110011;
ROM[35385] <= 32'b00000000101001001000001110110011;
ROM[35386] <= 32'b00000000000100111000001110010011;
ROM[35387] <= 32'b00000000000100111111001110010011;
ROM[35388] <= 32'b00000000011100010010000000100011;
ROM[35389] <= 32'b00000000010000010000000100010011;
ROM[35390] <= 32'b11111111110000010000000100010011;
ROM[35391] <= 32'b00000000000000010010001110000011;
ROM[35392] <= 32'b00000000000000111000101001100011;
ROM[35393] <= 32'b00000000000000100011001110110111;
ROM[35394] <= 32'b10010001100000111000001110010011;
ROM[35395] <= 32'b00000000111000111000001110110011;
ROM[35396] <= 32'b00000000000000111000000011100111;
ROM[35397] <= 32'b00000111100000000000000011101111;
ROM[35398] <= 32'b00000000110100101000010000110011;
ROM[35399] <= 32'b00000000000001000010001110000011;
ROM[35400] <= 32'b00000000011100010010000000100011;
ROM[35401] <= 32'b00000000010000010000000100010011;
ROM[35402] <= 32'b00000000000100000000001110010011;
ROM[35403] <= 32'b00000000011100010010000000100011;
ROM[35404] <= 32'b00000000010000010000000100010011;
ROM[35405] <= 32'b00000000000000100011001110110111;
ROM[35406] <= 32'b10011000000000111000001110010011;
ROM[35407] <= 32'b00000000111000111000001110110011;
ROM[35408] <= 32'b00000000011100010010000000100011;
ROM[35409] <= 32'b00000000010000010000000100010011;
ROM[35410] <= 32'b00000000001100010010000000100011;
ROM[35411] <= 32'b00000000010000010000000100010011;
ROM[35412] <= 32'b00000000010000010010000000100011;
ROM[35413] <= 32'b00000000010000010000000100010011;
ROM[35414] <= 32'b00000000010100010010000000100011;
ROM[35415] <= 32'b00000000010000010000000100010011;
ROM[35416] <= 32'b00000000011000010010000000100011;
ROM[35417] <= 32'b00000000010000010000000100010011;
ROM[35418] <= 32'b00000001010000000000001110010011;
ROM[35419] <= 32'b00000000100000111000001110010011;
ROM[35420] <= 32'b01000000011100010000001110110011;
ROM[35421] <= 32'b00000000011100000000001000110011;
ROM[35422] <= 32'b00000000001000000000000110110011;
ROM[35423] <= 32'b11100110000111111101000011101111;
ROM[35424] <= 32'b11111111110000010000000100010011;
ROM[35425] <= 32'b00000000000000010010001110000011;
ROM[35426] <= 32'b00000000011101100010000000100011;
ROM[35427] <= 32'b00000000110100101000010000110011;
ROM[35428] <= 32'b00000000000001000010001110000011;
ROM[35429] <= 32'b00000000011100010010000000100011;
ROM[35430] <= 32'b00000000010000010000000100010011;
ROM[35431] <= 32'b00000000000000100011001110110111;
ROM[35432] <= 32'b10011110100000111000001110010011;
ROM[35433] <= 32'b00000000111000111000001110110011;
ROM[35434] <= 32'b00000000011100010010000000100011;
ROM[35435] <= 32'b00000000010000010000000100010011;
ROM[35436] <= 32'b00000000001100010010000000100011;
ROM[35437] <= 32'b00000000010000010000000100010011;
ROM[35438] <= 32'b00000000010000010010000000100011;
ROM[35439] <= 32'b00000000010000010000000100010011;
ROM[35440] <= 32'b00000000010100010010000000100011;
ROM[35441] <= 32'b00000000010000010000000100010011;
ROM[35442] <= 32'b00000000011000010010000000100011;
ROM[35443] <= 32'b00000000010000010000000100010011;
ROM[35444] <= 32'b00000001010000000000001110010011;
ROM[35445] <= 32'b00000000010000111000001110010011;
ROM[35446] <= 32'b01000000011100010000001110110011;
ROM[35447] <= 32'b00000000011100000000001000110011;
ROM[35448] <= 32'b00000000001000000000000110110011;
ROM[35449] <= 32'b11011001100111111101000011101111;
ROM[35450] <= 32'b00000000010000000000001110010011;
ROM[35451] <= 32'b00000000011100010010000000100011;
ROM[35452] <= 32'b00000000010000010000000100010011;
ROM[35453] <= 32'b11111111110000010000000100010011;
ROM[35454] <= 32'b00000000000000010010001110000011;
ROM[35455] <= 32'b11111111110000010000000100010011;
ROM[35456] <= 32'b00000000000000010010010000000011;
ROM[35457] <= 32'b00000000011101000010010010110011;
ROM[35458] <= 32'b00000000100000111010010100110011;
ROM[35459] <= 32'b00000000101001001000001110110011;
ROM[35460] <= 32'b00000000000100111000001110010011;
ROM[35461] <= 32'b00000000000100111111001110010011;
ROM[35462] <= 32'b00000000011100010010000000100011;
ROM[35463] <= 32'b00000000010000010000000100010011;
ROM[35464] <= 32'b11111111110000010000000100010011;
ROM[35465] <= 32'b00000000000000010010001110000011;
ROM[35466] <= 32'b00000000000000111000101001100011;
ROM[35467] <= 32'b00000000000000100011001110110111;
ROM[35468] <= 32'b10100100000000111000001110010011;
ROM[35469] <= 32'b00000000111000111000001110110011;
ROM[35470] <= 32'b00000000000000111000000011100111;
ROM[35471] <= 32'b00000111100000000000000011101111;
ROM[35472] <= 32'b00000000110100101000010000110011;
ROM[35473] <= 32'b00000000000001000010001110000011;
ROM[35474] <= 32'b00000000011100010010000000100011;
ROM[35475] <= 32'b00000000010000010000000100010011;
ROM[35476] <= 32'b00000000000100000000001110010011;
ROM[35477] <= 32'b00000000011100010010000000100011;
ROM[35478] <= 32'b00000000010000010000000100010011;
ROM[35479] <= 32'b00000000000000100011001110110111;
ROM[35480] <= 32'b10101010100000111000001110010011;
ROM[35481] <= 32'b00000000111000111000001110110011;
ROM[35482] <= 32'b00000000011100010010000000100011;
ROM[35483] <= 32'b00000000010000010000000100010011;
ROM[35484] <= 32'b00000000001100010010000000100011;
ROM[35485] <= 32'b00000000010000010000000100010011;
ROM[35486] <= 32'b00000000010000010010000000100011;
ROM[35487] <= 32'b00000000010000010000000100010011;
ROM[35488] <= 32'b00000000010100010010000000100011;
ROM[35489] <= 32'b00000000010000010000000100010011;
ROM[35490] <= 32'b00000000011000010010000000100011;
ROM[35491] <= 32'b00000000010000010000000100010011;
ROM[35492] <= 32'b00000001010000000000001110010011;
ROM[35493] <= 32'b00000000100000111000001110010011;
ROM[35494] <= 32'b01000000011100010000001110110011;
ROM[35495] <= 32'b00000000011100000000001000110011;
ROM[35496] <= 32'b00000000001000000000000110110011;
ROM[35497] <= 32'b11010011100111111101000011101111;
ROM[35498] <= 32'b11111111110000010000000100010011;
ROM[35499] <= 32'b00000000000000010010001110000011;
ROM[35500] <= 32'b00000000011101100010000000100011;
ROM[35501] <= 32'b00000000100000011010001110000011;
ROM[35502] <= 32'b00000000011100010010000000100011;
ROM[35503] <= 32'b00000000010000010000000100010011;
ROM[35504] <= 32'b00001000010000000000001110010011;
ROM[35505] <= 32'b00000000011100010010000000100011;
ROM[35506] <= 32'b00000000010000010000000100010011;
ROM[35507] <= 32'b11111111110000010000000100010011;
ROM[35508] <= 32'b00000000000000010010001110000011;
ROM[35509] <= 32'b11111111110000010000000100010011;
ROM[35510] <= 32'b00000000000000010010010000000011;
ROM[35511] <= 32'b00000000011101000010010010110011;
ROM[35512] <= 32'b00000000100000111010010100110011;
ROM[35513] <= 32'b00000000101001001000001110110011;
ROM[35514] <= 32'b00000000000100111000001110010011;
ROM[35515] <= 32'b00000000000100111111001110010011;
ROM[35516] <= 32'b00000000011100010010000000100011;
ROM[35517] <= 32'b00000000010000010000000100010011;
ROM[35518] <= 32'b11111111110000010000000100010011;
ROM[35519] <= 32'b00000000000000010010001110000011;
ROM[35520] <= 32'b00000000000000111000101001100011;
ROM[35521] <= 32'b00000000000000100011001110110111;
ROM[35522] <= 32'b10110001100000111000001110010011;
ROM[35523] <= 32'b00000000111000111000001110110011;
ROM[35524] <= 32'b00000000000000111000000011100111;
ROM[35525] <= 32'b00100101010000000000000011101111;
ROM[35526] <= 32'b00000000110100101000010000110011;
ROM[35527] <= 32'b00000000000001000010001110000011;
ROM[35528] <= 32'b00000000011100010010000000100011;
ROM[35529] <= 32'b00000000010000010000000100010011;
ROM[35530] <= 32'b00000000000000100011001110110111;
ROM[35531] <= 32'b10110111010000111000001110010011;
ROM[35532] <= 32'b00000000111000111000001110110011;
ROM[35533] <= 32'b00000000011100010010000000100011;
ROM[35534] <= 32'b00000000010000010000000100010011;
ROM[35535] <= 32'b00000000001100010010000000100011;
ROM[35536] <= 32'b00000000010000010000000100010011;
ROM[35537] <= 32'b00000000010000010010000000100011;
ROM[35538] <= 32'b00000000010000010000000100010011;
ROM[35539] <= 32'b00000000010100010010000000100011;
ROM[35540] <= 32'b00000000010000010000000100010011;
ROM[35541] <= 32'b00000000011000010010000000100011;
ROM[35542] <= 32'b00000000010000010000000100010011;
ROM[35543] <= 32'b00000001010000000000001110010011;
ROM[35544] <= 32'b00000000010000111000001110010011;
ROM[35545] <= 32'b01000000011100010000001110110011;
ROM[35546] <= 32'b00000000011100000000001000110011;
ROM[35547] <= 32'b00000000001000000000000110110011;
ROM[35548] <= 32'b11000000110111111101000011101111;
ROM[35549] <= 32'b00000000000100000000001110010011;
ROM[35550] <= 32'b00000000011100010010000000100011;
ROM[35551] <= 32'b00000000010000010000000100010011;
ROM[35552] <= 32'b11111111110000010000000100010011;
ROM[35553] <= 32'b00000000000000010010001110000011;
ROM[35554] <= 32'b11111111110000010000000100010011;
ROM[35555] <= 32'b00000000000000010010010000000011;
ROM[35556] <= 32'b00000000011101000010010010110011;
ROM[35557] <= 32'b00000000100000111010010100110011;
ROM[35558] <= 32'b00000000101001001000001110110011;
ROM[35559] <= 32'b00000000000100111000001110010011;
ROM[35560] <= 32'b00000000000100111111001110010011;
ROM[35561] <= 32'b00000000011100010010000000100011;
ROM[35562] <= 32'b00000000010000010000000100010011;
ROM[35563] <= 32'b11111111110000010000000100010011;
ROM[35564] <= 32'b00000000000000010010001110000011;
ROM[35565] <= 32'b00000000000000111000101001100011;
ROM[35566] <= 32'b00000000000000100011001110110111;
ROM[35567] <= 32'b10111100110000111000001110010011;
ROM[35568] <= 32'b00000000111000111000001110110011;
ROM[35569] <= 32'b00000000000000111000000011100111;
ROM[35570] <= 32'b00000111100000000000000011101111;
ROM[35571] <= 32'b00000000110100101000010000110011;
ROM[35572] <= 32'b00000000000001000010001110000011;
ROM[35573] <= 32'b00000000011100010010000000100011;
ROM[35574] <= 32'b00000000010000010000000100010011;
ROM[35575] <= 32'b00000000010000000000001110010011;
ROM[35576] <= 32'b00000000011100010010000000100011;
ROM[35577] <= 32'b00000000010000010000000100010011;
ROM[35578] <= 32'b00000000000000100011001110110111;
ROM[35579] <= 32'b11000011010000111000001110010011;
ROM[35580] <= 32'b00000000111000111000001110110011;
ROM[35581] <= 32'b00000000011100010010000000100011;
ROM[35582] <= 32'b00000000010000010000000100010011;
ROM[35583] <= 32'b00000000001100010010000000100011;
ROM[35584] <= 32'b00000000010000010000000100010011;
ROM[35585] <= 32'b00000000010000010010000000100011;
ROM[35586] <= 32'b00000000010000010000000100010011;
ROM[35587] <= 32'b00000000010100010010000000100011;
ROM[35588] <= 32'b00000000010000010000000100010011;
ROM[35589] <= 32'b00000000011000010010000000100011;
ROM[35590] <= 32'b00000000010000010000000100010011;
ROM[35591] <= 32'b00000001010000000000001110010011;
ROM[35592] <= 32'b00000000100000111000001110010011;
ROM[35593] <= 32'b01000000011100010000001110110011;
ROM[35594] <= 32'b00000000011100000000001000110011;
ROM[35595] <= 32'b00000000001000000000000110110011;
ROM[35596] <= 32'b10111010110111111101000011101111;
ROM[35597] <= 32'b11111111110000010000000100010011;
ROM[35598] <= 32'b00000000000000010010001110000011;
ROM[35599] <= 32'b00000000011101100010000000100011;
ROM[35600] <= 32'b00000000110100101000010000110011;
ROM[35601] <= 32'b00000000000001000010001110000011;
ROM[35602] <= 32'b00000000011100010010000000100011;
ROM[35603] <= 32'b00000000010000010000000100010011;
ROM[35604] <= 32'b00000000000000100011001110110111;
ROM[35605] <= 32'b11001001110000111000001110010011;
ROM[35606] <= 32'b00000000111000111000001110110011;
ROM[35607] <= 32'b00000000011100010010000000100011;
ROM[35608] <= 32'b00000000010000010000000100010011;
ROM[35609] <= 32'b00000000001100010010000000100011;
ROM[35610] <= 32'b00000000010000010000000100010011;
ROM[35611] <= 32'b00000000010000010010000000100011;
ROM[35612] <= 32'b00000000010000010000000100010011;
ROM[35613] <= 32'b00000000010100010010000000100011;
ROM[35614] <= 32'b00000000010000010000000100010011;
ROM[35615] <= 32'b00000000011000010010000000100011;
ROM[35616] <= 32'b00000000010000010000000100010011;
ROM[35617] <= 32'b00000001010000000000001110010011;
ROM[35618] <= 32'b00000000010000111000001110010011;
ROM[35619] <= 32'b01000000011100010000001110110011;
ROM[35620] <= 32'b00000000011100000000001000110011;
ROM[35621] <= 32'b00000000001000000000000110110011;
ROM[35622] <= 32'b10101110010111111101000011101111;
ROM[35623] <= 32'b00000000001000000000001110010011;
ROM[35624] <= 32'b00000000011100010010000000100011;
ROM[35625] <= 32'b00000000010000010000000100010011;
ROM[35626] <= 32'b11111111110000010000000100010011;
ROM[35627] <= 32'b00000000000000010010001110000011;
ROM[35628] <= 32'b11111111110000010000000100010011;
ROM[35629] <= 32'b00000000000000010010010000000011;
ROM[35630] <= 32'b00000000011101000010010010110011;
ROM[35631] <= 32'b00000000100000111010010100110011;
ROM[35632] <= 32'b00000000101001001000001110110011;
ROM[35633] <= 32'b00000000000100111000001110010011;
ROM[35634] <= 32'b00000000000100111111001110010011;
ROM[35635] <= 32'b00000000011100010010000000100011;
ROM[35636] <= 32'b00000000010000010000000100010011;
ROM[35637] <= 32'b11111111110000010000000100010011;
ROM[35638] <= 32'b00000000000000010010001110000011;
ROM[35639] <= 32'b00000000000000111000101001100011;
ROM[35640] <= 32'b00000000000000100011001110110111;
ROM[35641] <= 32'b11001111010000111000001110010011;
ROM[35642] <= 32'b00000000111000111000001110110011;
ROM[35643] <= 32'b00000000000000111000000011100111;
ROM[35644] <= 32'b00000111100000000000000011101111;
ROM[35645] <= 32'b00000000110100101000010000110011;
ROM[35646] <= 32'b00000000000001000010001110000011;
ROM[35647] <= 32'b00000000011100010010000000100011;
ROM[35648] <= 32'b00000000010000010000000100010011;
ROM[35649] <= 32'b00000000010000000000001110010011;
ROM[35650] <= 32'b00000000011100010010000000100011;
ROM[35651] <= 32'b00000000010000010000000100010011;
ROM[35652] <= 32'b00000000000000100011001110110111;
ROM[35653] <= 32'b11010101110000111000001110010011;
ROM[35654] <= 32'b00000000111000111000001110110011;
ROM[35655] <= 32'b00000000011100010010000000100011;
ROM[35656] <= 32'b00000000010000010000000100010011;
ROM[35657] <= 32'b00000000001100010010000000100011;
ROM[35658] <= 32'b00000000010000010000000100010011;
ROM[35659] <= 32'b00000000010000010010000000100011;
ROM[35660] <= 32'b00000000010000010000000100010011;
ROM[35661] <= 32'b00000000010100010010000000100011;
ROM[35662] <= 32'b00000000010000010000000100010011;
ROM[35663] <= 32'b00000000011000010010000000100011;
ROM[35664] <= 32'b00000000010000010000000100010011;
ROM[35665] <= 32'b00000001010000000000001110010011;
ROM[35666] <= 32'b00000000100000111000001110010011;
ROM[35667] <= 32'b01000000011100010000001110110011;
ROM[35668] <= 32'b00000000011100000000001000110011;
ROM[35669] <= 32'b00000000001000000000000110110011;
ROM[35670] <= 32'b10101000010111111101000011101111;
ROM[35671] <= 32'b11111111110000010000000100010011;
ROM[35672] <= 32'b00000000000000010010001110000011;
ROM[35673] <= 32'b00000000011101100010000000100011;
ROM[35674] <= 32'b00000000100000011010001110000011;
ROM[35675] <= 32'b00000000011100010010000000100011;
ROM[35676] <= 32'b00000000010000010000000100010011;
ROM[35677] <= 32'b00001000010100000000001110010011;
ROM[35678] <= 32'b00000000011100010010000000100011;
ROM[35679] <= 32'b00000000010000010000000100010011;
ROM[35680] <= 32'b11111111110000010000000100010011;
ROM[35681] <= 32'b00000000000000010010001110000011;
ROM[35682] <= 32'b11111111110000010000000100010011;
ROM[35683] <= 32'b00000000000000010010010000000011;
ROM[35684] <= 32'b00000000011101000010010010110011;
ROM[35685] <= 32'b00000000100000111010010100110011;
ROM[35686] <= 32'b00000000101001001000001110110011;
ROM[35687] <= 32'b00000000000100111000001110010011;
ROM[35688] <= 32'b00000000000100111111001110010011;
ROM[35689] <= 32'b00000000011100010010000000100011;
ROM[35690] <= 32'b00000000010000010000000100010011;
ROM[35691] <= 32'b11111111110000010000000100010011;
ROM[35692] <= 32'b00000000000000010010001110000011;
ROM[35693] <= 32'b00000000000000111000101001100011;
ROM[35694] <= 32'b00000000000000100011001110110111;
ROM[35695] <= 32'b11011100110000111000001110010011;
ROM[35696] <= 32'b00000000111000111000001110110011;
ROM[35697] <= 32'b00000000000000111000000011100111;
ROM[35698] <= 32'b00100101010000000000000011101111;
ROM[35699] <= 32'b00000000110100101000010000110011;
ROM[35700] <= 32'b00000000000001000010001110000011;
ROM[35701] <= 32'b00000000011100010010000000100011;
ROM[35702] <= 32'b00000000010000010000000100010011;
ROM[35703] <= 32'b00000000000000100011001110110111;
ROM[35704] <= 32'b11100010100000111000001110010011;
ROM[35705] <= 32'b00000000111000111000001110110011;
ROM[35706] <= 32'b00000000011100010010000000100011;
ROM[35707] <= 32'b00000000010000010000000100010011;
ROM[35708] <= 32'b00000000001100010010000000100011;
ROM[35709] <= 32'b00000000010000010000000100010011;
ROM[35710] <= 32'b00000000010000010010000000100011;
ROM[35711] <= 32'b00000000010000010000000100010011;
ROM[35712] <= 32'b00000000010100010010000000100011;
ROM[35713] <= 32'b00000000010000010000000100010011;
ROM[35714] <= 32'b00000000011000010010000000100011;
ROM[35715] <= 32'b00000000010000010000000100010011;
ROM[35716] <= 32'b00000001010000000000001110010011;
ROM[35717] <= 32'b00000000010000111000001110010011;
ROM[35718] <= 32'b01000000011100010000001110110011;
ROM[35719] <= 32'b00000000011100000000001000110011;
ROM[35720] <= 32'b00000000001000000000000110110011;
ROM[35721] <= 32'b10010101100111111101000011101111;
ROM[35722] <= 32'b00000000001100000000001110010011;
ROM[35723] <= 32'b00000000011100010010000000100011;
ROM[35724] <= 32'b00000000010000010000000100010011;
ROM[35725] <= 32'b11111111110000010000000100010011;
ROM[35726] <= 32'b00000000000000010010001110000011;
ROM[35727] <= 32'b11111111110000010000000100010011;
ROM[35728] <= 32'b00000000000000010010010000000011;
ROM[35729] <= 32'b00000000011101000010010010110011;
ROM[35730] <= 32'b00000000100000111010010100110011;
ROM[35731] <= 32'b00000000101001001000001110110011;
ROM[35732] <= 32'b00000000000100111000001110010011;
ROM[35733] <= 32'b00000000000100111111001110010011;
ROM[35734] <= 32'b00000000011100010010000000100011;
ROM[35735] <= 32'b00000000010000010000000100010011;
ROM[35736] <= 32'b11111111110000010000000100010011;
ROM[35737] <= 32'b00000000000000010010001110000011;
ROM[35738] <= 32'b00000000000000111000101001100011;
ROM[35739] <= 32'b00000000000000100011001110110111;
ROM[35740] <= 32'b11101000000000111000001110010011;
ROM[35741] <= 32'b00000000111000111000001110110011;
ROM[35742] <= 32'b00000000000000111000000011100111;
ROM[35743] <= 32'b00000111100000000000000011101111;
ROM[35744] <= 32'b00000000110100101000010000110011;
ROM[35745] <= 32'b00000000000001000010001110000011;
ROM[35746] <= 32'b00000000011100010010000000100011;
ROM[35747] <= 32'b00000000010000010000000100010011;
ROM[35748] <= 32'b00000000001000000000001110010011;
ROM[35749] <= 32'b00000000011100010010000000100011;
ROM[35750] <= 32'b00000000010000010000000100010011;
ROM[35751] <= 32'b00000000000000100011001110110111;
ROM[35752] <= 32'b11101110100000111000001110010011;
ROM[35753] <= 32'b00000000111000111000001110110011;
ROM[35754] <= 32'b00000000011100010010000000100011;
ROM[35755] <= 32'b00000000010000010000000100010011;
ROM[35756] <= 32'b00000000001100010010000000100011;
ROM[35757] <= 32'b00000000010000010000000100010011;
ROM[35758] <= 32'b00000000010000010010000000100011;
ROM[35759] <= 32'b00000000010000010000000100010011;
ROM[35760] <= 32'b00000000010100010010000000100011;
ROM[35761] <= 32'b00000000010000010000000100010011;
ROM[35762] <= 32'b00000000011000010010000000100011;
ROM[35763] <= 32'b00000000010000010000000100010011;
ROM[35764] <= 32'b00000001010000000000001110010011;
ROM[35765] <= 32'b00000000100000111000001110010011;
ROM[35766] <= 32'b01000000011100010000001110110011;
ROM[35767] <= 32'b00000000011100000000001000110011;
ROM[35768] <= 32'b00000000001000000000000110110011;
ROM[35769] <= 32'b10001111100111111101000011101111;
ROM[35770] <= 32'b11111111110000010000000100010011;
ROM[35771] <= 32'b00000000000000010010001110000011;
ROM[35772] <= 32'b00000000011101100010000000100011;
ROM[35773] <= 32'b00000000110100101000010000110011;
ROM[35774] <= 32'b00000000000001000010001110000011;
ROM[35775] <= 32'b00000000011100010010000000100011;
ROM[35776] <= 32'b00000000010000010000000100010011;
ROM[35777] <= 32'b00000000000000100011001110110111;
ROM[35778] <= 32'b11110101000000111000001110010011;
ROM[35779] <= 32'b00000000111000111000001110110011;
ROM[35780] <= 32'b00000000011100010010000000100011;
ROM[35781] <= 32'b00000000010000010000000100010011;
ROM[35782] <= 32'b00000000001100010010000000100011;
ROM[35783] <= 32'b00000000010000010000000100010011;
ROM[35784] <= 32'b00000000010000010010000000100011;
ROM[35785] <= 32'b00000000010000010000000100010011;
ROM[35786] <= 32'b00000000010100010010000000100011;
ROM[35787] <= 32'b00000000010000010000000100010011;
ROM[35788] <= 32'b00000000011000010010000000100011;
ROM[35789] <= 32'b00000000010000010000000100010011;
ROM[35790] <= 32'b00000001010000000000001110010011;
ROM[35791] <= 32'b00000000010000111000001110010011;
ROM[35792] <= 32'b01000000011100010000001110110011;
ROM[35793] <= 32'b00000000011100000000001000110011;
ROM[35794] <= 32'b00000000001000000000000110110011;
ROM[35795] <= 32'b10000011000111111101000011101111;
ROM[35796] <= 32'b00000000010000000000001110010011;
ROM[35797] <= 32'b00000000011100010010000000100011;
ROM[35798] <= 32'b00000000010000010000000100010011;
ROM[35799] <= 32'b11111111110000010000000100010011;
ROM[35800] <= 32'b00000000000000010010001110000011;
ROM[35801] <= 32'b11111111110000010000000100010011;
ROM[35802] <= 32'b00000000000000010010010000000011;
ROM[35803] <= 32'b00000000011101000010010010110011;
ROM[35804] <= 32'b00000000100000111010010100110011;
ROM[35805] <= 32'b00000000101001001000001110110011;
ROM[35806] <= 32'b00000000000100111000001110010011;
ROM[35807] <= 32'b00000000000100111111001110010011;
ROM[35808] <= 32'b00000000011100010010000000100011;
ROM[35809] <= 32'b00000000010000010000000100010011;
ROM[35810] <= 32'b11111111110000010000000100010011;
ROM[35811] <= 32'b00000000000000010010001110000011;
ROM[35812] <= 32'b00000000000000111000101001100011;
ROM[35813] <= 32'b00000000000000100011001110110111;
ROM[35814] <= 32'b11111010100000111000001110010011;
ROM[35815] <= 32'b00000000111000111000001110110011;
ROM[35816] <= 32'b00000000000000111000000011100111;
ROM[35817] <= 32'b00000111100000000000000011101111;
ROM[35818] <= 32'b00000000110100101000010000110011;
ROM[35819] <= 32'b00000000000001000010001110000011;
ROM[35820] <= 32'b00000000011100010010000000100011;
ROM[35821] <= 32'b00000000010000010000000100010011;
ROM[35822] <= 32'b00000000001000000000001110010011;
ROM[35823] <= 32'b00000000011100010010000000100011;
ROM[35824] <= 32'b00000000010000010000000100010011;
ROM[35825] <= 32'b00000000000000100011001110110111;
ROM[35826] <= 32'b00000001000000111000001110010011;
ROM[35827] <= 32'b00000000111000111000001110110011;
ROM[35828] <= 32'b00000000011100010010000000100011;
ROM[35829] <= 32'b00000000010000010000000100010011;
ROM[35830] <= 32'b00000000001100010010000000100011;
ROM[35831] <= 32'b00000000010000010000000100010011;
ROM[35832] <= 32'b00000000010000010010000000100011;
ROM[35833] <= 32'b00000000010000010000000100010011;
ROM[35834] <= 32'b00000000010100010010000000100011;
ROM[35835] <= 32'b00000000010000010000000100010011;
ROM[35836] <= 32'b00000000011000010010000000100011;
ROM[35837] <= 32'b00000000010000010000000100010011;
ROM[35838] <= 32'b00000001010000000000001110010011;
ROM[35839] <= 32'b00000000100000111000001110010011;
ROM[35840] <= 32'b01000000011100010000001110110011;
ROM[35841] <= 32'b00000000011100000000001000110011;
ROM[35842] <= 32'b00000000001000000000000110110011;
ROM[35843] <= 32'b11111101000011111101000011101111;
ROM[35844] <= 32'b11111111110000010000000100010011;
ROM[35845] <= 32'b00000000000000010010001110000011;
ROM[35846] <= 32'b00000000011101100010000000100011;
ROM[35847] <= 32'b00000000110100101000010000110011;
ROM[35848] <= 32'b00000000000001000010001110000011;
ROM[35849] <= 32'b00000000011100010010000000100011;
ROM[35850] <= 32'b00000000010000010000000100010011;
ROM[35851] <= 32'b00000000000000100011001110110111;
ROM[35852] <= 32'b00000111100000111000001110010011;
ROM[35853] <= 32'b00000000111000111000001110110011;
ROM[35854] <= 32'b00000000011100010010000000100011;
ROM[35855] <= 32'b00000000010000010000000100010011;
ROM[35856] <= 32'b00000000001100010010000000100011;
ROM[35857] <= 32'b00000000010000010000000100010011;
ROM[35858] <= 32'b00000000010000010010000000100011;
ROM[35859] <= 32'b00000000010000010000000100010011;
ROM[35860] <= 32'b00000000010100010010000000100011;
ROM[35861] <= 32'b00000000010000010000000100010011;
ROM[35862] <= 32'b00000000011000010010000000100011;
ROM[35863] <= 32'b00000000010000010000000100010011;
ROM[35864] <= 32'b00000001010000000000001110010011;
ROM[35865] <= 32'b00000000010000111000001110010011;
ROM[35866] <= 32'b01000000011100010000001110110011;
ROM[35867] <= 32'b00000000011100000000001000110011;
ROM[35868] <= 32'b00000000001000000000000110110011;
ROM[35869] <= 32'b10000101110111111101000011101111;
ROM[35870] <= 32'b11111111110000010000000100010011;
ROM[35871] <= 32'b00000000000000010010001110000011;
ROM[35872] <= 32'b01000000011100000000001110110011;
ROM[35873] <= 32'b00000000000100111000001110010011;
ROM[35874] <= 32'b00000000011100010010000000100011;
ROM[35875] <= 32'b00000000010000010000000100010011;
ROM[35876] <= 32'b11111111110000010000000100010011;
ROM[35877] <= 32'b00000000000000010010001110000011;
ROM[35878] <= 32'b00000000000000111000101001100011;
ROM[35879] <= 32'b00000000000000100011001110110111;
ROM[35880] <= 32'b00001011000000111000001110010011;
ROM[35881] <= 32'b00000000111000111000001110110011;
ROM[35882] <= 32'b00000000000000111000000011100111;
ROM[35883] <= 32'b00001100010000000000000011101111;
ROM[35884] <= 32'b00000000110100101000010000110011;
ROM[35885] <= 32'b00000000010001000010001110000011;
ROM[35886] <= 32'b00000000011100010010000000100011;
ROM[35887] <= 32'b00000000010000010000000100010011;
ROM[35888] <= 32'b00000000000000100011001110110111;
ROM[35889] <= 32'b00010000110000111000001110010011;
ROM[35890] <= 32'b00000000111000111000001110110011;
ROM[35891] <= 32'b00000000011100010010000000100011;
ROM[35892] <= 32'b00000000010000010000000100010011;
ROM[35893] <= 32'b00000000001100010010000000100011;
ROM[35894] <= 32'b00000000010000010000000100010011;
ROM[35895] <= 32'b00000000010000010010000000100011;
ROM[35896] <= 32'b00000000010000010000000100010011;
ROM[35897] <= 32'b00000000010100010010000000100011;
ROM[35898] <= 32'b00000000010000010000000100010011;
ROM[35899] <= 32'b00000000011000010010000000100011;
ROM[35900] <= 32'b00000000010000010000000100010011;
ROM[35901] <= 32'b00000001010000000000001110010011;
ROM[35902] <= 32'b00000000010000111000001110010011;
ROM[35903] <= 32'b01000000011100010000001110110011;
ROM[35904] <= 32'b00000000011100000000001000110011;
ROM[35905] <= 32'b00000000001000000000000110110011;
ROM[35906] <= 32'b00010001110000000110000011101111;
ROM[35907] <= 32'b11111111110000010000000100010011;
ROM[35908] <= 32'b00000000000000010010001110000011;
ROM[35909] <= 32'b00000000011101100010000000100011;
ROM[35910] <= 32'b00000000000000100011001110110111;
ROM[35911] <= 32'b00010110010000111000001110010011;
ROM[35912] <= 32'b00000000111000111000001110110011;
ROM[35913] <= 32'b00000000011100010010000000100011;
ROM[35914] <= 32'b00000000010000010000000100010011;
ROM[35915] <= 32'b00000000001100010010000000100011;
ROM[35916] <= 32'b00000000010000010000000100010011;
ROM[35917] <= 32'b00000000010000010010000000100011;
ROM[35918] <= 32'b00000000010000010000000100010011;
ROM[35919] <= 32'b00000000010100010010000000100011;
ROM[35920] <= 32'b00000000010000010000000100010011;
ROM[35921] <= 32'b00000000011000010010000000100011;
ROM[35922] <= 32'b00000000010000010000000100010011;
ROM[35923] <= 32'b00000001010000000000001110010011;
ROM[35924] <= 32'b00000000000000111000001110010011;
ROM[35925] <= 32'b01000000011100010000001110110011;
ROM[35926] <= 32'b00000000011100000000001000110011;
ROM[35927] <= 32'b00000000001000000000000110110011;
ROM[35928] <= 32'b01101100100100000111000011101111;
ROM[35929] <= 32'b11111111110000010000000100010011;
ROM[35930] <= 32'b00000000000000010010001110000011;
ROM[35931] <= 32'b00000000011101100010000000100011;
ROM[35932] <= 32'b00000000110100101000010000110011;
ROM[35933] <= 32'b00000000010001000010001110000011;
ROM[35934] <= 32'b00000000011100010010000000100011;
ROM[35935] <= 32'b00000000010000010000000100010011;
ROM[35936] <= 32'b00000000110100101000010000110011;
ROM[35937] <= 32'b00000000000001000010001110000011;
ROM[35938] <= 32'b00000000011100010010000000100011;
ROM[35939] <= 32'b00000000010000010000000100010011;
ROM[35940] <= 32'b00000000000000100011001110110111;
ROM[35941] <= 32'b00011101110000111000001110010011;
ROM[35942] <= 32'b00000000111000111000001110110011;
ROM[35943] <= 32'b00000000011100010010000000100011;
ROM[35944] <= 32'b00000000010000010000000100010011;
ROM[35945] <= 32'b00000000001100010010000000100011;
ROM[35946] <= 32'b00000000010000010000000100010011;
ROM[35947] <= 32'b00000000010000010010000000100011;
ROM[35948] <= 32'b00000000010000010000000100010011;
ROM[35949] <= 32'b00000000010100010010000000100011;
ROM[35950] <= 32'b00000000010000010000000100010011;
ROM[35951] <= 32'b00000000011000010010000000100011;
ROM[35952] <= 32'b00000000010000010000000100010011;
ROM[35953] <= 32'b00000001010000000000001110010011;
ROM[35954] <= 32'b00000000010000111000001110010011;
ROM[35955] <= 32'b01000000011100010000001110110011;
ROM[35956] <= 32'b00000000011100000000001000110011;
ROM[35957] <= 32'b00000000001000000000000110110011;
ROM[35958] <= 32'b11000010010011111101000011101111;
ROM[35959] <= 32'b00000000110100101000010000110011;
ROM[35960] <= 32'b00000000000001000010001110000011;
ROM[35961] <= 32'b00000000011100010010000000100011;
ROM[35962] <= 32'b00000000010000010000000100010011;
ROM[35963] <= 32'b00000000000000100011001110110111;
ROM[35964] <= 32'b00100011100000111000001110010011;
ROM[35965] <= 32'b00000000111000111000001110110011;
ROM[35966] <= 32'b00000000011100010010000000100011;
ROM[35967] <= 32'b00000000010000010000000100010011;
ROM[35968] <= 32'b00000000001100010010000000100011;
ROM[35969] <= 32'b00000000010000010000000100010011;
ROM[35970] <= 32'b00000000010000010010000000100011;
ROM[35971] <= 32'b00000000010000010000000100010011;
ROM[35972] <= 32'b00000000010100010010000000100011;
ROM[35973] <= 32'b00000000010000010000000100010011;
ROM[35974] <= 32'b00000000011000010010000000100011;
ROM[35975] <= 32'b00000000010000010000000100010011;
ROM[35976] <= 32'b00000001010000000000001110010011;
ROM[35977] <= 32'b00000000010000111000001110010011;
ROM[35978] <= 32'b01000000011100010000001110110011;
ROM[35979] <= 32'b00000000011100000000001000110011;
ROM[35980] <= 32'b00000000001000000000000110110011;
ROM[35981] <= 32'b11000010100011111101000011101111;
ROM[35982] <= 32'b00000000000000100011001110110111;
ROM[35983] <= 32'b00101000010000111000001110010011;
ROM[35984] <= 32'b00000000111000111000001110110011;
ROM[35985] <= 32'b00000000011100010010000000100011;
ROM[35986] <= 32'b00000000010000010000000100010011;
ROM[35987] <= 32'b00000000001100010010000000100011;
ROM[35988] <= 32'b00000000010000010000000100010011;
ROM[35989] <= 32'b00000000010000010010000000100011;
ROM[35990] <= 32'b00000000010000010000000100010011;
ROM[35991] <= 32'b00000000010100010010000000100011;
ROM[35992] <= 32'b00000000010000010000000100010011;
ROM[35993] <= 32'b00000000011000010010000000100011;
ROM[35994] <= 32'b00000000010000010000000100010011;
ROM[35995] <= 32'b00000001010000000000001110010011;
ROM[35996] <= 32'b00000000110000111000001110010011;
ROM[35997] <= 32'b01000000011100010000001110110011;
ROM[35998] <= 32'b00000000011100000000001000110011;
ROM[35999] <= 32'b00000000001000000000000110110011;
ROM[36000] <= 32'b00101010010000000011000011101111;
ROM[36001] <= 32'b11111111110000010000000100010011;
ROM[36002] <= 32'b00000000000000010010001110000011;
ROM[36003] <= 32'b00000000000000111000101001100011;
ROM[36004] <= 32'b00000000000000100011001110110111;
ROM[36005] <= 32'b00101010010000111000001110010011;
ROM[36006] <= 32'b00000000111000111000001110110011;
ROM[36007] <= 32'b00000000000000111000000011100111;
ROM[36008] <= 32'b00010011010000000000000011101111;
ROM[36009] <= 32'b00000000110100101000010000110011;
ROM[36010] <= 32'b00000000000001000010001110000011;
ROM[36011] <= 32'b00000000011100010010000000100011;
ROM[36012] <= 32'b00000000010000010000000100010011;
ROM[36013] <= 32'b00000000000000100011001110110111;
ROM[36014] <= 32'b00110000000000111000001110010011;
ROM[36015] <= 32'b00000000111000111000001110110011;
ROM[36016] <= 32'b00000000011100010010000000100011;
ROM[36017] <= 32'b00000000010000010000000100010011;
ROM[36018] <= 32'b00000000001100010010000000100011;
ROM[36019] <= 32'b00000000010000010000000100010011;
ROM[36020] <= 32'b00000000010000010010000000100011;
ROM[36021] <= 32'b00000000010000010000000100010011;
ROM[36022] <= 32'b00000000010100010010000000100011;
ROM[36023] <= 32'b00000000010000010000000100010011;
ROM[36024] <= 32'b00000000011000010010000000100011;
ROM[36025] <= 32'b00000000010000010000000100010011;
ROM[36026] <= 32'b00000001010000000000001110010011;
ROM[36027] <= 32'b00000000010000111000001110010011;
ROM[36028] <= 32'b01000000011100010000001110110011;
ROM[36029] <= 32'b00000000011100000000001000110011;
ROM[36030] <= 32'b00000000001000000000000110110011;
ROM[36031] <= 32'b11011001000011111110000011101111;
ROM[36032] <= 32'b11111111110000010000000100010011;
ROM[36033] <= 32'b00000000000000010010001110000011;
ROM[36034] <= 32'b00000000011101100010000000100011;
ROM[36035] <= 32'b00000000010100010010000000100011;
ROM[36036] <= 32'b00000000010000010000000100010011;
ROM[36037] <= 32'b00000000000000100011001110110111;
ROM[36038] <= 32'b00110110000000111000001110010011;
ROM[36039] <= 32'b00000000111000111000001110110011;
ROM[36040] <= 32'b00000000011100010010000000100011;
ROM[36041] <= 32'b00000000010000010000000100010011;
ROM[36042] <= 32'b00000000001100010010000000100011;
ROM[36043] <= 32'b00000000010000010000000100010011;
ROM[36044] <= 32'b00000000010000010010000000100011;
ROM[36045] <= 32'b00000000010000010000000100010011;
ROM[36046] <= 32'b00000000010100010010000000100011;
ROM[36047] <= 32'b00000000010000010000000100010011;
ROM[36048] <= 32'b00000000011000010010000000100011;
ROM[36049] <= 32'b00000000010000010000000100010011;
ROM[36050] <= 32'b00000001010000000000001110010011;
ROM[36051] <= 32'b00000000010000111000001110010011;
ROM[36052] <= 32'b01000000011100010000001110110011;
ROM[36053] <= 32'b00000000011100000000001000110011;
ROM[36054] <= 32'b00000000001000000000000110110011;
ROM[36055] <= 32'b01000111100000000000000011101111;
ROM[36056] <= 32'b11111111110000010000000100010011;
ROM[36057] <= 32'b00000000000000010010001110000011;
ROM[36058] <= 32'b00000000011101100010000000100011;
ROM[36059] <= 32'b00000000110100101000010000110011;
ROM[36060] <= 32'b00000000010001000010001110000011;
ROM[36061] <= 32'b00000000011100010010000000100011;
ROM[36062] <= 32'b00000000010000010000000100010011;
ROM[36063] <= 32'b00000000000000100011001110110111;
ROM[36064] <= 32'b00111100100000111000001110010011;
ROM[36065] <= 32'b00000000111000111000001110110011;
ROM[36066] <= 32'b00000000011100010010000000100011;
ROM[36067] <= 32'b00000000010000010000000100010011;
ROM[36068] <= 32'b00000000001100010010000000100011;
ROM[36069] <= 32'b00000000010000010000000100010011;
ROM[36070] <= 32'b00000000010000010010000000100011;
ROM[36071] <= 32'b00000000010000010000000100010011;
ROM[36072] <= 32'b00000000010100010010000000100011;
ROM[36073] <= 32'b00000000010000010000000100010011;
ROM[36074] <= 32'b00000000011000010010000000100011;
ROM[36075] <= 32'b00000000010000010000000100010011;
ROM[36076] <= 32'b00000001010000000000001110010011;
ROM[36077] <= 32'b00000000010000111000001110010011;
ROM[36078] <= 32'b01000000011100010000001110110011;
ROM[36079] <= 32'b00000000011100000000001000110011;
ROM[36080] <= 32'b00000000001000000000000110110011;
ROM[36081] <= 32'b01100111100100000001000011101111;
ROM[36082] <= 32'b11111111110000010000000100010011;
ROM[36083] <= 32'b00000000000000010010001110000011;
ROM[36084] <= 32'b00000000011101100010000000100011;
ROM[36085] <= 32'b00000000110100101000010000110011;
ROM[36086] <= 32'b00000000000001000010001110000011;
ROM[36087] <= 32'b00000000011100010010000000100011;
ROM[36088] <= 32'b00000000010000010000000100010011;
ROM[36089] <= 32'b00000000110100101000010000110011;
ROM[36090] <= 32'b00000001010001000010001110000011;
ROM[36091] <= 32'b00000000011100010010000000100011;
ROM[36092] <= 32'b00000000010000010000000100010011;
ROM[36093] <= 32'b00000000000000100011001110110111;
ROM[36094] <= 32'b01000100000000111000001110010011;
ROM[36095] <= 32'b00000000111000111000001110110011;
ROM[36096] <= 32'b00000000011100010010000000100011;
ROM[36097] <= 32'b00000000010000010000000100010011;
ROM[36098] <= 32'b00000000001100010010000000100011;
ROM[36099] <= 32'b00000000010000010000000100010011;
ROM[36100] <= 32'b00000000010000010010000000100011;
ROM[36101] <= 32'b00000000010000010000000100010011;
ROM[36102] <= 32'b00000000010100010010000000100011;
ROM[36103] <= 32'b00000000010000010000000100010011;
ROM[36104] <= 32'b00000000011000010010000000100011;
ROM[36105] <= 32'b00000000010000010000000100010011;
ROM[36106] <= 32'b00000001010000000000001110010011;
ROM[36107] <= 32'b00000000100000111000001110010011;
ROM[36108] <= 32'b01000000011100010000001110110011;
ROM[36109] <= 32'b00000000011100000000001000110011;
ROM[36110] <= 32'b00000000001000000000000110110011;
ROM[36111] <= 32'b11000101100111111101000011101111;
ROM[36112] <= 32'b11111111110000010000000100010011;
ROM[36113] <= 32'b00000000000000010010001110000011;
ROM[36114] <= 32'b00000000011101100010000000100011;
ROM[36115] <= 32'b00000000110100101000010000110011;
ROM[36116] <= 32'b00000000010001000010001110000011;
ROM[36117] <= 32'b00000000011100010010000000100011;
ROM[36118] <= 32'b00000000010000010000000100010011;
ROM[36119] <= 32'b00000000000000100011001110110111;
ROM[36120] <= 32'b01001010100000111000001110010011;
ROM[36121] <= 32'b00000000111000111000001110110011;
ROM[36122] <= 32'b00000000011100010010000000100011;
ROM[36123] <= 32'b00000000010000010000000100010011;
ROM[36124] <= 32'b00000000001100010010000000100011;
ROM[36125] <= 32'b00000000010000010000000100010011;
ROM[36126] <= 32'b00000000010000010010000000100011;
ROM[36127] <= 32'b00000000010000010000000100010011;
ROM[36128] <= 32'b00000000010100010010000000100011;
ROM[36129] <= 32'b00000000010000010000000100010011;
ROM[36130] <= 32'b00000000011000010010000000100011;
ROM[36131] <= 32'b00000000010000010000000100010011;
ROM[36132] <= 32'b00000001010000000000001110010011;
ROM[36133] <= 32'b00000000010000111000001110010011;
ROM[36134] <= 32'b01000000011100010000001110110011;
ROM[36135] <= 32'b00000000011100000000001000110011;
ROM[36136] <= 32'b00000000001000000000000110110011;
ROM[36137] <= 32'b00011100110000000010000011101111;
ROM[36138] <= 32'b11111111110000010000000100010011;
ROM[36139] <= 32'b00000000000000010010001110000011;
ROM[36140] <= 32'b00000000011101100010000000100011;
ROM[36141] <= 32'b00000000110100101000010000110011;
ROM[36142] <= 32'b00000000010001000010001110000011;
ROM[36143] <= 32'b00000000011100010010000000100011;
ROM[36144] <= 32'b00000000010000010000000100010011;
ROM[36145] <= 32'b00000000000000100011001110110111;
ROM[36146] <= 32'b01010001000000111000001110010011;
ROM[36147] <= 32'b00000000111000111000001110110011;
ROM[36148] <= 32'b00000000011100010010000000100011;
ROM[36149] <= 32'b00000000010000010000000100010011;
ROM[36150] <= 32'b00000000001100010010000000100011;
ROM[36151] <= 32'b00000000010000010000000100010011;
ROM[36152] <= 32'b00000000010000010010000000100011;
ROM[36153] <= 32'b00000000010000010000000100010011;
ROM[36154] <= 32'b00000000010100010010000000100011;
ROM[36155] <= 32'b00000000010000010000000100010011;
ROM[36156] <= 32'b00000000011000010010000000100011;
ROM[36157] <= 32'b00000000010000010000000100010011;
ROM[36158] <= 32'b00000001010000000000001110010011;
ROM[36159] <= 32'b00000000010000111000001110010011;
ROM[36160] <= 32'b01000000011100010000001110110011;
ROM[36161] <= 32'b00000000011100000000001000110011;
ROM[36162] <= 32'b00000000001000000000000110110011;
ROM[36163] <= 32'b00111110010100000011000011101111;
ROM[36164] <= 32'b11111111110000010000000100010011;
ROM[36165] <= 32'b00000000000000010010001110000011;
ROM[36166] <= 32'b00000000011101100010000000100011;
ROM[36167] <= 32'b00000000110100101000010000110011;
ROM[36168] <= 32'b00000001100001000010001110000011;
ROM[36169] <= 32'b00000000011100010010000000100011;
ROM[36170] <= 32'b00000000010000010000000100010011;
ROM[36171] <= 32'b00000000000000100011001110110111;
ROM[36172] <= 32'b01010111100000111000001110010011;
ROM[36173] <= 32'b00000000111000111000001110110011;
ROM[36174] <= 32'b00000000011100010010000000100011;
ROM[36175] <= 32'b00000000010000010000000100010011;
ROM[36176] <= 32'b00000000001100010010000000100011;
ROM[36177] <= 32'b00000000010000010000000100010011;
ROM[36178] <= 32'b00000000010000010010000000100011;
ROM[36179] <= 32'b00000000010000010000000100010011;
ROM[36180] <= 32'b00000000010100010010000000100011;
ROM[36181] <= 32'b00000000010000010000000100010011;
ROM[36182] <= 32'b00000000011000010010000000100011;
ROM[36183] <= 32'b00000000010000010000000100010011;
ROM[36184] <= 32'b00000001010000000000001110010011;
ROM[36185] <= 32'b00000000010000111000001110010011;
ROM[36186] <= 32'b01000000011100010000001110110011;
ROM[36187] <= 32'b00000000011100000000001000110011;
ROM[36188] <= 32'b00000000001000000000000110110011;
ROM[36189] <= 32'b00110101000100000111000011101111;
ROM[36190] <= 32'b11111111110000010000000100010011;
ROM[36191] <= 32'b00000000000000010010001110000011;
ROM[36192] <= 32'b00000000011101100010000000100011;
ROM[36193] <= 32'b00000000010100010010000000100011;
ROM[36194] <= 32'b00000000010000010000000100010011;
ROM[36195] <= 32'b00000000000000100011001110110111;
ROM[36196] <= 32'b01011101100000111000001110010011;
ROM[36197] <= 32'b00000000111000111000001110110011;
ROM[36198] <= 32'b00000000011100010010000000100011;
ROM[36199] <= 32'b00000000010000010000000100010011;
ROM[36200] <= 32'b00000000001100010010000000100011;
ROM[36201] <= 32'b00000000010000010000000100010011;
ROM[36202] <= 32'b00000000010000010010000000100011;
ROM[36203] <= 32'b00000000010000010000000100010011;
ROM[36204] <= 32'b00000000010100010010000000100011;
ROM[36205] <= 32'b00000000010000010000000100010011;
ROM[36206] <= 32'b00000000011000010010000000100011;
ROM[36207] <= 32'b00000000010000010000000100010011;
ROM[36208] <= 32'b00000001010000000000001110010011;
ROM[36209] <= 32'b00000000010000111000001110010011;
ROM[36210] <= 32'b01000000011100010000001110110011;
ROM[36211] <= 32'b00000000011100000000001000110011;
ROM[36212] <= 32'b00000000001000000000000110110011;
ROM[36213] <= 32'b00111110100000000000000011101111;
ROM[36214] <= 32'b11111111110000010000000100010011;
ROM[36215] <= 32'b00000000000000010010001110000011;
ROM[36216] <= 32'b00000000011101100010000000100011;
ROM[36217] <= 32'b00000000110100101000010000110011;
ROM[36218] <= 32'b00000000000001000010001110000011;
ROM[36219] <= 32'b00000000011100010010000000100011;
ROM[36220] <= 32'b00000000010000010000000100010011;
ROM[36221] <= 32'b00000000000000100011001110110111;
ROM[36222] <= 32'b01100100000000111000001110010011;
ROM[36223] <= 32'b00000000111000111000001110110011;
ROM[36224] <= 32'b00000000011100010010000000100011;
ROM[36225] <= 32'b00000000010000010000000100010011;
ROM[36226] <= 32'b00000000001100010010000000100011;
ROM[36227] <= 32'b00000000010000010000000100010011;
ROM[36228] <= 32'b00000000010000010010000000100011;
ROM[36229] <= 32'b00000000010000010000000100010011;
ROM[36230] <= 32'b00000000010100010010000000100011;
ROM[36231] <= 32'b00000000010000010000000100010011;
ROM[36232] <= 32'b00000000011000010010000000100011;
ROM[36233] <= 32'b00000000010000010000000100010011;
ROM[36234] <= 32'b00000001010000000000001110010011;
ROM[36235] <= 32'b00000000010000111000001110010011;
ROM[36236] <= 32'b01000000011100010000001110110011;
ROM[36237] <= 32'b00000000011100000000001000110011;
ROM[36238] <= 32'b00000000001000000000000110110011;
ROM[36239] <= 32'b10010010100111111100000011101111;
ROM[36240] <= 32'b11111111110000010000000100010011;
ROM[36241] <= 32'b00000000000000010010001110000011;
ROM[36242] <= 32'b00000000000000111000101001100011;
ROM[36243] <= 32'b00000000000000100011001110110111;
ROM[36244] <= 32'b01100110000000111000001110010011;
ROM[36245] <= 32'b00000000111000111000001110110011;
ROM[36246] <= 32'b00000000000000111000000011100111;
ROM[36247] <= 32'b00000111000000000000000011101111;
ROM[36248] <= 32'b00000000110100101000010000110011;
ROM[36249] <= 32'b00000000000001000010001110000011;
ROM[36250] <= 32'b00000000011100010010000000100011;
ROM[36251] <= 32'b00000000010000010000000100010011;
ROM[36252] <= 32'b00000000000000100011001110110111;
ROM[36253] <= 32'b01101011110000111000001110010011;
ROM[36254] <= 32'b00000000111000111000001110110011;
ROM[36255] <= 32'b00000000011100010010000000100011;
ROM[36256] <= 32'b00000000010000010000000100010011;
ROM[36257] <= 32'b00000000001100010010000000100011;
ROM[36258] <= 32'b00000000010000010000000100010011;
ROM[36259] <= 32'b00000000010000010010000000100011;
ROM[36260] <= 32'b00000000010000010000000100010011;
ROM[36261] <= 32'b00000000010100010010000000100011;
ROM[36262] <= 32'b00000000010000010000000100010011;
ROM[36263] <= 32'b00000000011000010010000000100011;
ROM[36264] <= 32'b00000000010000010000000100010011;
ROM[36265] <= 32'b00000001010000000000001110010011;
ROM[36266] <= 32'b00000000010000111000001110010011;
ROM[36267] <= 32'b01000000011100010000001110110011;
ROM[36268] <= 32'b00000000011100000000001000110011;
ROM[36269] <= 32'b00000000001000000000000110110011;
ROM[36270] <= 32'b10000000010011111101000011101111;
ROM[36271] <= 32'b11111111110000010000000100010011;
ROM[36272] <= 32'b00000000000000010010001110000011;
ROM[36273] <= 32'b00000000110100101000010000110011;
ROM[36274] <= 32'b00000000011101000010101000100011;
ROM[36275] <= 32'b10001001110111111110000011101111;
ROM[36276] <= 32'b00000000110100101000010000110011;
ROM[36277] <= 32'b00000000010001000010001110000011;
ROM[36278] <= 32'b00000000011100010010000000100011;
ROM[36279] <= 32'b00000000010000010000000100010011;
ROM[36280] <= 32'b00000000000000100011001110110111;
ROM[36281] <= 32'b01110010110000111000001110010011;
ROM[36282] <= 32'b00000000111000111000001110110011;
ROM[36283] <= 32'b00000000011100010010000000100011;
ROM[36284] <= 32'b00000000010000010000000100010011;
ROM[36285] <= 32'b00000000001100010010000000100011;
ROM[36286] <= 32'b00000000010000010000000100010011;
ROM[36287] <= 32'b00000000010000010010000000100011;
ROM[36288] <= 32'b00000000010000010000000100010011;
ROM[36289] <= 32'b00000000010100010010000000100011;
ROM[36290] <= 32'b00000000010000010000000100010011;
ROM[36291] <= 32'b00000000011000010010000000100011;
ROM[36292] <= 32'b00000000010000010000000100010011;
ROM[36293] <= 32'b00000001010000000000001110010011;
ROM[36294] <= 32'b00000000010000111000001110010011;
ROM[36295] <= 32'b01000000011100010000001110110011;
ROM[36296] <= 32'b00000000011100000000001000110011;
ROM[36297] <= 32'b00000000001000000000000110110011;
ROM[36298] <= 32'b01010011010000000101000011101111;
ROM[36299] <= 32'b11111111110000010000000100010011;
ROM[36300] <= 32'b00000000000000010010001110000011;
ROM[36301] <= 32'b00000000011101100010000000100011;
ROM[36302] <= 32'b00000000000000100011001110110111;
ROM[36303] <= 32'b01111000010000111000001110010011;
ROM[36304] <= 32'b00000000111000111000001110110011;
ROM[36305] <= 32'b00000000011100010010000000100011;
ROM[36306] <= 32'b00000000010000010000000100010011;
ROM[36307] <= 32'b00000000001100010010000000100011;
ROM[36308] <= 32'b00000000010000010000000100010011;
ROM[36309] <= 32'b00000000010000010010000000100011;
ROM[36310] <= 32'b00000000010000010000000100010011;
ROM[36311] <= 32'b00000000010100010010000000100011;
ROM[36312] <= 32'b00000000010000010000000100010011;
ROM[36313] <= 32'b00000000011000010010000000100011;
ROM[36314] <= 32'b00000000010000010000000100010011;
ROM[36315] <= 32'b00000001010000000000001110010011;
ROM[36316] <= 32'b00000000000000111000001110010011;
ROM[36317] <= 32'b01000000011100010000001110110011;
ROM[36318] <= 32'b00000000011100000000001000110011;
ROM[36319] <= 32'b00000000001000000000000110110011;
ROM[36320] <= 32'b00001010100100000111000011101111;
ROM[36321] <= 32'b11111111110000010000000100010011;
ROM[36322] <= 32'b00000000000000010010001110000011;
ROM[36323] <= 32'b00000000011101100010000000100011;
ROM[36324] <= 32'b00000000000000000000001110010011;
ROM[36325] <= 32'b00000000011100010010000000100011;
ROM[36326] <= 32'b00000000010000010000000100010011;
ROM[36327] <= 32'b00000001010000000000001110010011;
ROM[36328] <= 32'b01000000011100011000001110110011;
ROM[36329] <= 32'b00000000000000111010000010000011;
ROM[36330] <= 32'b11111111110000010000000100010011;
ROM[36331] <= 32'b00000000000000010010001110000011;
ROM[36332] <= 32'b00000000011100100010000000100011;
ROM[36333] <= 32'b00000000010000100000000100010011;
ROM[36334] <= 32'b00000001010000000000001110010011;
ROM[36335] <= 32'b01000000011100011000001110110011;
ROM[36336] <= 32'b00000000010000111010000110000011;
ROM[36337] <= 32'b00000000100000111010001000000011;
ROM[36338] <= 32'b00000000110000111010001010000011;
ROM[36339] <= 32'b00000001000000111010001100000011;
ROM[36340] <= 32'b00000000000000001000000011100111;
ROM[36341] <= 32'b00000000000000100010001110000011;
ROM[36342] <= 32'b00000000011100010010000000100011;
ROM[36343] <= 32'b00000000010000010000000100010011;
ROM[36344] <= 32'b11111111110000010000000100010011;
ROM[36345] <= 32'b00000000000000010010001110000011;
ROM[36346] <= 32'b00000000000000111000001010010011;
ROM[36347] <= 32'b00000000110100101000010000110011;
ROM[36348] <= 32'b00000000100001000010001110000011;
ROM[36349] <= 32'b00000000011100010010000000100011;
ROM[36350] <= 32'b00000000010000010000000100010011;
ROM[36351] <= 32'b00000000101000000000001110010011;
ROM[36352] <= 32'b00000000011100010010000000100011;
ROM[36353] <= 32'b00000000010000010000000100010011;
ROM[36354] <= 32'b00000000110100101000010000110011;
ROM[36355] <= 32'b00000000110001000010001110000011;
ROM[36356] <= 32'b00000000011100010010000000100011;
ROM[36357] <= 32'b00000000010000010000000100010011;
ROM[36358] <= 32'b00000000000000100100001110110111;
ROM[36359] <= 32'b10000110010000111000001110010011;
ROM[36360] <= 32'b00000000111000111000001110110011;
ROM[36361] <= 32'b00000000011100010010000000100011;
ROM[36362] <= 32'b00000000010000010000000100010011;
ROM[36363] <= 32'b00000000001100010010000000100011;
ROM[36364] <= 32'b00000000010000010000000100010011;
ROM[36365] <= 32'b00000000010000010010000000100011;
ROM[36366] <= 32'b00000000010000010000000100010011;
ROM[36367] <= 32'b00000000010100010010000000100011;
ROM[36368] <= 32'b00000000010000010000000100010011;
ROM[36369] <= 32'b00000000011000010010000000100011;
ROM[36370] <= 32'b00000000010000010000000100010011;
ROM[36371] <= 32'b00000001010000000000001110010011;
ROM[36372] <= 32'b00000000100000111000001110010011;
ROM[36373] <= 32'b01000000011100010000001110110011;
ROM[36374] <= 32'b00000000011100000000001000110011;
ROM[36375] <= 32'b00000000001000000000000110110011;
ROM[36376] <= 32'b11111100110111101101000011101111;
ROM[36377] <= 32'b11111111110000010000000100010011;
ROM[36378] <= 32'b00000000000000010010001110000011;
ROM[36379] <= 32'b11111111110000010000000100010011;
ROM[36380] <= 32'b00000000000000010010010000000011;
ROM[36381] <= 32'b00000000011101000000001110110011;
ROM[36382] <= 32'b00000000011100010010000000100011;
ROM[36383] <= 32'b00000000010000010000000100010011;
ROM[36384] <= 32'b11111111110000010000000100010011;
ROM[36385] <= 32'b00000000000000010010001110000011;
ROM[36386] <= 32'b00000000110100101000010000110011;
ROM[36387] <= 32'b00000000011101000010010000100011;
ROM[36388] <= 32'b00000000110100101000010000110011;
ROM[36389] <= 32'b00000000110001000010001110000011;
ROM[36390] <= 32'b00000000011100010010000000100011;
ROM[36391] <= 32'b00000000010000010000000100010011;
ROM[36392] <= 32'b00000000000100000000001110010011;
ROM[36393] <= 32'b00000000011100010010000000100011;
ROM[36394] <= 32'b00000000010000010000000100010011;
ROM[36395] <= 32'b11111111110000010000000100010011;
ROM[36396] <= 32'b00000000000000010010001110000011;
ROM[36397] <= 32'b11111111110000010000000100010011;
ROM[36398] <= 32'b00000000000000010010010000000011;
ROM[36399] <= 32'b00000000011101000000001110110011;
ROM[36400] <= 32'b00000000011100010010000000100011;
ROM[36401] <= 32'b00000000010000010000000100010011;
ROM[36402] <= 32'b11111111110000010000000100010011;
ROM[36403] <= 32'b00000000000000010010001110000011;
ROM[36404] <= 32'b00000000110100101000010000110011;
ROM[36405] <= 32'b00000000011101000010011000100011;
ROM[36406] <= 32'b00000000110100101000010000110011;
ROM[36407] <= 32'b00000001100001000010001110000011;
ROM[36408] <= 32'b00000000011100010010000000100011;
ROM[36409] <= 32'b00000000010000010000000100010011;
ROM[36410] <= 32'b00000001111000000000001110010011;
ROM[36411] <= 32'b00000000011100010010000000100011;
ROM[36412] <= 32'b00000000010000010000000100010011;
ROM[36413] <= 32'b11111111110000010000000100010011;
ROM[36414] <= 32'b00000000000000010010001110000011;
ROM[36415] <= 32'b11111111110000010000000100010011;
ROM[36416] <= 32'b00000000000000010010010000000011;
ROM[36417] <= 32'b00000000100000111010001110110011;
ROM[36418] <= 32'b00000000011100010010000000100011;
ROM[36419] <= 32'b00000000010000010000000100010011;
ROM[36420] <= 32'b11111111110000010000000100010011;
ROM[36421] <= 32'b00000000000000010010001110000011;
ROM[36422] <= 32'b00000000000000111000101001100011;
ROM[36423] <= 32'b00000000000000100100001110110111;
ROM[36424] <= 32'b10010011000000111000001110010011;
ROM[36425] <= 32'b00000000111000111000001110110011;
ROM[36426] <= 32'b00000000000000111000000011100111;
ROM[36427] <= 32'b00000100110000000000000011101111;
ROM[36428] <= 32'b00000000110100101000010000110011;
ROM[36429] <= 32'b00000001100001000010001110000011;
ROM[36430] <= 32'b00000000011100010010000000100011;
ROM[36431] <= 32'b00000000010000010000000100010011;
ROM[36432] <= 32'b00000000010100000000001110010011;
ROM[36433] <= 32'b00000000011100010010000000100011;
ROM[36434] <= 32'b00000000010000010000000100010011;
ROM[36435] <= 32'b11111111110000010000000100010011;
ROM[36436] <= 32'b00000000000000010010001110000011;
ROM[36437] <= 32'b11111111110000010000000100010011;
ROM[36438] <= 32'b00000000000000010010010000000011;
ROM[36439] <= 32'b01000000011101000000001110110011;
ROM[36440] <= 32'b00000000011100010010000000100011;
ROM[36441] <= 32'b00000000010000010000000100010011;
ROM[36442] <= 32'b11111111110000010000000100010011;
ROM[36443] <= 32'b00000000000000010010001110000011;
ROM[36444] <= 32'b00000000110100101000010000110011;
ROM[36445] <= 32'b00000000011101000010110000100011;
ROM[36446] <= 32'b00000000000000000000001110010011;
ROM[36447] <= 32'b00000000011100010010000000100011;
ROM[36448] <= 32'b00000000010000010000000100010011;
ROM[36449] <= 32'b00000001010000000000001110010011;
ROM[36450] <= 32'b01000000011100011000001110110011;
ROM[36451] <= 32'b00000000000000111010000010000011;
ROM[36452] <= 32'b11111111110000010000000100010011;
ROM[36453] <= 32'b00000000000000010010001110000011;
ROM[36454] <= 32'b00000000011100100010000000100011;
ROM[36455] <= 32'b00000000010000100000000100010011;
ROM[36456] <= 32'b00000001010000000000001110010011;
ROM[36457] <= 32'b01000000011100011000001110110011;
ROM[36458] <= 32'b00000000010000111010000110000011;
ROM[36459] <= 32'b00000000100000111010001000000011;
ROM[36460] <= 32'b00000000110000111010001010000011;
ROM[36461] <= 32'b00000001000000111010001100000011;
ROM[36462] <= 32'b00000000000000001000000011100111;
ROM[36463] <= 32'b00000000000000100010001110000011;
ROM[36464] <= 32'b00000000011100010010000000100011;
ROM[36465] <= 32'b00000000010000010000000100010011;
ROM[36466] <= 32'b11111111110000010000000100010011;
ROM[36467] <= 32'b00000000000000010010001110000011;
ROM[36468] <= 32'b00000000000000111000001010010011;
ROM[36469] <= 32'b00000000110100101000010000110011;
ROM[36470] <= 32'b00000001010001000010001110000011;
ROM[36471] <= 32'b00000000011100010010000000100011;
ROM[36472] <= 32'b00000000010000010000000100010011;
ROM[36473] <= 32'b00000000000100000000001110010011;
ROM[36474] <= 32'b00000000011100010010000000100011;
ROM[36475] <= 32'b00000000010000010000000100010011;
ROM[36476] <= 32'b11111111110000010000000100010011;
ROM[36477] <= 32'b00000000000000010010001110000011;
ROM[36478] <= 32'b11111111110000010000000100010011;
ROM[36479] <= 32'b00000000000000010010010000000011;
ROM[36480] <= 32'b00000000011101000000001110110011;
ROM[36481] <= 32'b00000000011100010010000000100011;
ROM[36482] <= 32'b00000000010000010000000100010011;
ROM[36483] <= 32'b11111111110000010000000100010011;
ROM[36484] <= 32'b00000000000000010010001110000011;
ROM[36485] <= 32'b00000000110100101000010000110011;
ROM[36486] <= 32'b00000000011101000010101000100011;
ROM[36487] <= 32'b00000000110100101000010000110011;
ROM[36488] <= 32'b00000001010001000010001110000011;
ROM[36489] <= 32'b00000000011100010010000000100011;
ROM[36490] <= 32'b00000000010000010000000100010011;
ROM[36491] <= 32'b00000001010000000000001110010011;
ROM[36492] <= 32'b01000000011100011000001110110011;
ROM[36493] <= 32'b00000000000000111010000010000011;
ROM[36494] <= 32'b11111111110000010000000100010011;
ROM[36495] <= 32'b00000000000000010010001110000011;
ROM[36496] <= 32'b00000000011100100010000000100011;
ROM[36497] <= 32'b00000000010000100000000100010011;
ROM[36498] <= 32'b00000001010000000000001110010011;
ROM[36499] <= 32'b01000000011100011000001110110011;
ROM[36500] <= 32'b00000000010000111010000110000011;
ROM[36501] <= 32'b00000000100000111010001000000011;
ROM[36502] <= 32'b00000000110000111010001010000011;
ROM[36503] <= 32'b00000001000000111010001100000011;
ROM[36504] <= 32'b00000000000000001000000011100111;
ROM[36505] <= 32'b00000000000000100010001110000011;
ROM[36506] <= 32'b00000000011100010010000000100011;
ROM[36507] <= 32'b00000000010000010000000100010011;
ROM[36508] <= 32'b11111111110000010000000100010011;
ROM[36509] <= 32'b00000000000000010010001110000011;
ROM[36510] <= 32'b00000000000000111000001010010011;
ROM[36511] <= 32'b00000000110100101000010000110011;
ROM[36512] <= 32'b00000000010001000010001110000011;
ROM[36513] <= 32'b00000000011100010010000000100011;
ROM[36514] <= 32'b00000000010000010000000100010011;
ROM[36515] <= 32'b00000001010000000000001110010011;
ROM[36516] <= 32'b01000000011100011000001110110011;
ROM[36517] <= 32'b00000000000000111010000010000011;
ROM[36518] <= 32'b11111111110000010000000100010011;
ROM[36519] <= 32'b00000000000000010010001110000011;
ROM[36520] <= 32'b00000000011100100010000000100011;
ROM[36521] <= 32'b00000000010000100000000100010011;
ROM[36522] <= 32'b00000001010000000000001110010011;
ROM[36523] <= 32'b01000000011100011000001110110011;
ROM[36524] <= 32'b00000000010000111010000110000011;
ROM[36525] <= 32'b00000000100000111010001000000011;
ROM[36526] <= 32'b00000000110000111010001010000011;
ROM[36527] <= 32'b00000001000000111010001100000011;
ROM[36528] <= 32'b00000000000000001000000011100111;
ROM[36529] <= 32'b00000000000000100010001110000011;
ROM[36530] <= 32'b00000000011100010010000000100011;
ROM[36531] <= 32'b00000000010000010000000100010011;
ROM[36532] <= 32'b11111111110000010000000100010011;
ROM[36533] <= 32'b00000000000000010010001110000011;
ROM[36534] <= 32'b00000000000000111000001010010011;
ROM[36535] <= 32'b00000000110100101000010000110011;
ROM[36536] <= 32'b00000000000001000010001110000011;
ROM[36537] <= 32'b00000000011100010010000000100011;
ROM[36538] <= 32'b00000000010000010000000100010011;
ROM[36539] <= 32'b00000001010000000000001110010011;
ROM[36540] <= 32'b01000000011100011000001110110011;
ROM[36541] <= 32'b00000000000000111010000010000011;
ROM[36542] <= 32'b11111111110000010000000100010011;
ROM[36543] <= 32'b00000000000000010010001110000011;
ROM[36544] <= 32'b00000000011100100010000000100011;
ROM[36545] <= 32'b00000000010000100000000100010011;
ROM[36546] <= 32'b00000001010000000000001110010011;
ROM[36547] <= 32'b01000000011100011000001110110011;
ROM[36548] <= 32'b00000000010000111010000110000011;
ROM[36549] <= 32'b00000000100000111010001000000011;
ROM[36550] <= 32'b00000000110000111010001010000011;
ROM[36551] <= 32'b00000001000000111010001100000011;
ROM[36552] <= 32'b00000000000000001000000011100111;
ROM[36553] <= 32'b00000000000000100010001110000011;
ROM[36554] <= 32'b00000000011100010010000000100011;
ROM[36555] <= 32'b00000000010000010000000100010011;
ROM[36556] <= 32'b11111111110000010000000100010011;
ROM[36557] <= 32'b00000000000000010010001110000011;
ROM[36558] <= 32'b00000000000000111000001010010011;
ROM[36559] <= 32'b00000000110100101000010000110011;
ROM[36560] <= 32'b00000001010001000010001110000011;
ROM[36561] <= 32'b00000000011100010010000000100011;
ROM[36562] <= 32'b00000000010000010000000100010011;
ROM[36563] <= 32'b00000001010000000000001110010011;
ROM[36564] <= 32'b01000000011100011000001110110011;
ROM[36565] <= 32'b00000000000000111010000010000011;
ROM[36566] <= 32'b11111111110000010000000100010011;
ROM[36567] <= 32'b00000000000000010010001110000011;
ROM[36568] <= 32'b00000000011100100010000000100011;
ROM[36569] <= 32'b00000000010000100000000100010011;
ROM[36570] <= 32'b00000001010000000000001110010011;
ROM[36571] <= 32'b01000000011100011000001110110011;
ROM[36572] <= 32'b00000000010000111010000110000011;
ROM[36573] <= 32'b00000000100000111010001000000011;
ROM[36574] <= 32'b00000000110000111010001010000011;
ROM[36575] <= 32'b00000001000000111010001100000011;
ROM[36576] <= 32'b00000000000000001000000011100111;
ROM[36577] <= 32'b00000000000000100010001110000011;
ROM[36578] <= 32'b00000000011100010010000000100011;
ROM[36579] <= 32'b00000000010000010000000100010011;
ROM[36580] <= 32'b11111111110000010000000100010011;
ROM[36581] <= 32'b00000000000000010010001110000011;
ROM[36582] <= 32'b00000000000000111000001010010011;
ROM[36583] <= 32'b00000000110100101000010000110011;
ROM[36584] <= 32'b00000000100001000010001110000011;
ROM[36585] <= 32'b00000000011100010010000000100011;
ROM[36586] <= 32'b00000000010000010000000100010011;
ROM[36587] <= 32'b00000001010000000000001110010011;
ROM[36588] <= 32'b01000000011100011000001110110011;
ROM[36589] <= 32'b00000000000000111010000010000011;
ROM[36590] <= 32'b11111111110000010000000100010011;
ROM[36591] <= 32'b00000000000000010010001110000011;
ROM[36592] <= 32'b00000000011100100010000000100011;
ROM[36593] <= 32'b00000000010000100000000100010011;
ROM[36594] <= 32'b00000001010000000000001110010011;
ROM[36595] <= 32'b01000000011100011000001110110011;
ROM[36596] <= 32'b00000000010000111010000110000011;
ROM[36597] <= 32'b00000000100000111010001000000011;
ROM[36598] <= 32'b00000000110000111010001010000011;
ROM[36599] <= 32'b00000001000000111010001100000011;
ROM[36600] <= 32'b00000000000000001000000011100111;
ROM[36601] <= 32'b00000000000000100010001110000011;
ROM[36602] <= 32'b00000000011100010010000000100011;
ROM[36603] <= 32'b00000000010000010000000100010011;
ROM[36604] <= 32'b11111111110000010000000100010011;
ROM[36605] <= 32'b00000000000000010010001110000011;
ROM[36606] <= 32'b00000000000000111000001010010011;
ROM[36607] <= 32'b00000000110100101000010000110011;
ROM[36608] <= 32'b00000000110001000010001110000011;
ROM[36609] <= 32'b00000000011100010010000000100011;
ROM[36610] <= 32'b00000000010000010000000100010011;
ROM[36611] <= 32'b00000001010000000000001110010011;
ROM[36612] <= 32'b01000000011100011000001110110011;
ROM[36613] <= 32'b00000000000000111010000010000011;
ROM[36614] <= 32'b11111111110000010000000100010011;
ROM[36615] <= 32'b00000000000000010010001110000011;
ROM[36616] <= 32'b00000000011100100010000000100011;
ROM[36617] <= 32'b00000000010000100000000100010011;
ROM[36618] <= 32'b00000001010000000000001110010011;
ROM[36619] <= 32'b01000000011100011000001110110011;
ROM[36620] <= 32'b00000000010000111010000110000011;
ROM[36621] <= 32'b00000000100000111010001000000011;
ROM[36622] <= 32'b00000000110000111010001010000011;
ROM[36623] <= 32'b00000001000000111010001100000011;
ROM[36624] <= 32'b00000000000000001000000011100111;
ROM[36625] <= 32'b00000000000000100010001110000011;
ROM[36626] <= 32'b00000000011100010010000000100011;
ROM[36627] <= 32'b00000000010000010000000100010011;
ROM[36628] <= 32'b11111111110000010000000100010011;
ROM[36629] <= 32'b00000000000000010010001110000011;
ROM[36630] <= 32'b00000000000000111000001010010011;
ROM[36631] <= 32'b00000000110100101000010000110011;
ROM[36632] <= 32'b00000001000001000010001110000011;
ROM[36633] <= 32'b00000000011100010010000000100011;
ROM[36634] <= 32'b00000000010000010000000100010011;
ROM[36635] <= 32'b00000001010000000000001110010011;
ROM[36636] <= 32'b01000000011100011000001110110011;
ROM[36637] <= 32'b00000000000000111010000010000011;
ROM[36638] <= 32'b11111111110000010000000100010011;
ROM[36639] <= 32'b00000000000000010010001110000011;
ROM[36640] <= 32'b00000000011100100010000000100011;
ROM[36641] <= 32'b00000000010000100000000100010011;
ROM[36642] <= 32'b00000001010000000000001110010011;
ROM[36643] <= 32'b01000000011100011000001110110011;
ROM[36644] <= 32'b00000000010000111010000110000011;
ROM[36645] <= 32'b00000000100000111010001000000011;
ROM[36646] <= 32'b00000000110000111010001010000011;
ROM[36647] <= 32'b00000001000000111010001100000011;
ROM[36648] <= 32'b00000000000000001000000011100111;
ROM[36649] <= 32'b00000000000000010010000000100011;
ROM[36650] <= 32'b00000000010000010000000100010011;
ROM[36651] <= 32'b00000000000000100100001110110111;
ROM[36652] <= 32'b11001111100000111000001110010011;
ROM[36653] <= 32'b00000000111000111000001110110011;
ROM[36654] <= 32'b00000000011100010010000000100011;
ROM[36655] <= 32'b00000000010000010000000100010011;
ROM[36656] <= 32'b00000000001100010010000000100011;
ROM[36657] <= 32'b00000000010000010000000100010011;
ROM[36658] <= 32'b00000000010000010010000000100011;
ROM[36659] <= 32'b00000000010000010000000100010011;
ROM[36660] <= 32'b00000000010100010010000000100011;
ROM[36661] <= 32'b00000000010000010000000100010011;
ROM[36662] <= 32'b00000000011000010010000000100011;
ROM[36663] <= 32'b00000000010000010000000100010011;
ROM[36664] <= 32'b00000001010000000000001110010011;
ROM[36665] <= 32'b00000000000000111000001110010011;
ROM[36666] <= 32'b01000000011100010000001110110011;
ROM[36667] <= 32'b00000000011100000000001000110011;
ROM[36668] <= 32'b00000000001000000000000110110011;
ROM[36669] <= 32'b11000100000111111101000011101111;
ROM[36670] <= 32'b11111111110000010000000100010011;
ROM[36671] <= 32'b00000000000000010010001110000011;
ROM[36672] <= 32'b00000000011100011010000000100011;
ROM[36673] <= 32'b00000000000000011010001110000011;
ROM[36674] <= 32'b00000000011100010010000000100011;
ROM[36675] <= 32'b00000000010000010000000100010011;
ROM[36676] <= 32'b00000000000000100100001110110111;
ROM[36677] <= 32'b11010101110000111000001110010011;
ROM[36678] <= 32'b00000000111000111000001110110011;
ROM[36679] <= 32'b00000000011100010010000000100011;
ROM[36680] <= 32'b00000000010000010000000100010011;
ROM[36681] <= 32'b00000000001100010010000000100011;
ROM[36682] <= 32'b00000000010000010000000100010011;
ROM[36683] <= 32'b00000000010000010010000000100011;
ROM[36684] <= 32'b00000000010000010000000100010011;
ROM[36685] <= 32'b00000000010100010010000000100011;
ROM[36686] <= 32'b00000000010000010000000100010011;
ROM[36687] <= 32'b00000000011000010010000000100011;
ROM[36688] <= 32'b00000000010000010000000100010011;
ROM[36689] <= 32'b00000001010000000000001110010011;
ROM[36690] <= 32'b00000000010000111000001110010011;
ROM[36691] <= 32'b01000000011100010000001110110011;
ROM[36692] <= 32'b00000000011100000000001000110011;
ROM[36693] <= 32'b00000000001000000000000110110011;
ROM[36694] <= 32'b10011100100011111110000011101111;
ROM[36695] <= 32'b11111111110000010000000100010011;
ROM[36696] <= 32'b00000000000000010010001110000011;
ROM[36697] <= 32'b00000000011101100010000000100011;
ROM[36698] <= 32'b00000000000000011010001110000011;
ROM[36699] <= 32'b00000000011100010010000000100011;
ROM[36700] <= 32'b00000000010000010000000100010011;
ROM[36701] <= 32'b00000000000000100100001110110111;
ROM[36702] <= 32'b11011100000000111000001110010011;
ROM[36703] <= 32'b00000000111000111000001110110011;
ROM[36704] <= 32'b00000000011100010010000000100011;
ROM[36705] <= 32'b00000000010000010000000100010011;
ROM[36706] <= 32'b00000000001100010010000000100011;
ROM[36707] <= 32'b00000000010000010000000100010011;
ROM[36708] <= 32'b00000000010000010010000000100011;
ROM[36709] <= 32'b00000000010000010000000100010011;
ROM[36710] <= 32'b00000000010100010010000000100011;
ROM[36711] <= 32'b00000000010000010000000100010011;
ROM[36712] <= 32'b00000000011000010010000000100011;
ROM[36713] <= 32'b00000000010000010000000100010011;
ROM[36714] <= 32'b00000001010000000000001110010011;
ROM[36715] <= 32'b00000000010000111000001110010011;
ROM[36716] <= 32'b01000000011100010000001110110011;
ROM[36717] <= 32'b00000000011100000000001000110011;
ROM[36718] <= 32'b00000000001000000000000110110011;
ROM[36719] <= 32'b11111101100111111101000011101111;
ROM[36720] <= 32'b11111111110000010000000100010011;
ROM[36721] <= 32'b00000000000000010010001110000011;
ROM[36722] <= 32'b00000000011101100010000000100011;
ROM[36723] <= 32'b00000000000000000000001110010011;
ROM[36724] <= 32'b00000000011100010010000000100011;
ROM[36725] <= 32'b00000000010000010000000100010011;
ROM[36726] <= 32'b00000001010000000000001110010011;
ROM[36727] <= 32'b01000000011100011000001110110011;
ROM[36728] <= 32'b00000000000000111010000010000011;
ROM[36729] <= 32'b11111111110000010000000100010011;
ROM[36730] <= 32'b00000000000000010010001110000011;
ROM[36731] <= 32'b00000000011100100010000000100011;
ROM[36732] <= 32'b00000000010000100000000100010011;
ROM[36733] <= 32'b00000001010000000000001110010011;
ROM[36734] <= 32'b01000000011100011000001110110011;
ROM[36735] <= 32'b00000000010000111010000110000011;
ROM[36736] <= 32'b00000000100000111010001000000011;
ROM[36737] <= 32'b00000000110000111010001010000011;
ROM[36738] <= 32'b00000001000000111010001100000011;
ROM[36739] <= 32'b00000000000000001000000011100111;
ROM[36740] <= 32'b00000000100100000000001110010011;
ROM[36741] <= 32'b00000000011100010010000000100011;
ROM[36742] <= 32'b00000000010000010000000100010011;
ROM[36743] <= 32'b00000000000000100100001110110111;
ROM[36744] <= 32'b11100110100000111000001110010011;
ROM[36745] <= 32'b00000000111000111000001110110011;
ROM[36746] <= 32'b00000000011100010010000000100011;
ROM[36747] <= 32'b00000000010000010000000100010011;
ROM[36748] <= 32'b00000000001100010010000000100011;
ROM[36749] <= 32'b00000000010000010000000100010011;
ROM[36750] <= 32'b00000000010000010010000000100011;
ROM[36751] <= 32'b00000000010000010000000100010011;
ROM[36752] <= 32'b00000000010100010010000000100011;
ROM[36753] <= 32'b00000000010000010000000100010011;
ROM[36754] <= 32'b00000000011000010010000000100011;
ROM[36755] <= 32'b00000000010000010000000100010011;
ROM[36756] <= 32'b00000001010000000000001110010011;
ROM[36757] <= 32'b00000000010000111000001110010011;
ROM[36758] <= 32'b01000000011100010000001110110011;
ROM[36759] <= 32'b00000000011100000000001000110011;
ROM[36760] <= 32'b00000000001000000000000110110011;
ROM[36761] <= 32'b10000111000111110000000011101111;
ROM[36762] <= 32'b11111111110000010000000100010011;
ROM[36763] <= 32'b00000000000000010010001110000011;
ROM[36764] <= 32'b00000000000000111000001010010011;
ROM[36765] <= 32'b00000000000000100010001110000011;
ROM[36766] <= 32'b00000000011100010010000000100011;
ROM[36767] <= 32'b00000000010000010000000100010011;
ROM[36768] <= 32'b11111111110000010000000100010011;
ROM[36769] <= 32'b00000000000000010010001110000011;
ROM[36770] <= 32'b00000000110100101000010000110011;
ROM[36771] <= 32'b00000000011101000010000000100011;
ROM[36772] <= 32'b00000000010000100010001110000011;
ROM[36773] <= 32'b00000000011100010010000000100011;
ROM[36774] <= 32'b00000000010000010000000100010011;
ROM[36775] <= 32'b00000000010000000000001110010011;
ROM[36776] <= 32'b00000000011100010010000000100011;
ROM[36777] <= 32'b00000000010000010000000100010011;
ROM[36778] <= 32'b00000000000000100100001110110111;
ROM[36779] <= 32'b11101111010000111000001110010011;
ROM[36780] <= 32'b00000000111000111000001110110011;
ROM[36781] <= 32'b00000000011100010010000000100011;
ROM[36782] <= 32'b00000000010000010000000100010011;
ROM[36783] <= 32'b00000000001100010010000000100011;
ROM[36784] <= 32'b00000000010000010000000100010011;
ROM[36785] <= 32'b00000000010000010010000000100011;
ROM[36786] <= 32'b00000000010000010000000100010011;
ROM[36787] <= 32'b00000000010100010010000000100011;
ROM[36788] <= 32'b00000000010000010000000100010011;
ROM[36789] <= 32'b00000000011000010010000000100011;
ROM[36790] <= 32'b00000000010000010000000100010011;
ROM[36791] <= 32'b00000001010000000000001110010011;
ROM[36792] <= 32'b00000000100000111000001110010011;
ROM[36793] <= 32'b01000000011100010000001110110011;
ROM[36794] <= 32'b00000000011100000000001000110011;
ROM[36795] <= 32'b00000000001000000000000110110011;
ROM[36796] <= 32'b11001011100111101101000011101111;
ROM[36797] <= 32'b11111111110000010000000100010011;
ROM[36798] <= 32'b00000000000000010010001110000011;
ROM[36799] <= 32'b00000000110100101000010000110011;
ROM[36800] <= 32'b00000000011101000010001000100011;
ROM[36801] <= 32'b00000000100000100010001110000011;
ROM[36802] <= 32'b00000000011100010010000000100011;
ROM[36803] <= 32'b00000000010000010000000100010011;
ROM[36804] <= 32'b00000001000000000000001110010011;
ROM[36805] <= 32'b00000000011100010010000000100011;
ROM[36806] <= 32'b00000000010000010000000100010011;
ROM[36807] <= 32'b11111111110000010000000100010011;
ROM[36808] <= 32'b00000000000000010010001110000011;
ROM[36809] <= 32'b11111111110000010000000100010011;
ROM[36810] <= 32'b00000000000000010010010000000011;
ROM[36811] <= 32'b01000000011101000000001110110011;
ROM[36812] <= 32'b00000000011100010010000000100011;
ROM[36813] <= 32'b00000000010000010000000100010011;
ROM[36814] <= 32'b00000000010000000000001110010011;
ROM[36815] <= 32'b00000000011100010010000000100011;
ROM[36816] <= 32'b00000000010000010000000100010011;
ROM[36817] <= 32'b00000000000000100100001110110111;
ROM[36818] <= 32'b11111001000000111000001110010011;
ROM[36819] <= 32'b00000000111000111000001110110011;
ROM[36820] <= 32'b00000000011100010010000000100011;
ROM[36821] <= 32'b00000000010000010000000100010011;
ROM[36822] <= 32'b00000000001100010010000000100011;
ROM[36823] <= 32'b00000000010000010000000100010011;
ROM[36824] <= 32'b00000000010000010010000000100011;
ROM[36825] <= 32'b00000000010000010000000100010011;
ROM[36826] <= 32'b00000000010100010010000000100011;
ROM[36827] <= 32'b00000000010000010000000100010011;
ROM[36828] <= 32'b00000000011000010010000000100011;
ROM[36829] <= 32'b00000000010000010000000100010011;
ROM[36830] <= 32'b00000001010000000000001110010011;
ROM[36831] <= 32'b00000000100000111000001110010011;
ROM[36832] <= 32'b01000000011100010000001110110011;
ROM[36833] <= 32'b00000000011100000000001000110011;
ROM[36834] <= 32'b00000000001000000000000110110011;
ROM[36835] <= 32'b11000001110111101101000011101111;
ROM[36836] <= 32'b11111111110000010000000100010011;
ROM[36837] <= 32'b00000000000000010010001110000011;
ROM[36838] <= 32'b00000000110100101000010000110011;
ROM[36839] <= 32'b00000000011101000010010000100011;
ROM[36840] <= 32'b00000000101000000000001110010011;
ROM[36841] <= 32'b00000000011100010010000000100011;
ROM[36842] <= 32'b00000000010000010000000100010011;
ROM[36843] <= 32'b00000000000000100100001110110111;
ROM[36844] <= 32'b11111111100000111000001110010011;
ROM[36845] <= 32'b00000000111000111000001110110011;
ROM[36846] <= 32'b00000000011100010010000000100011;
ROM[36847] <= 32'b00000000010000010000000100010011;
ROM[36848] <= 32'b00000000001100010010000000100011;
ROM[36849] <= 32'b00000000010000010000000100010011;
ROM[36850] <= 32'b00000000010000010010000000100011;
ROM[36851] <= 32'b00000000010000010000000100010011;
ROM[36852] <= 32'b00000000010100010010000000100011;
ROM[36853] <= 32'b00000000010000010000000100010011;
ROM[36854] <= 32'b00000000011000010010000000100011;
ROM[36855] <= 32'b00000000010000010000000100010011;
ROM[36856] <= 32'b00000001010000000000001110010011;
ROM[36857] <= 32'b00000000010000111000001110010011;
ROM[36858] <= 32'b01000000011100010000001110110011;
ROM[36859] <= 32'b00000000011100000000001000110011;
ROM[36860] <= 32'b00000000001000000000000110110011;
ROM[36861] <= 32'b10001000110011011100000011101111;
ROM[36862] <= 32'b11111111110000010000000100010011;
ROM[36863] <= 32'b00000000000000010010001110000011;
ROM[36864] <= 32'b00000000110100101000010000110011;
ROM[36865] <= 32'b00000000011101000010110000100011;
ROM[36866] <= 32'b00000000101000000000001110010011;
ROM[36867] <= 32'b00000000011100010010000000100011;
ROM[36868] <= 32'b00000000010000010000000100010011;
ROM[36869] <= 32'b00000000000000100100001110110111;
ROM[36870] <= 32'b00000110000000111000001110010011;
ROM[36871] <= 32'b00000000111000111000001110110011;
ROM[36872] <= 32'b00000000011100010010000000100011;
ROM[36873] <= 32'b00000000010000010000000100010011;
ROM[36874] <= 32'b00000000001100010010000000100011;
ROM[36875] <= 32'b00000000010000010000000100010011;
ROM[36876] <= 32'b00000000010000010010000000100011;
ROM[36877] <= 32'b00000000010000010000000100010011;
ROM[36878] <= 32'b00000000010100010010000000100011;
ROM[36879] <= 32'b00000000010000010000000100010011;
ROM[36880] <= 32'b00000000011000010010000000100011;
ROM[36881] <= 32'b00000000010000010000000100010011;
ROM[36882] <= 32'b00000001010000000000001110010011;
ROM[36883] <= 32'b00000000010000111000001110010011;
ROM[36884] <= 32'b01000000011100010000001110110011;
ROM[36885] <= 32'b00000000011100000000001000110011;
ROM[36886] <= 32'b00000000001000000000000110110011;
ROM[36887] <= 32'b10000010010011011100000011101111;
ROM[36888] <= 32'b11111111110000010000000100010011;
ROM[36889] <= 32'b00000000000000010010001110000011;
ROM[36890] <= 32'b00000000110100101000010000110011;
ROM[36891] <= 32'b00000000011101000010111000100011;
ROM[36892] <= 32'b00000011100100000000001110010011;
ROM[36893] <= 32'b00000000011100010010000000100011;
ROM[36894] <= 32'b00000000010000010000000100010011;
ROM[36895] <= 32'b00000000110100101000010000110011;
ROM[36896] <= 32'b00000001110001000010001110000011;
ROM[36897] <= 32'b00000000011100010010000000100011;
ROM[36898] <= 32'b00000000010000010000000100010011;
ROM[36899] <= 32'b00000000000000000000001110010011;
ROM[36900] <= 32'b00000000011100010010000000100011;
ROM[36901] <= 32'b00000000010000010000000100010011;
ROM[36902] <= 32'b00000000010000000000001110010011;
ROM[36903] <= 32'b00000000011100010010000000100011;
ROM[36904] <= 32'b00000000010000010000000100010011;
ROM[36905] <= 32'b00000000000000100100001110110111;
ROM[36906] <= 32'b00001111000000111000001110010011;
ROM[36907] <= 32'b00000000111000111000001110110011;
ROM[36908] <= 32'b00000000011100010010000000100011;
ROM[36909] <= 32'b00000000010000010000000100010011;
ROM[36910] <= 32'b00000000001100010010000000100011;
ROM[36911] <= 32'b00000000010000010000000100010011;
ROM[36912] <= 32'b00000000010000010010000000100011;
ROM[36913] <= 32'b00000000010000010000000100010011;
ROM[36914] <= 32'b00000000010100010010000000100011;
ROM[36915] <= 32'b00000000010000010000000100010011;
ROM[36916] <= 32'b00000000011000010010000000100011;
ROM[36917] <= 32'b00000000010000010000000100010011;
ROM[36918] <= 32'b00000001010000000000001110010011;
ROM[36919] <= 32'b00000000100000111000001110010011;
ROM[36920] <= 32'b01000000011100010000001110110011;
ROM[36921] <= 32'b00000000011100000000001000110011;
ROM[36922] <= 32'b00000000001000000000000110110011;
ROM[36923] <= 32'b11110100000011101101000011101111;
ROM[36924] <= 32'b11111111110000010000000100010011;
ROM[36925] <= 32'b00000000000000010010001110000011;
ROM[36926] <= 32'b11111111110000010000000100010011;
ROM[36927] <= 32'b00000000000000010010010000000011;
ROM[36928] <= 32'b00000000011101000000001110110011;
ROM[36929] <= 32'b00000000011100010010000000100011;
ROM[36930] <= 32'b00000000010000010000000100010011;
ROM[36931] <= 32'b11111111110000010000000100010011;
ROM[36932] <= 32'b00000000000000010010001110000011;
ROM[36933] <= 32'b00000000000000111000001100010011;
ROM[36934] <= 32'b11111111110000010000000100010011;
ROM[36935] <= 32'b00000000000000010010001110000011;
ROM[36936] <= 32'b00000000110100110000010000110011;
ROM[36937] <= 32'b00000000011101000010000000100011;
ROM[36938] <= 32'b00000001100000000000001110010011;
ROM[36939] <= 32'b00000000011100010010000000100011;
ROM[36940] <= 32'b00000000010000010000000100010011;
ROM[36941] <= 32'b00000000110100101000010000110011;
ROM[36942] <= 32'b00000001110001000010001110000011;
ROM[36943] <= 32'b00000000011100010010000000100011;
ROM[36944] <= 32'b00000000010000010000000100010011;
ROM[36945] <= 32'b00000000000100000000001110010011;
ROM[36946] <= 32'b00000000011100010010000000100011;
ROM[36947] <= 32'b00000000010000010000000100010011;
ROM[36948] <= 32'b00000000010000000000001110010011;
ROM[36949] <= 32'b00000000011100010010000000100011;
ROM[36950] <= 32'b00000000010000010000000100010011;
ROM[36951] <= 32'b00000000000000100100001110110111;
ROM[36952] <= 32'b00011010100000111000001110010011;
ROM[36953] <= 32'b00000000111000111000001110110011;
ROM[36954] <= 32'b00000000011100010010000000100011;
ROM[36955] <= 32'b00000000010000010000000100010011;
ROM[36956] <= 32'b00000000001100010010000000100011;
ROM[36957] <= 32'b00000000010000010000000100010011;
ROM[36958] <= 32'b00000000010000010010000000100011;
ROM[36959] <= 32'b00000000010000010000000100010011;
ROM[36960] <= 32'b00000000010100010010000000100011;
ROM[36961] <= 32'b00000000010000010000000100010011;
ROM[36962] <= 32'b00000000011000010010000000100011;
ROM[36963] <= 32'b00000000010000010000000100010011;
ROM[36964] <= 32'b00000001010000000000001110010011;
ROM[36965] <= 32'b00000000100000111000001110010011;
ROM[36966] <= 32'b01000000011100010000001110110011;
ROM[36967] <= 32'b00000000011100000000001000110011;
ROM[36968] <= 32'b00000000001000000000000110110011;
ROM[36969] <= 32'b11101000100011101101000011101111;
ROM[36970] <= 32'b11111111110000010000000100010011;
ROM[36971] <= 32'b00000000000000010010001110000011;
ROM[36972] <= 32'b11111111110000010000000100010011;
ROM[36973] <= 32'b00000000000000010010010000000011;
ROM[36974] <= 32'b00000000011101000000001110110011;
ROM[36975] <= 32'b00000000011100010010000000100011;
ROM[36976] <= 32'b00000000010000010000000100010011;
ROM[36977] <= 32'b11111111110000010000000100010011;
ROM[36978] <= 32'b00000000000000010010001110000011;
ROM[36979] <= 32'b00000000000000111000001100010011;
ROM[36980] <= 32'b11111111110000010000000100010011;
ROM[36981] <= 32'b00000000000000010010001110000011;
ROM[36982] <= 32'b00000000110100110000010000110011;
ROM[36983] <= 32'b00000000011101000010000000100011;
ROM[36984] <= 32'b00000101001100000000001110010011;
ROM[36985] <= 32'b00000000011100010010000000100011;
ROM[36986] <= 32'b00000000010000010000000100010011;
ROM[36987] <= 32'b00000000110100101000010000110011;
ROM[36988] <= 32'b00000001110001000010001110000011;
ROM[36989] <= 32'b00000000011100010010000000100011;
ROM[36990] <= 32'b00000000010000010000000100010011;
ROM[36991] <= 32'b00000000001000000000001110010011;
ROM[36992] <= 32'b00000000011100010010000000100011;
ROM[36993] <= 32'b00000000010000010000000100010011;
ROM[36994] <= 32'b00000000010000000000001110010011;
ROM[36995] <= 32'b00000000011100010010000000100011;
ROM[36996] <= 32'b00000000010000010000000100010011;
ROM[36997] <= 32'b00000000000000100100001110110111;
ROM[36998] <= 32'b00100110000000111000001110010011;
ROM[36999] <= 32'b00000000111000111000001110110011;
ROM[37000] <= 32'b00000000011100010010000000100011;
ROM[37001] <= 32'b00000000010000010000000100010011;
ROM[37002] <= 32'b00000000001100010010000000100011;
ROM[37003] <= 32'b00000000010000010000000100010011;
ROM[37004] <= 32'b00000000010000010010000000100011;
ROM[37005] <= 32'b00000000010000010000000100010011;
ROM[37006] <= 32'b00000000010100010010000000100011;
ROM[37007] <= 32'b00000000010000010000000100010011;
ROM[37008] <= 32'b00000000011000010010000000100011;
ROM[37009] <= 32'b00000000010000010000000100010011;
ROM[37010] <= 32'b00000001010000000000001110010011;
ROM[37011] <= 32'b00000000100000111000001110010011;
ROM[37012] <= 32'b01000000011100010000001110110011;
ROM[37013] <= 32'b00000000011100000000001000110011;
ROM[37014] <= 32'b00000000001000000000000110110011;
ROM[37015] <= 32'b11011101000011101101000011101111;
ROM[37016] <= 32'b11111111110000010000000100010011;
ROM[37017] <= 32'b00000000000000010010001110000011;
ROM[37018] <= 32'b11111111110000010000000100010011;
ROM[37019] <= 32'b00000000000000010010010000000011;
ROM[37020] <= 32'b00000000011101000000001110110011;
ROM[37021] <= 32'b00000000011100010010000000100011;
ROM[37022] <= 32'b00000000010000010000000100010011;
ROM[37023] <= 32'b11111111110000010000000100010011;
ROM[37024] <= 32'b00000000000000010010001110000011;
ROM[37025] <= 32'b00000000000000111000001100010011;
ROM[37026] <= 32'b11111111110000010000000100010011;
ROM[37027] <= 32'b00000000000000010010001110000011;
ROM[37028] <= 32'b00000000110100110000010000110011;
ROM[37029] <= 32'b00000000011101000010000000100011;
ROM[37030] <= 32'b00000100101100000000001110010011;
ROM[37031] <= 32'b00000000011100010010000000100011;
ROM[37032] <= 32'b00000000010000010000000100010011;
ROM[37033] <= 32'b00000000110100101000010000110011;
ROM[37034] <= 32'b00000001110001000010001110000011;
ROM[37035] <= 32'b00000000011100010010000000100011;
ROM[37036] <= 32'b00000000010000010000000100010011;
ROM[37037] <= 32'b00000000001100000000001110010011;
ROM[37038] <= 32'b00000000011100010010000000100011;
ROM[37039] <= 32'b00000000010000010000000100010011;
ROM[37040] <= 32'b00000000010000000000001110010011;
ROM[37041] <= 32'b00000000011100010010000000100011;
ROM[37042] <= 32'b00000000010000010000000100010011;
ROM[37043] <= 32'b00000000000000100100001110110111;
ROM[37044] <= 32'b00110001100000111000001110010011;
ROM[37045] <= 32'b00000000111000111000001110110011;
ROM[37046] <= 32'b00000000011100010010000000100011;
ROM[37047] <= 32'b00000000010000010000000100010011;
ROM[37048] <= 32'b00000000001100010010000000100011;
ROM[37049] <= 32'b00000000010000010000000100010011;
ROM[37050] <= 32'b00000000010000010010000000100011;
ROM[37051] <= 32'b00000000010000010000000100010011;
ROM[37052] <= 32'b00000000010100010010000000100011;
ROM[37053] <= 32'b00000000010000010000000100010011;
ROM[37054] <= 32'b00000000011000010010000000100011;
ROM[37055] <= 32'b00000000010000010000000100010011;
ROM[37056] <= 32'b00000001010000000000001110010011;
ROM[37057] <= 32'b00000000100000111000001110010011;
ROM[37058] <= 32'b01000000011100010000001110110011;
ROM[37059] <= 32'b00000000011100000000001000110011;
ROM[37060] <= 32'b00000000001000000000000110110011;
ROM[37061] <= 32'b11010001100011101101000011101111;
ROM[37062] <= 32'b11111111110000010000000100010011;
ROM[37063] <= 32'b00000000000000010010001110000011;
ROM[37064] <= 32'b11111111110000010000000100010011;
ROM[37065] <= 32'b00000000000000010010010000000011;
ROM[37066] <= 32'b00000000011101000000001110110011;
ROM[37067] <= 32'b00000000011100010010000000100011;
ROM[37068] <= 32'b00000000010000010000000100010011;
ROM[37069] <= 32'b11111111110000010000000100010011;
ROM[37070] <= 32'b00000000000000010010001110000011;
ROM[37071] <= 32'b00000000000000111000001100010011;
ROM[37072] <= 32'b11111111110000010000000100010011;
ROM[37073] <= 32'b00000000000000010010001110000011;
ROM[37074] <= 32'b00000000110100110000010000110011;
ROM[37075] <= 32'b00000000011101000010000000100011;
ROM[37076] <= 32'b00000010010000000000001110010011;
ROM[37077] <= 32'b00000000011100010010000000100011;
ROM[37078] <= 32'b00000000010000010000000100010011;
ROM[37079] <= 32'b00000000110100101000010000110011;
ROM[37080] <= 32'b00000001110001000010001110000011;
ROM[37081] <= 32'b00000000011100010010000000100011;
ROM[37082] <= 32'b00000000010000010000000100010011;
ROM[37083] <= 32'b00000000010000000000001110010011;
ROM[37084] <= 32'b00000000011100010010000000100011;
ROM[37085] <= 32'b00000000010000010000000100010011;
ROM[37086] <= 32'b00000000010000000000001110010011;
ROM[37087] <= 32'b00000000011100010010000000100011;
ROM[37088] <= 32'b00000000010000010000000100010011;
ROM[37089] <= 32'b00000000000000100100001110110111;
ROM[37090] <= 32'b00111101000000111000001110010011;
ROM[37091] <= 32'b00000000111000111000001110110011;
ROM[37092] <= 32'b00000000011100010010000000100011;
ROM[37093] <= 32'b00000000010000010000000100010011;
ROM[37094] <= 32'b00000000001100010010000000100011;
ROM[37095] <= 32'b00000000010000010000000100010011;
ROM[37096] <= 32'b00000000010000010010000000100011;
ROM[37097] <= 32'b00000000010000010000000100010011;
ROM[37098] <= 32'b00000000010100010010000000100011;
ROM[37099] <= 32'b00000000010000010000000100010011;
ROM[37100] <= 32'b00000000011000010010000000100011;
ROM[37101] <= 32'b00000000010000010000000100010011;
ROM[37102] <= 32'b00000001010000000000001110010011;
ROM[37103] <= 32'b00000000100000111000001110010011;
ROM[37104] <= 32'b01000000011100010000001110110011;
ROM[37105] <= 32'b00000000011100000000001000110011;
ROM[37106] <= 32'b00000000001000000000000110110011;
ROM[37107] <= 32'b11000110000011101101000011101111;
ROM[37108] <= 32'b11111111110000010000000100010011;
ROM[37109] <= 32'b00000000000000010010001110000011;
ROM[37110] <= 32'b11111111110000010000000100010011;
ROM[37111] <= 32'b00000000000000010010010000000011;
ROM[37112] <= 32'b00000000011101000000001110110011;
ROM[37113] <= 32'b00000000011100010010000000100011;
ROM[37114] <= 32'b00000000010000010000000100010011;
ROM[37115] <= 32'b11111111110000010000000100010011;
ROM[37116] <= 32'b00000000000000010010001110000011;
ROM[37117] <= 32'b00000000000000111000001100010011;
ROM[37118] <= 32'b11111111110000010000000100010011;
ROM[37119] <= 32'b00000000000000010010001110000011;
ROM[37120] <= 32'b00000000110100110000010000110011;
ROM[37121] <= 32'b00000000011101000010000000100011;
ROM[37122] <= 32'b00000110001100000000001110010011;
ROM[37123] <= 32'b00000000011100010010000000100011;
ROM[37124] <= 32'b00000000010000010000000100010011;
ROM[37125] <= 32'b00000000110100101000010000110011;
ROM[37126] <= 32'b00000001110001000010001110000011;
ROM[37127] <= 32'b00000000011100010010000000100011;
ROM[37128] <= 32'b00000000010000010000000100010011;
ROM[37129] <= 32'b00000000010100000000001110010011;
ROM[37130] <= 32'b00000000011100010010000000100011;
ROM[37131] <= 32'b00000000010000010000000100010011;
ROM[37132] <= 32'b00000000010000000000001110010011;
ROM[37133] <= 32'b00000000011100010010000000100011;
ROM[37134] <= 32'b00000000010000010000000100010011;
ROM[37135] <= 32'b00000000000000100100001110110111;
ROM[37136] <= 32'b01001000100000111000001110010011;
ROM[37137] <= 32'b00000000111000111000001110110011;
ROM[37138] <= 32'b00000000011100010010000000100011;
ROM[37139] <= 32'b00000000010000010000000100010011;
ROM[37140] <= 32'b00000000001100010010000000100011;
ROM[37141] <= 32'b00000000010000010000000100010011;
ROM[37142] <= 32'b00000000010000010010000000100011;
ROM[37143] <= 32'b00000000010000010000000100010011;
ROM[37144] <= 32'b00000000010100010010000000100011;
ROM[37145] <= 32'b00000000010000010000000100010011;
ROM[37146] <= 32'b00000000011000010010000000100011;
ROM[37147] <= 32'b00000000010000010000000100010011;
ROM[37148] <= 32'b00000001010000000000001110010011;
ROM[37149] <= 32'b00000000100000111000001110010011;
ROM[37150] <= 32'b01000000011100010000001110110011;
ROM[37151] <= 32'b00000000011100000000001000110011;
ROM[37152] <= 32'b00000000001000000000000110110011;
ROM[37153] <= 32'b10111010100011101101000011101111;
ROM[37154] <= 32'b11111111110000010000000100010011;
ROM[37155] <= 32'b00000000000000010010001110000011;
ROM[37156] <= 32'b11111111110000010000000100010011;
ROM[37157] <= 32'b00000000000000010010010000000011;
ROM[37158] <= 32'b00000000011101000000001110110011;
ROM[37159] <= 32'b00000000011100010010000000100011;
ROM[37160] <= 32'b00000000010000010000000100010011;
ROM[37161] <= 32'b11111111110000010000000100010011;
ROM[37162] <= 32'b00000000000000010010001110000011;
ROM[37163] <= 32'b00000000000000111000001100010011;
ROM[37164] <= 32'b11111111110000010000000100010011;
ROM[37165] <= 32'b00000000000000010010001110000011;
ROM[37166] <= 32'b00000000110100110000010000110011;
ROM[37167] <= 32'b00000000011101000010000000100011;
ROM[37168] <= 32'b00000100010000000000001110010011;
ROM[37169] <= 32'b00000000011100010010000000100011;
ROM[37170] <= 32'b00000000010000010000000100010011;
ROM[37171] <= 32'b00000000110100101000010000110011;
ROM[37172] <= 32'b00000001110001000010001110000011;
ROM[37173] <= 32'b00000000011100010010000000100011;
ROM[37174] <= 32'b00000000010000010000000100010011;
ROM[37175] <= 32'b00000000011000000000001110010011;
ROM[37176] <= 32'b00000000011100010010000000100011;
ROM[37177] <= 32'b00000000010000010000000100010011;
ROM[37178] <= 32'b00000000010000000000001110010011;
ROM[37179] <= 32'b00000000011100010010000000100011;
ROM[37180] <= 32'b00000000010000010000000100010011;
ROM[37181] <= 32'b00000000000000100100001110110111;
ROM[37182] <= 32'b01010100000000111000001110010011;
ROM[37183] <= 32'b00000000111000111000001110110011;
ROM[37184] <= 32'b00000000011100010010000000100011;
ROM[37185] <= 32'b00000000010000010000000100010011;
ROM[37186] <= 32'b00000000001100010010000000100011;
ROM[37187] <= 32'b00000000010000010000000100010011;
ROM[37188] <= 32'b00000000010000010010000000100011;
ROM[37189] <= 32'b00000000010000010000000100010011;
ROM[37190] <= 32'b00000000010100010010000000100011;
ROM[37191] <= 32'b00000000010000010000000100010011;
ROM[37192] <= 32'b00000000011000010010000000100011;
ROM[37193] <= 32'b00000000010000010000000100010011;
ROM[37194] <= 32'b00000001010000000000001110010011;
ROM[37195] <= 32'b00000000100000111000001110010011;
ROM[37196] <= 32'b01000000011100010000001110110011;
ROM[37197] <= 32'b00000000011100000000001000110011;
ROM[37198] <= 32'b00000000001000000000000110110011;
ROM[37199] <= 32'b10101111000011101101000011101111;
ROM[37200] <= 32'b11111111110000010000000100010011;
ROM[37201] <= 32'b00000000000000010010001110000011;
ROM[37202] <= 32'b11111111110000010000000100010011;
ROM[37203] <= 32'b00000000000000010010010000000011;
ROM[37204] <= 32'b00000000011101000000001110110011;
ROM[37205] <= 32'b00000000011100010010000000100011;
ROM[37206] <= 32'b00000000010000010000000100010011;
ROM[37207] <= 32'b11111111110000010000000100010011;
ROM[37208] <= 32'b00000000000000010010001110000011;
ROM[37209] <= 32'b00000000000000111000001100010011;
ROM[37210] <= 32'b11111111110000010000000100010011;
ROM[37211] <= 32'b00000000000000010010001110000011;
ROM[37212] <= 32'b00000000110100110000010000110011;
ROM[37213] <= 32'b00000000011101000010000000100011;
ROM[37214] <= 32'b00000010101000000000001110010011;
ROM[37215] <= 32'b00000000011100010010000000100011;
ROM[37216] <= 32'b00000000010000010000000100010011;
ROM[37217] <= 32'b00000000110100101000010000110011;
ROM[37218] <= 32'b00000001110001000010001110000011;
ROM[37219] <= 32'b00000000011100010010000000100011;
ROM[37220] <= 32'b00000000010000010000000100010011;
ROM[37221] <= 32'b00000000011100000000001110010011;
ROM[37222] <= 32'b00000000011100010010000000100011;
ROM[37223] <= 32'b00000000010000010000000100010011;
ROM[37224] <= 32'b00000000010000000000001110010011;
ROM[37225] <= 32'b00000000011100010010000000100011;
ROM[37226] <= 32'b00000000010000010000000100010011;
ROM[37227] <= 32'b00000000000000100100001110110111;
ROM[37228] <= 32'b01011111100000111000001110010011;
ROM[37229] <= 32'b00000000111000111000001110110011;
ROM[37230] <= 32'b00000000011100010010000000100011;
ROM[37231] <= 32'b00000000010000010000000100010011;
ROM[37232] <= 32'b00000000001100010010000000100011;
ROM[37233] <= 32'b00000000010000010000000100010011;
ROM[37234] <= 32'b00000000010000010010000000100011;
ROM[37235] <= 32'b00000000010000010000000100010011;
ROM[37236] <= 32'b00000000010100010010000000100011;
ROM[37237] <= 32'b00000000010000010000000100010011;
ROM[37238] <= 32'b00000000011000010010000000100011;
ROM[37239] <= 32'b00000000010000010000000100010011;
ROM[37240] <= 32'b00000001010000000000001110010011;
ROM[37241] <= 32'b00000000100000111000001110010011;
ROM[37242] <= 32'b01000000011100010000001110110011;
ROM[37243] <= 32'b00000000011100000000001000110011;
ROM[37244] <= 32'b00000000001000000000000110110011;
ROM[37245] <= 32'b10100011100011101101000011101111;
ROM[37246] <= 32'b11111111110000010000000100010011;
ROM[37247] <= 32'b00000000000000010010001110000011;
ROM[37248] <= 32'b11111111110000010000000100010011;
ROM[37249] <= 32'b00000000000000010010010000000011;
ROM[37250] <= 32'b00000000011101000000001110110011;
ROM[37251] <= 32'b00000000011100010010000000100011;
ROM[37252] <= 32'b00000000010000010000000100010011;
ROM[37253] <= 32'b11111111110000010000000100010011;
ROM[37254] <= 32'b00000000000000010010001110000011;
ROM[37255] <= 32'b00000000000000111000001100010011;
ROM[37256] <= 32'b11111111110000010000000100010011;
ROM[37257] <= 32'b00000000000000010010001110000011;
ROM[37258] <= 32'b00000000110100110000010000110011;
ROM[37259] <= 32'b00000000011101000010000000100011;
ROM[37260] <= 32'b00000101101000000000001110010011;
ROM[37261] <= 32'b00000000011100010010000000100011;
ROM[37262] <= 32'b00000000010000010000000100010011;
ROM[37263] <= 32'b00000000110100101000010000110011;
ROM[37264] <= 32'b00000001110001000010001110000011;
ROM[37265] <= 32'b00000000011100010010000000100011;
ROM[37266] <= 32'b00000000010000010000000100010011;
ROM[37267] <= 32'b00000000100000000000001110010011;
ROM[37268] <= 32'b00000000011100010010000000100011;
ROM[37269] <= 32'b00000000010000010000000100010011;
ROM[37270] <= 32'b00000000010000000000001110010011;
ROM[37271] <= 32'b00000000011100010010000000100011;
ROM[37272] <= 32'b00000000010000010000000100010011;
ROM[37273] <= 32'b00000000000000100100001110110111;
ROM[37274] <= 32'b01101011000000111000001110010011;
ROM[37275] <= 32'b00000000111000111000001110110011;
ROM[37276] <= 32'b00000000011100010010000000100011;
ROM[37277] <= 32'b00000000010000010000000100010011;
ROM[37278] <= 32'b00000000001100010010000000100011;
ROM[37279] <= 32'b00000000010000010000000100010011;
ROM[37280] <= 32'b00000000010000010010000000100011;
ROM[37281] <= 32'b00000000010000010000000100010011;
ROM[37282] <= 32'b00000000010100010010000000100011;
ROM[37283] <= 32'b00000000010000010000000100010011;
ROM[37284] <= 32'b00000000011000010010000000100011;
ROM[37285] <= 32'b00000000010000010000000100010011;
ROM[37286] <= 32'b00000001010000000000001110010011;
ROM[37287] <= 32'b00000000100000111000001110010011;
ROM[37288] <= 32'b01000000011100010000001110110011;
ROM[37289] <= 32'b00000000011100000000001000110011;
ROM[37290] <= 32'b00000000001000000000000110110011;
ROM[37291] <= 32'b10011000000011101101000011101111;
ROM[37292] <= 32'b11111111110000010000000100010011;
ROM[37293] <= 32'b00000000000000010010001110000011;
ROM[37294] <= 32'b11111111110000010000000100010011;
ROM[37295] <= 32'b00000000000000010010010000000011;
ROM[37296] <= 32'b00000000011101000000001110110011;
ROM[37297] <= 32'b00000000011100010010000000100011;
ROM[37298] <= 32'b00000000010000010000000100010011;
ROM[37299] <= 32'b11111111110000010000000100010011;
ROM[37300] <= 32'b00000000000000010010001110000011;
ROM[37301] <= 32'b00000000000000111000001100010011;
ROM[37302] <= 32'b11111111110000010000000100010011;
ROM[37303] <= 32'b00000000000000010010001110000011;
ROM[37304] <= 32'b00000000110100110000010000110011;
ROM[37305] <= 32'b00000000011101000010000000100011;
ROM[37306] <= 32'b00000100100000000000001110010011;
ROM[37307] <= 32'b00000000011100010010000000100011;
ROM[37308] <= 32'b00000000010000010000000100010011;
ROM[37309] <= 32'b00000000110100101000010000110011;
ROM[37310] <= 32'b00000001110001000010001110000011;
ROM[37311] <= 32'b00000000011100010010000000100011;
ROM[37312] <= 32'b00000000010000010000000100010011;
ROM[37313] <= 32'b00000000100100000000001110010011;
ROM[37314] <= 32'b00000000011100010010000000100011;
ROM[37315] <= 32'b00000000010000010000000100010011;
ROM[37316] <= 32'b00000000010000000000001110010011;
ROM[37317] <= 32'b00000000011100010010000000100011;
ROM[37318] <= 32'b00000000010000010000000100010011;
ROM[37319] <= 32'b00000000000000100100001110110111;
ROM[37320] <= 32'b01110110100000111000001110010011;
ROM[37321] <= 32'b00000000111000111000001110110011;
ROM[37322] <= 32'b00000000011100010010000000100011;
ROM[37323] <= 32'b00000000010000010000000100010011;
ROM[37324] <= 32'b00000000001100010010000000100011;
ROM[37325] <= 32'b00000000010000010000000100010011;
ROM[37326] <= 32'b00000000010000010010000000100011;
ROM[37327] <= 32'b00000000010000010000000100010011;
ROM[37328] <= 32'b00000000010100010010000000100011;
ROM[37329] <= 32'b00000000010000010000000100010011;
ROM[37330] <= 32'b00000000011000010010000000100011;
ROM[37331] <= 32'b00000000010000010000000100010011;
ROM[37332] <= 32'b00000001010000000000001110010011;
ROM[37333] <= 32'b00000000100000111000001110010011;
ROM[37334] <= 32'b01000000011100010000001110110011;
ROM[37335] <= 32'b00000000011100000000001000110011;
ROM[37336] <= 32'b00000000001000000000000110110011;
ROM[37337] <= 32'b10001100100011101101000011101111;
ROM[37338] <= 32'b11111111110000010000000100010011;
ROM[37339] <= 32'b00000000000000010010001110000011;
ROM[37340] <= 32'b11111111110000010000000100010011;
ROM[37341] <= 32'b00000000000000010010010000000011;
ROM[37342] <= 32'b00000000011101000000001110110011;
ROM[37343] <= 32'b00000000011100010010000000100011;
ROM[37344] <= 32'b00000000010000010000000100010011;
ROM[37345] <= 32'b11111111110000010000000100010011;
ROM[37346] <= 32'b00000000000000010010001110000011;
ROM[37347] <= 32'b00000000000000111000001100010011;
ROM[37348] <= 32'b11111111110000010000000100010011;
ROM[37349] <= 32'b00000000000000010010001110000011;
ROM[37350] <= 32'b00000000110100110000010000110011;
ROM[37351] <= 32'b00000000011101000010000000100011;
ROM[37352] <= 32'b00000011011000000000001110010011;
ROM[37353] <= 32'b00000000011100010010000000100011;
ROM[37354] <= 32'b00000000010000010000000100010011;
ROM[37355] <= 32'b00000000110100101000010000110011;
ROM[37356] <= 32'b00000001100001000010001110000011;
ROM[37357] <= 32'b00000000011100010010000000100011;
ROM[37358] <= 32'b00000000010000010000000100010011;
ROM[37359] <= 32'b00000000000000000000001110010011;
ROM[37360] <= 32'b00000000011100010010000000100011;
ROM[37361] <= 32'b00000000010000010000000100010011;
ROM[37362] <= 32'b00000000010000000000001110010011;
ROM[37363] <= 32'b00000000011100010010000000100011;
ROM[37364] <= 32'b00000000010000010000000100010011;
ROM[37365] <= 32'b00000000000000100101001110110111;
ROM[37366] <= 32'b10000010000000111000001110010011;
ROM[37367] <= 32'b00000000111000111000001110110011;
ROM[37368] <= 32'b00000000011100010010000000100011;
ROM[37369] <= 32'b00000000010000010000000100010011;
ROM[37370] <= 32'b00000000001100010010000000100011;
ROM[37371] <= 32'b00000000010000010000000100010011;
ROM[37372] <= 32'b00000000010000010010000000100011;
ROM[37373] <= 32'b00000000010000010000000100010011;
ROM[37374] <= 32'b00000000010100010010000000100011;
ROM[37375] <= 32'b00000000010000010000000100010011;
ROM[37376] <= 32'b00000000011000010010000000100011;
ROM[37377] <= 32'b00000000010000010000000100010011;
ROM[37378] <= 32'b00000001010000000000001110010011;
ROM[37379] <= 32'b00000000100000111000001110010011;
ROM[37380] <= 32'b01000000011100010000001110110011;
ROM[37381] <= 32'b00000000011100000000001000110011;
ROM[37382] <= 32'b00000000001000000000000110110011;
ROM[37383] <= 32'b10000001000011101101000011101111;
ROM[37384] <= 32'b11111111110000010000000100010011;
ROM[37385] <= 32'b00000000000000010010001110000011;
ROM[37386] <= 32'b11111111110000010000000100010011;
ROM[37387] <= 32'b00000000000000010010010000000011;
ROM[37388] <= 32'b00000000011101000000001110110011;
ROM[37389] <= 32'b00000000011100010010000000100011;
ROM[37390] <= 32'b00000000010000010000000100010011;
ROM[37391] <= 32'b11111111110000010000000100010011;
ROM[37392] <= 32'b00000000000000010010001110000011;
ROM[37393] <= 32'b00000000000000111000001100010011;
ROM[37394] <= 32'b11111111110000010000000100010011;
ROM[37395] <= 32'b00000000000000010010001110000011;
ROM[37396] <= 32'b00000000110100110000010000110011;
ROM[37397] <= 32'b00000000011101000010000000100011;
ROM[37398] <= 32'b00000010101100000000001110010011;
ROM[37399] <= 32'b00000000011100010010000000100011;
ROM[37400] <= 32'b00000000010000010000000100010011;
ROM[37401] <= 32'b00000000110100101000010000110011;
ROM[37402] <= 32'b00000001100001000010001110000011;
ROM[37403] <= 32'b00000000011100010010000000100011;
ROM[37404] <= 32'b00000000010000010000000100010011;
ROM[37405] <= 32'b00000000000100000000001110010011;
ROM[37406] <= 32'b00000000011100010010000000100011;
ROM[37407] <= 32'b00000000010000010000000100010011;
ROM[37408] <= 32'b00000000010000000000001110010011;
ROM[37409] <= 32'b00000000011100010010000000100011;
ROM[37410] <= 32'b00000000010000010000000100010011;
ROM[37411] <= 32'b00000000000000100101001110110111;
ROM[37412] <= 32'b10001101100000111000001110010011;
ROM[37413] <= 32'b00000000111000111000001110110011;
ROM[37414] <= 32'b00000000011100010010000000100011;
ROM[37415] <= 32'b00000000010000010000000100010011;
ROM[37416] <= 32'b00000000001100010010000000100011;
ROM[37417] <= 32'b00000000010000010000000100010011;
ROM[37418] <= 32'b00000000010000010010000000100011;
ROM[37419] <= 32'b00000000010000010000000100010011;
ROM[37420] <= 32'b00000000010100010010000000100011;
ROM[37421] <= 32'b00000000010000010000000100010011;
ROM[37422] <= 32'b00000000011000010010000000100011;
ROM[37423] <= 32'b00000000010000010000000100010011;
ROM[37424] <= 32'b00000001010000000000001110010011;
ROM[37425] <= 32'b00000000100000111000001110010011;
ROM[37426] <= 32'b01000000011100010000001110110011;
ROM[37427] <= 32'b00000000011100000000001000110011;
ROM[37428] <= 32'b00000000001000000000000110110011;
ROM[37429] <= 32'b11110101100111101100000011101111;
ROM[37430] <= 32'b11111111110000010000000100010011;
ROM[37431] <= 32'b00000000000000010010001110000011;
ROM[37432] <= 32'b11111111110000010000000100010011;
ROM[37433] <= 32'b00000000000000010010010000000011;
ROM[37434] <= 32'b00000000011101000000001110110011;
ROM[37435] <= 32'b00000000011100010010000000100011;
ROM[37436] <= 32'b00000000010000010000000100010011;
ROM[37437] <= 32'b11111111110000010000000100010011;
ROM[37438] <= 32'b00000000000000010010001110000011;
ROM[37439] <= 32'b00000000000000111000001100010011;
ROM[37440] <= 32'b11111111110000010000000100010011;
ROM[37441] <= 32'b00000000000000010010001110000011;
ROM[37442] <= 32'b00000000110100110000010000110011;
ROM[37443] <= 32'b00000000011101000010000000100011;
ROM[37444] <= 32'b00000101100000000000001110010011;
ROM[37445] <= 32'b00000000011100010010000000100011;
ROM[37446] <= 32'b00000000010000010000000100010011;
ROM[37447] <= 32'b00000000110100101000010000110011;
ROM[37448] <= 32'b00000001100001000010001110000011;
ROM[37449] <= 32'b00000000011100010010000000100011;
ROM[37450] <= 32'b00000000010000010000000100010011;
ROM[37451] <= 32'b00000000001000000000001110010011;
ROM[37452] <= 32'b00000000011100010010000000100011;
ROM[37453] <= 32'b00000000010000010000000100010011;
ROM[37454] <= 32'b00000000010000000000001110010011;
ROM[37455] <= 32'b00000000011100010010000000100011;
ROM[37456] <= 32'b00000000010000010000000100010011;
ROM[37457] <= 32'b00000000000000100101001110110111;
ROM[37458] <= 32'b10011001000000111000001110010011;
ROM[37459] <= 32'b00000000111000111000001110110011;
ROM[37460] <= 32'b00000000011100010010000000100011;
ROM[37461] <= 32'b00000000010000010000000100010011;
ROM[37462] <= 32'b00000000001100010010000000100011;
ROM[37463] <= 32'b00000000010000010000000100010011;
ROM[37464] <= 32'b00000000010000010010000000100011;
ROM[37465] <= 32'b00000000010000010000000100010011;
ROM[37466] <= 32'b00000000010100010010000000100011;
ROM[37467] <= 32'b00000000010000010000000100010011;
ROM[37468] <= 32'b00000000011000010010000000100011;
ROM[37469] <= 32'b00000000010000010000000100010011;
ROM[37470] <= 32'b00000001010000000000001110010011;
ROM[37471] <= 32'b00000000100000111000001110010011;
ROM[37472] <= 32'b01000000011100010000001110110011;
ROM[37473] <= 32'b00000000011100000000001000110011;
ROM[37474] <= 32'b00000000001000000000000110110011;
ROM[37475] <= 32'b11101010000111101100000011101111;
ROM[37476] <= 32'b11111111110000010000000100010011;
ROM[37477] <= 32'b00000000000000010010001110000011;
ROM[37478] <= 32'b11111111110000010000000100010011;
ROM[37479] <= 32'b00000000000000010010010000000011;
ROM[37480] <= 32'b00000000011101000000001110110011;
ROM[37481] <= 32'b00000000011100010010000000100011;
ROM[37482] <= 32'b00000000010000010000000100010011;
ROM[37483] <= 32'b11111111110000010000000100010011;
ROM[37484] <= 32'b00000000000000010010001110000011;
ROM[37485] <= 32'b00000000000000111000001100010011;
ROM[37486] <= 32'b11111111110000010000000100010011;
ROM[37487] <= 32'b00000000000000010010001110000011;
ROM[37488] <= 32'b00000000110100110000010000110011;
ROM[37489] <= 32'b00000000011101000010000000100011;
ROM[37490] <= 32'b00000100101100000000001110010011;
ROM[37491] <= 32'b00000000011100010010000000100011;
ROM[37492] <= 32'b00000000010000010000000100010011;
ROM[37493] <= 32'b00000000110100101000010000110011;
ROM[37494] <= 32'b00000001100001000010001110000011;
ROM[37495] <= 32'b00000000011100010010000000100011;
ROM[37496] <= 32'b00000000010000010000000100010011;
ROM[37497] <= 32'b00000000001100000000001110010011;
ROM[37498] <= 32'b00000000011100010010000000100011;
ROM[37499] <= 32'b00000000010000010000000100010011;
ROM[37500] <= 32'b00000000010000000000001110010011;
ROM[37501] <= 32'b00000000011100010010000000100011;
ROM[37502] <= 32'b00000000010000010000000100010011;
ROM[37503] <= 32'b00000000000000100101001110110111;
ROM[37504] <= 32'b10100100100000111000001110010011;
ROM[37505] <= 32'b00000000111000111000001110110011;
ROM[37506] <= 32'b00000000011100010010000000100011;
ROM[37507] <= 32'b00000000010000010000000100010011;
ROM[37508] <= 32'b00000000001100010010000000100011;
ROM[37509] <= 32'b00000000010000010000000100010011;
ROM[37510] <= 32'b00000000010000010010000000100011;
ROM[37511] <= 32'b00000000010000010000000100010011;
ROM[37512] <= 32'b00000000010100010010000000100011;
ROM[37513] <= 32'b00000000010000010000000100010011;
ROM[37514] <= 32'b00000000011000010010000000100011;
ROM[37515] <= 32'b00000000010000010000000100010011;
ROM[37516] <= 32'b00000001010000000000001110010011;
ROM[37517] <= 32'b00000000100000111000001110010011;
ROM[37518] <= 32'b01000000011100010000001110110011;
ROM[37519] <= 32'b00000000011100000000001000110011;
ROM[37520] <= 32'b00000000001000000000000110110011;
ROM[37521] <= 32'b11011110100111101100000011101111;
ROM[37522] <= 32'b11111111110000010000000100010011;
ROM[37523] <= 32'b00000000000000010010001110000011;
ROM[37524] <= 32'b11111111110000010000000100010011;
ROM[37525] <= 32'b00000000000000010010010000000011;
ROM[37526] <= 32'b00000000011101000000001110110011;
ROM[37527] <= 32'b00000000011100010010000000100011;
ROM[37528] <= 32'b00000000010000010000000100010011;
ROM[37529] <= 32'b11111111110000010000000100010011;
ROM[37530] <= 32'b00000000000000010010001110000011;
ROM[37531] <= 32'b00000000000000111000001100010011;
ROM[37532] <= 32'b11111111110000010000000100010011;
ROM[37533] <= 32'b00000000000000010010001110000011;
ROM[37534] <= 32'b00000000110100110000010000110011;
ROM[37535] <= 32'b00000000011101000010000000100011;
ROM[37536] <= 32'b00000101011100000000001110010011;
ROM[37537] <= 32'b00000000011100010010000000100011;
ROM[37538] <= 32'b00000000010000010000000100010011;
ROM[37539] <= 32'b00000000110100101000010000110011;
ROM[37540] <= 32'b00000001100001000010001110000011;
ROM[37541] <= 32'b00000000011100010010000000100011;
ROM[37542] <= 32'b00000000010000010000000100010011;
ROM[37543] <= 32'b00000000010000000000001110010011;
ROM[37544] <= 32'b00000000011100010010000000100011;
ROM[37545] <= 32'b00000000010000010000000100010011;
ROM[37546] <= 32'b00000000010000000000001110010011;
ROM[37547] <= 32'b00000000011100010010000000100011;
ROM[37548] <= 32'b00000000010000010000000100010011;
ROM[37549] <= 32'b00000000000000100101001110110111;
ROM[37550] <= 32'b10110000000000111000001110010011;
ROM[37551] <= 32'b00000000111000111000001110110011;
ROM[37552] <= 32'b00000000011100010010000000100011;
ROM[37553] <= 32'b00000000010000010000000100010011;
ROM[37554] <= 32'b00000000001100010010000000100011;
ROM[37555] <= 32'b00000000010000010000000100010011;
ROM[37556] <= 32'b00000000010000010010000000100011;
ROM[37557] <= 32'b00000000010000010000000100010011;
ROM[37558] <= 32'b00000000010100010010000000100011;
ROM[37559] <= 32'b00000000010000010000000100010011;
ROM[37560] <= 32'b00000000011000010010000000100011;
ROM[37561] <= 32'b00000000010000010000000100010011;
ROM[37562] <= 32'b00000001010000000000001110010011;
ROM[37563] <= 32'b00000000100000111000001110010011;
ROM[37564] <= 32'b01000000011100010000001110110011;
ROM[37565] <= 32'b00000000011100000000001000110011;
ROM[37566] <= 32'b00000000001000000000000110110011;
ROM[37567] <= 32'b11010011000111101100000011101111;
ROM[37568] <= 32'b11111111110000010000000100010011;
ROM[37569] <= 32'b00000000000000010010001110000011;
ROM[37570] <= 32'b11111111110000010000000100010011;
ROM[37571] <= 32'b00000000000000010010010000000011;
ROM[37572] <= 32'b00000000011101000000001110110011;
ROM[37573] <= 32'b00000000011100010010000000100011;
ROM[37574] <= 32'b00000000010000010000000100010011;
ROM[37575] <= 32'b11111111110000010000000100010011;
ROM[37576] <= 32'b00000000000000010010001110000011;
ROM[37577] <= 32'b00000000000000111000001100010011;
ROM[37578] <= 32'b11111111110000010000000100010011;
ROM[37579] <= 32'b00000000000000010010001110000011;
ROM[37580] <= 32'b00000000110100110000010000110011;
ROM[37581] <= 32'b00000000011101000010000000100011;
ROM[37582] <= 32'b00000001010100000000001110010011;
ROM[37583] <= 32'b00000000011100010010000000100011;
ROM[37584] <= 32'b00000000010000010000000100010011;
ROM[37585] <= 32'b00000000110100101000010000110011;
ROM[37586] <= 32'b00000001100001000010001110000011;
ROM[37587] <= 32'b00000000011100010010000000100011;
ROM[37588] <= 32'b00000000010000010000000100010011;
ROM[37589] <= 32'b00000000010100000000001110010011;
ROM[37590] <= 32'b00000000011100010010000000100011;
ROM[37591] <= 32'b00000000010000010000000100010011;
ROM[37592] <= 32'b00000000010000000000001110010011;
ROM[37593] <= 32'b00000000011100010010000000100011;
ROM[37594] <= 32'b00000000010000010000000100010011;
ROM[37595] <= 32'b00000000000000100101001110110111;
ROM[37596] <= 32'b10111011100000111000001110010011;
ROM[37597] <= 32'b00000000111000111000001110110011;
ROM[37598] <= 32'b00000000011100010010000000100011;
ROM[37599] <= 32'b00000000010000010000000100010011;
ROM[37600] <= 32'b00000000001100010010000000100011;
ROM[37601] <= 32'b00000000010000010000000100010011;
ROM[37602] <= 32'b00000000010000010010000000100011;
ROM[37603] <= 32'b00000000010000010000000100010011;
ROM[37604] <= 32'b00000000010100010010000000100011;
ROM[37605] <= 32'b00000000010000010000000100010011;
ROM[37606] <= 32'b00000000011000010010000000100011;
ROM[37607] <= 32'b00000000010000010000000100010011;
ROM[37608] <= 32'b00000001010000000000001110010011;
ROM[37609] <= 32'b00000000100000111000001110010011;
ROM[37610] <= 32'b01000000011100010000001110110011;
ROM[37611] <= 32'b00000000011100000000001000110011;
ROM[37612] <= 32'b00000000001000000000000110110011;
ROM[37613] <= 32'b11000111100111101100000011101111;
ROM[37614] <= 32'b11111111110000010000000100010011;
ROM[37615] <= 32'b00000000000000010010001110000011;
ROM[37616] <= 32'b11111111110000010000000100010011;
ROM[37617] <= 32'b00000000000000010010010000000011;
ROM[37618] <= 32'b00000000011101000000001110110011;
ROM[37619] <= 32'b00000000011100010010000000100011;
ROM[37620] <= 32'b00000000010000010000000100010011;
ROM[37621] <= 32'b11111111110000010000000100010011;
ROM[37622] <= 32'b00000000000000010010001110000011;
ROM[37623] <= 32'b00000000000000111000001100010011;
ROM[37624] <= 32'b11111111110000010000000100010011;
ROM[37625] <= 32'b00000000000000010010001110000011;
ROM[37626] <= 32'b00000000110100110000010000110011;
ROM[37627] <= 32'b00000000011101000010000000100011;
ROM[37628] <= 32'b00000000100100000000001110010011;
ROM[37629] <= 32'b00000000011100010010000000100011;
ROM[37630] <= 32'b00000000010000010000000100010011;
ROM[37631] <= 32'b00000000110100101000010000110011;
ROM[37632] <= 32'b00000001100001000010001110000011;
ROM[37633] <= 32'b00000000011100010010000000100011;
ROM[37634] <= 32'b00000000010000010000000100010011;
ROM[37635] <= 32'b00000000011000000000001110010011;
ROM[37636] <= 32'b00000000011100010010000000100011;
ROM[37637] <= 32'b00000000010000010000000100010011;
ROM[37638] <= 32'b00000000010000000000001110010011;
ROM[37639] <= 32'b00000000011100010010000000100011;
ROM[37640] <= 32'b00000000010000010000000100010011;
ROM[37641] <= 32'b00000000000000100101001110110111;
ROM[37642] <= 32'b11000111000000111000001110010011;
ROM[37643] <= 32'b00000000111000111000001110110011;
ROM[37644] <= 32'b00000000011100010010000000100011;
ROM[37645] <= 32'b00000000010000010000000100010011;
ROM[37646] <= 32'b00000000001100010010000000100011;
ROM[37647] <= 32'b00000000010000010000000100010011;
ROM[37648] <= 32'b00000000010000010010000000100011;
ROM[37649] <= 32'b00000000010000010000000100010011;
ROM[37650] <= 32'b00000000010100010010000000100011;
ROM[37651] <= 32'b00000000010000010000000100010011;
ROM[37652] <= 32'b00000000011000010010000000100011;
ROM[37653] <= 32'b00000000010000010000000100010011;
ROM[37654] <= 32'b00000001010000000000001110010011;
ROM[37655] <= 32'b00000000100000111000001110010011;
ROM[37656] <= 32'b01000000011100010000001110110011;
ROM[37657] <= 32'b00000000011100000000001000110011;
ROM[37658] <= 32'b00000000001000000000000110110011;
ROM[37659] <= 32'b10111100000111101100000011101111;
ROM[37660] <= 32'b11111111110000010000000100010011;
ROM[37661] <= 32'b00000000000000010010001110000011;
ROM[37662] <= 32'b11111111110000010000000100010011;
ROM[37663] <= 32'b00000000000000010010010000000011;
ROM[37664] <= 32'b00000000011101000000001110110011;
ROM[37665] <= 32'b00000000011100010010000000100011;
ROM[37666] <= 32'b00000000010000010000000100010011;
ROM[37667] <= 32'b11111111110000010000000100010011;
ROM[37668] <= 32'b00000000000000010010001110000011;
ROM[37669] <= 32'b00000000000000111000001100010011;
ROM[37670] <= 32'b11111111110000010000000100010011;
ROM[37671] <= 32'b00000000000000010010001110000011;
ROM[37672] <= 32'b00000000110100110000010000110011;
ROM[37673] <= 32'b00000000011101000010000000100011;
ROM[37674] <= 32'b00000100001000000000001110010011;
ROM[37675] <= 32'b00000000011100010010000000100011;
ROM[37676] <= 32'b00000000010000010000000100010011;
ROM[37677] <= 32'b00000000110100101000010000110011;
ROM[37678] <= 32'b00000001100001000010001110000011;
ROM[37679] <= 32'b00000000011100010010000000100011;
ROM[37680] <= 32'b00000000010000010000000100010011;
ROM[37681] <= 32'b00000000011100000000001110010011;
ROM[37682] <= 32'b00000000011100010010000000100011;
ROM[37683] <= 32'b00000000010000010000000100010011;
ROM[37684] <= 32'b00000000010000000000001110010011;
ROM[37685] <= 32'b00000000011100010010000000100011;
ROM[37686] <= 32'b00000000010000010000000100010011;
ROM[37687] <= 32'b00000000000000100101001110110111;
ROM[37688] <= 32'b11010010100000111000001110010011;
ROM[37689] <= 32'b00000000111000111000001110110011;
ROM[37690] <= 32'b00000000011100010010000000100011;
ROM[37691] <= 32'b00000000010000010000000100010011;
ROM[37692] <= 32'b00000000001100010010000000100011;
ROM[37693] <= 32'b00000000010000010000000100010011;
ROM[37694] <= 32'b00000000010000010010000000100011;
ROM[37695] <= 32'b00000000010000010000000100010011;
ROM[37696] <= 32'b00000000010100010010000000100011;
ROM[37697] <= 32'b00000000010000010000000100010011;
ROM[37698] <= 32'b00000000011000010010000000100011;
ROM[37699] <= 32'b00000000010000010000000100010011;
ROM[37700] <= 32'b00000001010000000000001110010011;
ROM[37701] <= 32'b00000000100000111000001110010011;
ROM[37702] <= 32'b01000000011100010000001110110011;
ROM[37703] <= 32'b00000000011100000000001000110011;
ROM[37704] <= 32'b00000000001000000000000110110011;
ROM[37705] <= 32'b10110000100111101100000011101111;
ROM[37706] <= 32'b11111111110000010000000100010011;
ROM[37707] <= 32'b00000000000000010010001110000011;
ROM[37708] <= 32'b11111111110000010000000100010011;
ROM[37709] <= 32'b00000000000000010010010000000011;
ROM[37710] <= 32'b00000000011101000000001110110011;
ROM[37711] <= 32'b00000000011100010010000000100011;
ROM[37712] <= 32'b00000000010000010000000100010011;
ROM[37713] <= 32'b11111111110000010000000100010011;
ROM[37714] <= 32'b00000000000000010010001110000011;
ROM[37715] <= 32'b00000000000000111000001100010011;
ROM[37716] <= 32'b11111111110000010000000100010011;
ROM[37717] <= 32'b00000000000000010010001110000011;
ROM[37718] <= 32'b00000000110100110000010000110011;
ROM[37719] <= 32'b00000000011101000010000000100011;
ROM[37720] <= 32'b00000011100000000000001110010011;
ROM[37721] <= 32'b00000000011100010010000000100011;
ROM[37722] <= 32'b00000000010000010000000100010011;
ROM[37723] <= 32'b00000000110100101000010000110011;
ROM[37724] <= 32'b00000001100001000010001110000011;
ROM[37725] <= 32'b00000000011100010010000000100011;
ROM[37726] <= 32'b00000000010000010000000100010011;
ROM[37727] <= 32'b00000000100000000000001110010011;
ROM[37728] <= 32'b00000000011100010010000000100011;
ROM[37729] <= 32'b00000000010000010000000100010011;
ROM[37730] <= 32'b00000000010000000000001110010011;
ROM[37731] <= 32'b00000000011100010010000000100011;
ROM[37732] <= 32'b00000000010000010000000100010011;
ROM[37733] <= 32'b00000000000000100101001110110111;
ROM[37734] <= 32'b11011110000000111000001110010011;
ROM[37735] <= 32'b00000000111000111000001110110011;
ROM[37736] <= 32'b00000000011100010010000000100011;
ROM[37737] <= 32'b00000000010000010000000100010011;
ROM[37738] <= 32'b00000000001100010010000000100011;
ROM[37739] <= 32'b00000000010000010000000100010011;
ROM[37740] <= 32'b00000000010000010010000000100011;
ROM[37741] <= 32'b00000000010000010000000100010011;
ROM[37742] <= 32'b00000000010100010010000000100011;
ROM[37743] <= 32'b00000000010000010000000100010011;
ROM[37744] <= 32'b00000000011000010010000000100011;
ROM[37745] <= 32'b00000000010000010000000100010011;
ROM[37746] <= 32'b00000001010000000000001110010011;
ROM[37747] <= 32'b00000000100000111000001110010011;
ROM[37748] <= 32'b01000000011100010000001110110011;
ROM[37749] <= 32'b00000000011100000000001000110011;
ROM[37750] <= 32'b00000000001000000000000110110011;
ROM[37751] <= 32'b10100101000111101100000011101111;
ROM[37752] <= 32'b11111111110000010000000100010011;
ROM[37753] <= 32'b00000000000000010010001110000011;
ROM[37754] <= 32'b11111111110000010000000100010011;
ROM[37755] <= 32'b00000000000000010010010000000011;
ROM[37756] <= 32'b00000000011101000000001110110011;
ROM[37757] <= 32'b00000000011100010010000000100011;
ROM[37758] <= 32'b00000000010000010000000100010011;
ROM[37759] <= 32'b11111111110000010000000100010011;
ROM[37760] <= 32'b00000000000000010010001110000011;
ROM[37761] <= 32'b00000000000000111000001100010011;
ROM[37762] <= 32'b11111111110000010000000100010011;
ROM[37763] <= 32'b00000000000000010010001110000011;
ROM[37764] <= 32'b00000000110100110000010000110011;
ROM[37765] <= 32'b00000000011101000010000000100011;
ROM[37766] <= 32'b00000010001100000000001110010011;
ROM[37767] <= 32'b00000000011100010010000000100011;
ROM[37768] <= 32'b00000000010000010000000100010011;
ROM[37769] <= 32'b00000000110100101000010000110011;
ROM[37770] <= 32'b00000001100001000010001110000011;
ROM[37771] <= 32'b00000000011100010010000000100011;
ROM[37772] <= 32'b00000000010000010000000100010011;
ROM[37773] <= 32'b00000000100100000000001110010011;
ROM[37774] <= 32'b00000000011100010010000000100011;
ROM[37775] <= 32'b00000000010000010000000100010011;
ROM[37776] <= 32'b00000000010000000000001110010011;
ROM[37777] <= 32'b00000000011100010010000000100011;
ROM[37778] <= 32'b00000000010000010000000100010011;
ROM[37779] <= 32'b00000000000000100101001110110111;
ROM[37780] <= 32'b11101001100000111000001110010011;
ROM[37781] <= 32'b00000000111000111000001110110011;
ROM[37782] <= 32'b00000000011100010010000000100011;
ROM[37783] <= 32'b00000000010000010000000100010011;
ROM[37784] <= 32'b00000000001100010010000000100011;
ROM[37785] <= 32'b00000000010000010000000100010011;
ROM[37786] <= 32'b00000000010000010010000000100011;
ROM[37787] <= 32'b00000000010000010000000100010011;
ROM[37788] <= 32'b00000000010100010010000000100011;
ROM[37789] <= 32'b00000000010000010000000100010011;
ROM[37790] <= 32'b00000000011000010010000000100011;
ROM[37791] <= 32'b00000000010000010000000100010011;
ROM[37792] <= 32'b00000001010000000000001110010011;
ROM[37793] <= 32'b00000000100000111000001110010011;
ROM[37794] <= 32'b01000000011100010000001110110011;
ROM[37795] <= 32'b00000000011100000000001000110011;
ROM[37796] <= 32'b00000000001000000000000110110011;
ROM[37797] <= 32'b10011001100111101100000011101111;
ROM[37798] <= 32'b11111111110000010000000100010011;
ROM[37799] <= 32'b00000000000000010010001110000011;
ROM[37800] <= 32'b11111111110000010000000100010011;
ROM[37801] <= 32'b00000000000000010010010000000011;
ROM[37802] <= 32'b00000000011101000000001110110011;
ROM[37803] <= 32'b00000000011100010010000000100011;
ROM[37804] <= 32'b00000000010000010000000100010011;
ROM[37805] <= 32'b11111111110000010000000100010011;
ROM[37806] <= 32'b00000000000000010010001110000011;
ROM[37807] <= 32'b00000000000000111000001100010011;
ROM[37808] <= 32'b11111111110000010000000100010011;
ROM[37809] <= 32'b00000000000000010010001110000011;
ROM[37810] <= 32'b00000000110100110000010000110011;
ROM[37811] <= 32'b00000000011101000010000000100011;
ROM[37812] <= 32'b00000000000000000000001110010011;
ROM[37813] <= 32'b00000000011100010010000000100011;
ROM[37814] <= 32'b00000000010000010000000100010011;
ROM[37815] <= 32'b11111111110000010000000100010011;
ROM[37816] <= 32'b00000000000000010010001110000011;
ROM[37817] <= 32'b00000000110100101000010000110011;
ROM[37818] <= 32'b00000010011101000010000000100011;
ROM[37819] <= 32'b00000000010100010010000000100011;
ROM[37820] <= 32'b00000000010000010000000100010011;
ROM[37821] <= 32'b00000000000000100101001110110111;
ROM[37822] <= 32'b11110100000000111000001110010011;
ROM[37823] <= 32'b00000000111000111000001110110011;
ROM[37824] <= 32'b00000000011100010010000000100011;
ROM[37825] <= 32'b00000000010000010000000100010011;
ROM[37826] <= 32'b00000000001100010010000000100011;
ROM[37827] <= 32'b00000000010000010000000100010011;
ROM[37828] <= 32'b00000000010000010010000000100011;
ROM[37829] <= 32'b00000000010000010000000100010011;
ROM[37830] <= 32'b00000000010100010010000000100011;
ROM[37831] <= 32'b00000000010000010000000100010011;
ROM[37832] <= 32'b00000000011000010010000000100011;
ROM[37833] <= 32'b00000000010000010000000100010011;
ROM[37834] <= 32'b00000001010000000000001110010011;
ROM[37835] <= 32'b00000000010000111000001110010011;
ROM[37836] <= 32'b01000000011100010000001110110011;
ROM[37837] <= 32'b00000000011100000000001000110011;
ROM[37838] <= 32'b00000000001000000000000110110011;
ROM[37839] <= 32'b00011000110100000000000011101111;
ROM[37840] <= 32'b11111111110000010000000100010011;
ROM[37841] <= 32'b00000000000000010010001110000011;
ROM[37842] <= 32'b00000000011101100010000000100011;
ROM[37843] <= 32'b00000000010100010010000000100011;
ROM[37844] <= 32'b00000000010000010000000100010011;
ROM[37845] <= 32'b00000001010000000000001110010011;
ROM[37846] <= 32'b01000000011100011000001110110011;
ROM[37847] <= 32'b00000000000000111010000010000011;
ROM[37848] <= 32'b11111111110000010000000100010011;
ROM[37849] <= 32'b00000000000000010010001110000011;
ROM[37850] <= 32'b00000000011100100010000000100011;
ROM[37851] <= 32'b00000000010000100000000100010011;
ROM[37852] <= 32'b00000001010000000000001110010011;
ROM[37853] <= 32'b01000000011100011000001110110011;
ROM[37854] <= 32'b00000000010000111010000110000011;
ROM[37855] <= 32'b00000000100000111010001000000011;
ROM[37856] <= 32'b00000000110000111010001010000011;
ROM[37857] <= 32'b00000001000000111010001100000011;
ROM[37858] <= 32'b00000000000000001000000011100111;
ROM[37859] <= 32'b00000000000000010010000000100011;
ROM[37860] <= 32'b00000000010000010000000100010011;
ROM[37861] <= 32'b00000000000000010010000000100011;
ROM[37862] <= 32'b00000000010000010000000100010011;
ROM[37863] <= 32'b00000000000000100010001110000011;
ROM[37864] <= 32'b00000000011100010010000000100011;
ROM[37865] <= 32'b00000000010000010000000100010011;
ROM[37866] <= 32'b11111111110000010000000100010011;
ROM[37867] <= 32'b00000000000000010010001110000011;
ROM[37868] <= 32'b00000000000000111000001010010011;
ROM[37869] <= 32'b00000000000000000000001110010011;
ROM[37870] <= 32'b00000000011100010010000000100011;
ROM[37871] <= 32'b00000000010000010000000100010011;
ROM[37872] <= 32'b11111111110000010000000100010011;
ROM[37873] <= 32'b00000000000000010010001110000011;
ROM[37874] <= 32'b00000000011100011010000000100011;
ROM[37875] <= 32'b00000000000000011010001110000011;
ROM[37876] <= 32'b00000000011100010010000000100011;
ROM[37877] <= 32'b00000000010000010000000100010011;
ROM[37878] <= 32'b00000000110100101000010000110011;
ROM[37879] <= 32'b00000000010001000010001110000011;
ROM[37880] <= 32'b00000000011100010010000000100011;
ROM[37881] <= 32'b00000000010000010000000100010011;
ROM[37882] <= 32'b11111111110000010000000100010011;
ROM[37883] <= 32'b00000000000000010010001110000011;
ROM[37884] <= 32'b11111111110000010000000100010011;
ROM[37885] <= 32'b00000000000000010010010000000011;
ROM[37886] <= 32'b00000000011101000010001110110011;
ROM[37887] <= 32'b00000000011100010010000000100011;
ROM[37888] <= 32'b00000000010000010000000100010011;
ROM[37889] <= 32'b11111111110000010000000100010011;
ROM[37890] <= 32'b00000000000000010010001110000011;
ROM[37891] <= 32'b01000000011100000000001110110011;
ROM[37892] <= 32'b00000000000100111000001110010011;
ROM[37893] <= 32'b00000000011100010010000000100011;
ROM[37894] <= 32'b00000000010000010000000100010011;
ROM[37895] <= 32'b11111111110000010000000100010011;
ROM[37896] <= 32'b00000000000000010010001110000011;
ROM[37897] <= 32'b00000000000000111000101001100011;
ROM[37898] <= 32'b00000000000000100101001110110111;
ROM[37899] <= 32'b00011001100000111000001110010011;
ROM[37900] <= 32'b00000000111000111000001110110011;
ROM[37901] <= 32'b00000000000000111000000011100111;
ROM[37902] <= 32'b00000000110100101000010000110011;
ROM[37903] <= 32'b00000001010001000010001110000011;
ROM[37904] <= 32'b00000000011100010010000000100011;
ROM[37905] <= 32'b00000000010000010000000100010011;
ROM[37906] <= 32'b00000000000000011010001110000011;
ROM[37907] <= 32'b00000000011100010010000000100011;
ROM[37908] <= 32'b00000000010000010000000100010011;
ROM[37909] <= 32'b00000000010000000000001110010011;
ROM[37910] <= 32'b00000000011100010010000000100011;
ROM[37911] <= 32'b00000000010000010000000100010011;
ROM[37912] <= 32'b00000000000000100101001110110111;
ROM[37913] <= 32'b00001010110000111000001110010011;
ROM[37914] <= 32'b00000000111000111000001110110011;
ROM[37915] <= 32'b00000000011100010010000000100011;
ROM[37916] <= 32'b00000000010000010000000100010011;
ROM[37917] <= 32'b00000000001100010010000000100011;
ROM[37918] <= 32'b00000000010000010000000100010011;
ROM[37919] <= 32'b00000000010000010010000000100011;
ROM[37920] <= 32'b00000000010000010000000100010011;
ROM[37921] <= 32'b00000000010100010010000000100011;
ROM[37922] <= 32'b00000000010000010000000100010011;
ROM[37923] <= 32'b00000000011000010010000000100011;
ROM[37924] <= 32'b00000000010000010000000100010011;
ROM[37925] <= 32'b00000001010000000000001110010011;
ROM[37926] <= 32'b00000000100000111000001110010011;
ROM[37927] <= 32'b01000000011100010000001110110011;
ROM[37928] <= 32'b00000000011100000000001000110011;
ROM[37929] <= 32'b00000000001000000000000110110011;
ROM[37930] <= 32'b11111000010011101100000011101111;
ROM[37931] <= 32'b11111111110000010000000100010011;
ROM[37932] <= 32'b00000000000000010010001110000011;
ROM[37933] <= 32'b11111111110000010000000100010011;
ROM[37934] <= 32'b00000000000000010010010000000011;
ROM[37935] <= 32'b00000000011101000000001110110011;
ROM[37936] <= 32'b00000000011100010010000000100011;
ROM[37937] <= 32'b00000000010000010000000100010011;
ROM[37938] <= 32'b11111111110000010000000100010011;
ROM[37939] <= 32'b00000000000000010010001110000011;
ROM[37940] <= 32'b00000000000000111000001100010011;
ROM[37941] <= 32'b00000000110100110000010000110011;
ROM[37942] <= 32'b00000000000001000010001110000011;
ROM[37943] <= 32'b00000000011100010010000000100011;
ROM[37944] <= 32'b00000000010000010000000100010011;
ROM[37945] <= 32'b11111111110000010000000100010011;
ROM[37946] <= 32'b00000000000000010010001110000011;
ROM[37947] <= 32'b00000000011100011010001000100011;
ROM[37948] <= 32'b00000000010000011010001110000011;
ROM[37949] <= 32'b00000000011100010010000000100011;
ROM[37950] <= 32'b00000000010000010000000100010011;
ROM[37951] <= 32'b00000000000000100101001110110111;
ROM[37952] <= 32'b00010100100000111000001110010011;
ROM[37953] <= 32'b00000000111000111000001110110011;
ROM[37954] <= 32'b00000000011100010010000000100011;
ROM[37955] <= 32'b00000000010000010000000100010011;
ROM[37956] <= 32'b00000000001100010010000000100011;
ROM[37957] <= 32'b00000000010000010000000100010011;
ROM[37958] <= 32'b00000000010000010010000000100011;
ROM[37959] <= 32'b00000000010000010000000100010011;
ROM[37960] <= 32'b00000000010100010010000000100011;
ROM[37961] <= 32'b00000000010000010000000100010011;
ROM[37962] <= 32'b00000000011000010010000000100011;
ROM[37963] <= 32'b00000000010000010000000100010011;
ROM[37964] <= 32'b00000001010000000000001110010011;
ROM[37965] <= 32'b00000000010000111000001110010011;
ROM[37966] <= 32'b01000000011100010000001110110011;
ROM[37967] <= 32'b00000000011100000000001000110011;
ROM[37968] <= 32'b00000000001000000000000110110011;
ROM[37969] <= 32'b11111100110111011010000011101111;
ROM[37970] <= 32'b11111111110000010000000100010011;
ROM[37971] <= 32'b00000000000000010010001110000011;
ROM[37972] <= 32'b00000000011101100010000000100011;
ROM[37973] <= 32'b00000000000000011010001110000011;
ROM[37974] <= 32'b00000000011100010010000000100011;
ROM[37975] <= 32'b00000000010000010000000100010011;
ROM[37976] <= 32'b00000000000100000000001110010011;
ROM[37977] <= 32'b00000000011100010010000000100011;
ROM[37978] <= 32'b00000000010000010000000100010011;
ROM[37979] <= 32'b11111111110000010000000100010011;
ROM[37980] <= 32'b00000000000000010010001110000011;
ROM[37981] <= 32'b11111111110000010000000100010011;
ROM[37982] <= 32'b00000000000000010010010000000011;
ROM[37983] <= 32'b00000000011101000000001110110011;
ROM[37984] <= 32'b00000000011100010010000000100011;
ROM[37985] <= 32'b00000000010000010000000100010011;
ROM[37986] <= 32'b11111111110000010000000100010011;
ROM[37987] <= 32'b00000000000000010010001110000011;
ROM[37988] <= 32'b00000000011100011010000000100011;
ROM[37989] <= 32'b11100011100111111111000011101111;
ROM[37990] <= 32'b00000000010100010010000000100011;
ROM[37991] <= 32'b00000000010000010000000100010011;
ROM[37992] <= 32'b00000000000000100101001110110111;
ROM[37993] <= 32'b00011110110000111000001110010011;
ROM[37994] <= 32'b00000000111000111000001110110011;
ROM[37995] <= 32'b00000000011100010010000000100011;
ROM[37996] <= 32'b00000000010000010000000100010011;
ROM[37997] <= 32'b00000000001100010010000000100011;
ROM[37998] <= 32'b00000000010000010000000100010011;
ROM[37999] <= 32'b00000000010000010010000000100011;
ROM[38000] <= 32'b00000000010000010000000100010011;
ROM[38001] <= 32'b00000000010100010010000000100011;
ROM[38002] <= 32'b00000000010000010000000100010011;
ROM[38003] <= 32'b00000000011000010010000000100011;
ROM[38004] <= 32'b00000000010000010000000100010011;
ROM[38005] <= 32'b00000001010000000000001110010011;
ROM[38006] <= 32'b00000000010000111000001110010011;
ROM[38007] <= 32'b01000000011100010000001110110011;
ROM[38008] <= 32'b00000000011100000000001000110011;
ROM[38009] <= 32'b00000000001000000000000110110011;
ROM[38010] <= 32'b10010111010111101110000011101111;
ROM[38011] <= 32'b11111111110000010000000100010011;
ROM[38012] <= 32'b00000000000000010010001110000011;
ROM[38013] <= 32'b00000000011101100010000000100011;
ROM[38014] <= 32'b00000000000000000000001110010011;
ROM[38015] <= 32'b00000000011100010010000000100011;
ROM[38016] <= 32'b00000000010000010000000100010011;
ROM[38017] <= 32'b00000001010000000000001110010011;
ROM[38018] <= 32'b01000000011100011000001110110011;
ROM[38019] <= 32'b00000000000000111010000010000011;
ROM[38020] <= 32'b11111111110000010000000100010011;
ROM[38021] <= 32'b00000000000000010010001110000011;
ROM[38022] <= 32'b00000000011100100010000000100011;
ROM[38023] <= 32'b00000000010000100000000100010011;
ROM[38024] <= 32'b00000001010000000000001110010011;
ROM[38025] <= 32'b01000000011100011000001110110011;
ROM[38026] <= 32'b00000000010000111010000110000011;
ROM[38027] <= 32'b00000000100000111010001000000011;
ROM[38028] <= 32'b00000000110000111010001010000011;
ROM[38029] <= 32'b00000001000000111010001100000011;
ROM[38030] <= 32'b00000000000000001000000011100111;
ROM[38031] <= 32'b00000000000000010010000000100011;
ROM[38032] <= 32'b00000000010000010000000100010011;
ROM[38033] <= 32'b00000000000000010010000000100011;
ROM[38034] <= 32'b00000000010000010000000100010011;
ROM[38035] <= 32'b00000000000000010010000000100011;
ROM[38036] <= 32'b00000000010000010000000100010011;
ROM[38037] <= 32'b00000000000000100010001110000011;
ROM[38038] <= 32'b00000000011100010010000000100011;
ROM[38039] <= 32'b00000000010000010000000100010011;
ROM[38040] <= 32'b11111111110000010000000100010011;
ROM[38041] <= 32'b00000000000000010010001110000011;
ROM[38042] <= 32'b00000000000000111000001010010011;
ROM[38043] <= 32'b00000000000000000000001110010011;
ROM[38044] <= 32'b00000000011100010010000000100011;
ROM[38045] <= 32'b00000000010000010000000100010011;
ROM[38046] <= 32'b11111111110000010000000100010011;
ROM[38047] <= 32'b00000000000000010010001110000011;
ROM[38048] <= 32'b00000000011100011010000000100011;
ROM[38049] <= 32'b00000000000000011010001110000011;
ROM[38050] <= 32'b00000000011100010010000000100011;
ROM[38051] <= 32'b00000000010000010000000100010011;
ROM[38052] <= 32'b11111111110000010000000100010011;
ROM[38053] <= 32'b00000000000000010010001110000011;
ROM[38054] <= 32'b01000000011100000000001110110011;
ROM[38055] <= 32'b00000000000100111000001110010011;
ROM[38056] <= 32'b00000000011100010010000000100011;
ROM[38057] <= 32'b00000000010000010000000100010011;
ROM[38058] <= 32'b11111111110000010000000100010011;
ROM[38059] <= 32'b00000000000000010010001110000011;
ROM[38060] <= 32'b01000000011100000000001110110011;
ROM[38061] <= 32'b00000000000100111000001110010011;
ROM[38062] <= 32'b00000000011100010010000000100011;
ROM[38063] <= 32'b00000000010000010000000100010011;
ROM[38064] <= 32'b11111111110000010000000100010011;
ROM[38065] <= 32'b00000000000000010010001110000011;
ROM[38066] <= 32'b00000000000000111000101001100011;
ROM[38067] <= 32'b00000000000000100101001110110111;
ROM[38068] <= 32'b01011111010000111000001110010011;
ROM[38069] <= 32'b00000000111000111000001110110011;
ROM[38070] <= 32'b00000000000000111000000011100111;
ROM[38071] <= 32'b00000000110100101000010000110011;
ROM[38072] <= 32'b00000001100001000010001110000011;
ROM[38073] <= 32'b00000000011100010010000000100011;
ROM[38074] <= 32'b00000000010000010000000100010011;
ROM[38075] <= 32'b00000000110100101000010000110011;
ROM[38076] <= 32'b00000010000001000010001110000011;
ROM[38077] <= 32'b00000000011100010010000000100011;
ROM[38078] <= 32'b00000000010000010000000100010011;
ROM[38079] <= 32'b00000000010000000000001110010011;
ROM[38080] <= 32'b00000000011100010010000000100011;
ROM[38081] <= 32'b00000000010000010000000100010011;
ROM[38082] <= 32'b00000000000000100101001110110111;
ROM[38083] <= 32'b00110101010000111000001110010011;
ROM[38084] <= 32'b00000000111000111000001110110011;
ROM[38085] <= 32'b00000000011100010010000000100011;
ROM[38086] <= 32'b00000000010000010000000100010011;
ROM[38087] <= 32'b00000000001100010010000000100011;
ROM[38088] <= 32'b00000000010000010000000100010011;
ROM[38089] <= 32'b00000000010000010010000000100011;
ROM[38090] <= 32'b00000000010000010000000100010011;
ROM[38091] <= 32'b00000000010100010010000000100011;
ROM[38092] <= 32'b00000000010000010000000100010011;
ROM[38093] <= 32'b00000000011000010010000000100011;
ROM[38094] <= 32'b00000000010000010000000100010011;
ROM[38095] <= 32'b00000001010000000000001110010011;
ROM[38096] <= 32'b00000000100000111000001110010011;
ROM[38097] <= 32'b01000000011100010000001110110011;
ROM[38098] <= 32'b00000000011100000000001000110011;
ROM[38099] <= 32'b00000000001000000000000110110011;
ROM[38100] <= 32'b11001101110011101100000011101111;
ROM[38101] <= 32'b11111111110000010000000100010011;
ROM[38102] <= 32'b00000000000000010010001110000011;
ROM[38103] <= 32'b11111111110000010000000100010011;
ROM[38104] <= 32'b00000000000000010010010000000011;
ROM[38105] <= 32'b00000000011101000000001110110011;
ROM[38106] <= 32'b00000000011100010010000000100011;
ROM[38107] <= 32'b00000000010000010000000100010011;
ROM[38108] <= 32'b11111111110000010000000100010011;
ROM[38109] <= 32'b00000000000000010010001110000011;
ROM[38110] <= 32'b00000000000000111000001100010011;
ROM[38111] <= 32'b00000000110100110000010000110011;
ROM[38112] <= 32'b00000000000001000010001110000011;
ROM[38113] <= 32'b00000000011100010010000000100011;
ROM[38114] <= 32'b00000000010000010000000100010011;
ROM[38115] <= 32'b11111111110000010000000100010011;
ROM[38116] <= 32'b00000000000000010010001110000011;
ROM[38117] <= 32'b00000000011100011010001000100011;
ROM[38118] <= 32'b00000000110100101000010000110011;
ROM[38119] <= 32'b00000001110001000010001110000011;
ROM[38120] <= 32'b00000000011100010010000000100011;
ROM[38121] <= 32'b00000000010000010000000100010011;
ROM[38122] <= 32'b00000000110100101000010000110011;
ROM[38123] <= 32'b00000010000001000010001110000011;
ROM[38124] <= 32'b00000000011100010010000000100011;
ROM[38125] <= 32'b00000000010000010000000100010011;
ROM[38126] <= 32'b00000000010000000000001110010011;
ROM[38127] <= 32'b00000000011100010010000000100011;
ROM[38128] <= 32'b00000000010000010000000100010011;
ROM[38129] <= 32'b00000000000000100101001110110111;
ROM[38130] <= 32'b01000001000000111000001110010011;
ROM[38131] <= 32'b00000000111000111000001110110011;
ROM[38132] <= 32'b00000000011100010010000000100011;
ROM[38133] <= 32'b00000000010000010000000100010011;
ROM[38134] <= 32'b00000000001100010010000000100011;
ROM[38135] <= 32'b00000000010000010000000100010011;
ROM[38136] <= 32'b00000000010000010010000000100011;
ROM[38137] <= 32'b00000000010000010000000100010011;
ROM[38138] <= 32'b00000000010100010010000000100011;
ROM[38139] <= 32'b00000000010000010000000100010011;
ROM[38140] <= 32'b00000000011000010010000000100011;
ROM[38141] <= 32'b00000000010000010000000100010011;
ROM[38142] <= 32'b00000001010000000000001110010011;
ROM[38143] <= 32'b00000000100000111000001110010011;
ROM[38144] <= 32'b01000000011100010000001110110011;
ROM[38145] <= 32'b00000000011100000000001000110011;
ROM[38146] <= 32'b00000000001000000000000110110011;
ROM[38147] <= 32'b11000010000011101100000011101111;
ROM[38148] <= 32'b11111111110000010000000100010011;
ROM[38149] <= 32'b00000000000000010010001110000011;
ROM[38150] <= 32'b11111111110000010000000100010011;
ROM[38151] <= 32'b00000000000000010010010000000011;
ROM[38152] <= 32'b00000000011101000000001110110011;
ROM[38153] <= 32'b00000000011100010010000000100011;
ROM[38154] <= 32'b00000000010000010000000100010011;
ROM[38155] <= 32'b11111111110000010000000100010011;
ROM[38156] <= 32'b00000000000000010010001110000011;
ROM[38157] <= 32'b00000000000000111000001100010011;
ROM[38158] <= 32'b00000000110100110000010000110011;
ROM[38159] <= 32'b00000000000001000010001110000011;
ROM[38160] <= 32'b00000000011100010010000000100011;
ROM[38161] <= 32'b00000000010000010000000100010011;
ROM[38162] <= 32'b11111111110000010000000100010011;
ROM[38163] <= 32'b00000000000000010010001110000011;
ROM[38164] <= 32'b00000000011100011010010000100011;
ROM[38165] <= 32'b00000000110100101000010000110011;
ROM[38166] <= 32'b00000010000001000010001110000011;
ROM[38167] <= 32'b00000000011100010010000000100011;
ROM[38168] <= 32'b00000000010000010000000100010011;
ROM[38169] <= 32'b00000000000100000000001110010011;
ROM[38170] <= 32'b00000000011100010010000000100011;
ROM[38171] <= 32'b00000000010000010000000100010011;
ROM[38172] <= 32'b11111111110000010000000100010011;
ROM[38173] <= 32'b00000000000000010010001110000011;
ROM[38174] <= 32'b11111111110000010000000100010011;
ROM[38175] <= 32'b00000000000000010010010000000011;
ROM[38176] <= 32'b00000000011101000000001110110011;
ROM[38177] <= 32'b00000000011100010010000000100011;
ROM[38178] <= 32'b00000000010000010000000100010011;
ROM[38179] <= 32'b11111111110000010000000100010011;
ROM[38180] <= 32'b00000000000000010010001110000011;
ROM[38181] <= 32'b00000000110100101000010000110011;
ROM[38182] <= 32'b00000010011101000010000000100011;
ROM[38183] <= 32'b00000000110100101000010000110011;
ROM[38184] <= 32'b00000010000001000010001110000011;
ROM[38185] <= 32'b00000000011100010010000000100011;
ROM[38186] <= 32'b00000000010000010000000100010011;
ROM[38187] <= 32'b00000000001000000000001110010011;
ROM[38188] <= 32'b00000000011100010010000000100011;
ROM[38189] <= 32'b00000000010000010000000100010011;
ROM[38190] <= 32'b11111111110000010000000100010011;
ROM[38191] <= 32'b00000000000000010010001110000011;
ROM[38192] <= 32'b11111111110000010000000100010011;
ROM[38193] <= 32'b00000000000000010010010000000011;
ROM[38194] <= 32'b00000000011101000010010010110011;
ROM[38195] <= 32'b00000000100000111010010100110011;
ROM[38196] <= 32'b00000000101001001000001110110011;
ROM[38197] <= 32'b00000000000100111000001110010011;
ROM[38198] <= 32'b00000000000100111111001110010011;
ROM[38199] <= 32'b00000000011100010010000000100011;
ROM[38200] <= 32'b00000000010000010000000100010011;
ROM[38201] <= 32'b11111111110000010000000100010011;
ROM[38202] <= 32'b00000000000000010010001110000011;
ROM[38203] <= 32'b00000000000000111000101001100011;
ROM[38204] <= 32'b00000000000000100101001110110111;
ROM[38205] <= 32'b01010000010000111000001110010011;
ROM[38206] <= 32'b00000000111000111000001110110011;
ROM[38207] <= 32'b00000000000000111000000011100111;
ROM[38208] <= 32'b00000010000000000000000011101111;
ROM[38209] <= 32'b00000000000000000000001110010011;
ROM[38210] <= 32'b00000000011100010010000000100011;
ROM[38211] <= 32'b00000000010000010000000100010011;
ROM[38212] <= 32'b11111111110000010000000100010011;
ROM[38213] <= 32'b00000000000000010010001110000011;
ROM[38214] <= 32'b00000000110100101000010000110011;
ROM[38215] <= 32'b00000010011101000010000000100011;
ROM[38216] <= 32'b00000000010100010010000000100011;
ROM[38217] <= 32'b00000000010000010000000100010011;
ROM[38218] <= 32'b00000000010000011010001110000011;
ROM[38219] <= 32'b00000000011100010010000000100011;
ROM[38220] <= 32'b00000000010000010000000100010011;
ROM[38221] <= 32'b00000000100000011010001110000011;
ROM[38222] <= 32'b00000000011100010010000000100011;
ROM[38223] <= 32'b00000000010000010000000100010011;
ROM[38224] <= 32'b00000000000000100101001110110111;
ROM[38225] <= 32'b01011000110000111000001110010011;
ROM[38226] <= 32'b00000000111000111000001110110011;
ROM[38227] <= 32'b00000000011100010010000000100011;
ROM[38228] <= 32'b00000000010000010000000100010011;
ROM[38229] <= 32'b00000000001100010010000000100011;
ROM[38230] <= 32'b00000000010000010000000100010011;
ROM[38231] <= 32'b00000000010000010010000000100011;
ROM[38232] <= 32'b00000000010000010000000100010011;
ROM[38233] <= 32'b00000000010100010010000000100011;
ROM[38234] <= 32'b00000000010000010000000100010011;
ROM[38235] <= 32'b00000000011000010010000000100011;
ROM[38236] <= 32'b00000000010000010000000100010011;
ROM[38237] <= 32'b00000001010000000000001110010011;
ROM[38238] <= 32'b00000000110000111000001110010011;
ROM[38239] <= 32'b01000000011100010000001110110011;
ROM[38240] <= 32'b00000000011100000000001000110011;
ROM[38241] <= 32'b00000000001000000000000110110011;
ROM[38242] <= 32'b01010110000100000000000011101111;
ROM[38243] <= 32'b11111111110000010000000100010011;
ROM[38244] <= 32'b00000000000000010010001110000011;
ROM[38245] <= 32'b01000000011100000000001110110011;
ROM[38246] <= 32'b00000000000100111000001110010011;
ROM[38247] <= 32'b00000000011100010010000000100011;
ROM[38248] <= 32'b00000000010000010000000100010011;
ROM[38249] <= 32'b11111111110000010000000100010011;
ROM[38250] <= 32'b00000000000000010010001110000011;
ROM[38251] <= 32'b00000000000000111000101001100011;
ROM[38252] <= 32'b00000000000000100101001110110111;
ROM[38253] <= 32'b01011100010000111000001110010011;
ROM[38254] <= 32'b00000000111000111000001110110011;
ROM[38255] <= 32'b00000000000000111000000011100111;
ROM[38256] <= 32'b00000011000000000000000011101111;
ROM[38257] <= 32'b00000000000100000000001110010011;
ROM[38258] <= 32'b00000000011100010010000000100011;
ROM[38259] <= 32'b00000000010000010000000100010011;
ROM[38260] <= 32'b11111111110000010000000100010011;
ROM[38261] <= 32'b00000000000000010010001110000011;
ROM[38262] <= 32'b01000000011100000000001110110011;
ROM[38263] <= 32'b00000000011100010010000000100011;
ROM[38264] <= 32'b00000000010000010000000100010011;
ROM[38265] <= 32'b11111111110000010000000100010011;
ROM[38266] <= 32'b00000000000000010010001110000011;
ROM[38267] <= 32'b00000000011100011010000000100011;
ROM[38268] <= 32'b11001001010111111111000011101111;
ROM[38269] <= 32'b00000000010000011010001110000011;
ROM[38270] <= 32'b00000000011100010010000000100011;
ROM[38271] <= 32'b00000000010000010000000100010011;
ROM[38272] <= 32'b11111111110000010000000100010011;
ROM[38273] <= 32'b00000000000000010010001110000011;
ROM[38274] <= 32'b00000000110100101000010000110011;
ROM[38275] <= 32'b00000000011101000010011000100011;
ROM[38276] <= 32'b00000000100000011010001110000011;
ROM[38277] <= 32'b00000000011100010010000000100011;
ROM[38278] <= 32'b00000000010000010000000100010011;
ROM[38279] <= 32'b11111111110000010000000100010011;
ROM[38280] <= 32'b00000000000000010010001110000011;
ROM[38281] <= 32'b00000000110100101000010000110011;
ROM[38282] <= 32'b00000000011101000010100000100011;
ROM[38283] <= 32'b00000000000000000000001110010011;
ROM[38284] <= 32'b00000000011100010010000000100011;
ROM[38285] <= 32'b00000000010000010000000100010011;
ROM[38286] <= 32'b00000001010000000000001110010011;
ROM[38287] <= 32'b01000000011100011000001110110011;
ROM[38288] <= 32'b00000000000000111010000010000011;
ROM[38289] <= 32'b11111111110000010000000100010011;
ROM[38290] <= 32'b00000000000000010010001110000011;
ROM[38291] <= 32'b00000000011100100010000000100011;
ROM[38292] <= 32'b00000000010000100000000100010011;
ROM[38293] <= 32'b00000001010000000000001110010011;
ROM[38294] <= 32'b01000000011100011000001110110011;
ROM[38295] <= 32'b00000000010000111010000110000011;
ROM[38296] <= 32'b00000000100000111010001000000011;
ROM[38297] <= 32'b00000000110000111010001010000011;
ROM[38298] <= 32'b00000001000000111010001100000011;
ROM[38299] <= 32'b00000000000000001000000011100111;
ROM[38300] <= 32'b00000000000000100010001110000011;
ROM[38301] <= 32'b00000000011100010010000000100011;
ROM[38302] <= 32'b00000000010000010000000100010011;
ROM[38303] <= 32'b11111111110000010000000100010011;
ROM[38304] <= 32'b00000000000000010010001110000011;
ROM[38305] <= 32'b00000000000000111000001010010011;
ROM[38306] <= 32'b00000000000100000000001110010011;
ROM[38307] <= 32'b00000000011100010010000000100011;
ROM[38308] <= 32'b00000000010000010000000100010011;
ROM[38309] <= 32'b11111111110000010000000100010011;
ROM[38310] <= 32'b00000000000000010010001110000011;
ROM[38311] <= 32'b01000000011100000000001110110011;
ROM[38312] <= 32'b00000000011100010010000000100011;
ROM[38313] <= 32'b00000000010000010000000100010011;
ROM[38314] <= 32'b00000000000000100101001110110111;
ROM[38315] <= 32'b01101111010000111000001110010011;
ROM[38316] <= 32'b00000000111000111000001110110011;
ROM[38317] <= 32'b00000000011100010010000000100011;
ROM[38318] <= 32'b00000000010000010000000100010011;
ROM[38319] <= 32'b00000000001100010010000000100011;
ROM[38320] <= 32'b00000000010000010000000100010011;
ROM[38321] <= 32'b00000000010000010010000000100011;
ROM[38322] <= 32'b00000000010000010000000100010011;
ROM[38323] <= 32'b00000000010100010010000000100011;
ROM[38324] <= 32'b00000000010000010000000100010011;
ROM[38325] <= 32'b00000000011000010010000000100011;
ROM[38326] <= 32'b00000000010000010000000100010011;
ROM[38327] <= 32'b00000001010000000000001110010011;
ROM[38328] <= 32'b00000000010000111000001110010011;
ROM[38329] <= 32'b01000000011100010000001110110011;
ROM[38330] <= 32'b00000000011100000000001000110011;
ROM[38331] <= 32'b00000000001000000000000110110011;
ROM[38332] <= 32'b10010110000111111000000011101111;
ROM[38333] <= 32'b11111111110000010000000100010011;
ROM[38334] <= 32'b00000000000000010010001110000011;
ROM[38335] <= 32'b00000000011101100010000000100011;
ROM[38336] <= 32'b00000000110100101000010000110011;
ROM[38337] <= 32'b00000000110001000010001110000011;
ROM[38338] <= 32'b00000000011100010010000000100011;
ROM[38339] <= 32'b00000000010000010000000100010011;
ROM[38340] <= 32'b00000000010000000000001110010011;
ROM[38341] <= 32'b00000000011100010010000000100011;
ROM[38342] <= 32'b00000000010000010000000100010011;
ROM[38343] <= 32'b00000000000000100101001110110111;
ROM[38344] <= 32'b01110110100000111000001110010011;
ROM[38345] <= 32'b00000000111000111000001110110011;
ROM[38346] <= 32'b00000000011100010010000000100011;
ROM[38347] <= 32'b00000000010000010000000100010011;
ROM[38348] <= 32'b00000000001100010010000000100011;
ROM[38349] <= 32'b00000000010000010000000100010011;
ROM[38350] <= 32'b00000000010000010010000000100011;
ROM[38351] <= 32'b00000000010000010000000100010011;
ROM[38352] <= 32'b00000000010100010010000000100011;
ROM[38353] <= 32'b00000000010000010000000100010011;
ROM[38354] <= 32'b00000000011000010010000000100011;
ROM[38355] <= 32'b00000000010000010000000100010011;
ROM[38356] <= 32'b00000001010000000000001110010011;
ROM[38357] <= 32'b00000000100000111000001110010011;
ROM[38358] <= 32'b01000000011100010000001110110011;
ROM[38359] <= 32'b00000000011100000000001000110011;
ROM[38360] <= 32'b00000000001000000000000110110011;
ROM[38361] <= 32'b10001100100011101100000011101111;
ROM[38362] <= 32'b00000000001000000000001110010011;
ROM[38363] <= 32'b00000000011100010010000000100011;
ROM[38364] <= 32'b00000000010000010000000100010011;
ROM[38365] <= 32'b11111111110000010000000100010011;
ROM[38366] <= 32'b00000000000000010010001110000011;
ROM[38367] <= 32'b11111111110000010000000100010011;
ROM[38368] <= 32'b00000000000000010010010000000011;
ROM[38369] <= 32'b00000000011101000000001110110011;
ROM[38370] <= 32'b00000000011100010010000000100011;
ROM[38371] <= 32'b00000000010000010000000100010011;
ROM[38372] <= 32'b00000000110100101000010000110011;
ROM[38373] <= 32'b00000001000001000010001110000011;
ROM[38374] <= 32'b00000000011100010010000000100011;
ROM[38375] <= 32'b00000000010000010000000100010011;
ROM[38376] <= 32'b00000000010000000000001110010011;
ROM[38377] <= 32'b00000000011100010010000000100011;
ROM[38378] <= 32'b00000000010000010000000100010011;
ROM[38379] <= 32'b00000000000000100101001110110111;
ROM[38380] <= 32'b01111111100000111000001110010011;
ROM[38381] <= 32'b00000000111000111000001110110011;
ROM[38382] <= 32'b00000000011100010010000000100011;
ROM[38383] <= 32'b00000000010000010000000100010011;
ROM[38384] <= 32'b00000000001100010010000000100011;
ROM[38385] <= 32'b00000000010000010000000100010011;
ROM[38386] <= 32'b00000000010000010010000000100011;
ROM[38387] <= 32'b00000000010000010000000100010011;
ROM[38388] <= 32'b00000000010100010010000000100011;
ROM[38389] <= 32'b00000000010000010000000100010011;
ROM[38390] <= 32'b00000000011000010010000000100011;
ROM[38391] <= 32'b00000000010000010000000100010011;
ROM[38392] <= 32'b00000001010000000000001110010011;
ROM[38393] <= 32'b00000000100000111000001110010011;
ROM[38394] <= 32'b01000000011100010000001110110011;
ROM[38395] <= 32'b00000000011100000000001000110011;
ROM[38396] <= 32'b00000000001000000000000110110011;
ROM[38397] <= 32'b10000011100011101100000011101111;
ROM[38398] <= 32'b00000000001000000000001110010011;
ROM[38399] <= 32'b00000000011100010010000000100011;
ROM[38400] <= 32'b00000000010000010000000100010011;
ROM[38401] <= 32'b11111111110000010000000100010011;
ROM[38402] <= 32'b00000000000000010010001110000011;
ROM[38403] <= 32'b11111111110000010000000100010011;
ROM[38404] <= 32'b00000000000000010010010000000011;
ROM[38405] <= 32'b00000000011101000000001110110011;
ROM[38406] <= 32'b00000000011100010010000000100011;
ROM[38407] <= 32'b00000000010000010000000100010011;
ROM[38408] <= 32'b00000000001000000000001110010011;
ROM[38409] <= 32'b00000000011100010010000000100011;
ROM[38410] <= 32'b00000000010000010000000100010011;
ROM[38411] <= 32'b00000000000000100110001110110111;
ROM[38412] <= 32'b10000111100000111000001110010011;
ROM[38413] <= 32'b00000000111000111000001110110011;
ROM[38414] <= 32'b00000000011100010010000000100011;
ROM[38415] <= 32'b00000000010000010000000100010011;
ROM[38416] <= 32'b00000000001100010010000000100011;
ROM[38417] <= 32'b00000000010000010000000100010011;
ROM[38418] <= 32'b00000000010000010010000000100011;
ROM[38419] <= 32'b00000000010000010000000100010011;
ROM[38420] <= 32'b00000000010100010010000000100011;
ROM[38421] <= 32'b00000000010000010000000100010011;
ROM[38422] <= 32'b00000000011000010010000000100011;
ROM[38423] <= 32'b00000000010000010000000100010011;
ROM[38424] <= 32'b00000001010000000000001110010011;
ROM[38425] <= 32'b00000000110000111000001110010011;
ROM[38426] <= 32'b01000000011100010000001110110011;
ROM[38427] <= 32'b00000000011100000000001000110011;
ROM[38428] <= 32'b00000000001000000000000110110011;
ROM[38429] <= 32'b11001111010111111001000011101111;
ROM[38430] <= 32'b11111111110000010000000100010011;
ROM[38431] <= 32'b00000000000000010010001110000011;
ROM[38432] <= 32'b00000000011101100010000000100011;
ROM[38433] <= 32'b00000000000000000000001110010011;
ROM[38434] <= 32'b00000000011100010010000000100011;
ROM[38435] <= 32'b00000000010000010000000100010011;
ROM[38436] <= 32'b00000001010000000000001110010011;
ROM[38437] <= 32'b01000000011100011000001110110011;
ROM[38438] <= 32'b00000000000000111010000010000011;
ROM[38439] <= 32'b11111111110000010000000100010011;
ROM[38440] <= 32'b00000000000000010010001110000011;
ROM[38441] <= 32'b00000000011100100010000000100011;
ROM[38442] <= 32'b00000000010000100000000100010011;
ROM[38443] <= 32'b00000001010000000000001110010011;
ROM[38444] <= 32'b01000000011100011000001110110011;
ROM[38445] <= 32'b00000000010000111010000110000011;
ROM[38446] <= 32'b00000000100000111010001000000011;
ROM[38447] <= 32'b00000000110000111010001010000011;
ROM[38448] <= 32'b00000001000000111010001100000011;
ROM[38449] <= 32'b00000000000000001000000011100111;
ROM[38450] <= 32'b00000000000000010010000000100011;
ROM[38451] <= 32'b00000000010000010000000100010011;
ROM[38452] <= 32'b00000000000000010010000000100011;
ROM[38453] <= 32'b00000000010000010000000100010011;
ROM[38454] <= 32'b00000000000000010010000000100011;
ROM[38455] <= 32'b00000000010000010000000100010011;
ROM[38456] <= 32'b00000000000000100010001110000011;
ROM[38457] <= 32'b00000000011100010010000000100011;
ROM[38458] <= 32'b00000000010000010000000100010011;
ROM[38459] <= 32'b11111111110000010000000100010011;
ROM[38460] <= 32'b00000000000000010010001110000011;
ROM[38461] <= 32'b00000000000000111000001010010011;
ROM[38462] <= 32'b00000000110100101000010000110011;
ROM[38463] <= 32'b00000000010001000010001110000011;
ROM[38464] <= 32'b00000000011100010010000000100011;
ROM[38465] <= 32'b00000000010000010000000100010011;
ROM[38466] <= 32'b00000000000000100110001110110111;
ROM[38467] <= 32'b10010101010000111000001110010011;
ROM[38468] <= 32'b00000000111000111000001110110011;
ROM[38469] <= 32'b00000000011100010010000000100011;
ROM[38470] <= 32'b00000000010000010000000100010011;
ROM[38471] <= 32'b00000000001100010010000000100011;
ROM[38472] <= 32'b00000000010000010000000100010011;
ROM[38473] <= 32'b00000000010000010010000000100011;
ROM[38474] <= 32'b00000000010000010000000100010011;
ROM[38475] <= 32'b00000000010100010010000000100011;
ROM[38476] <= 32'b00000000010000010000000100010011;
ROM[38477] <= 32'b00000000011000010010000000100011;
ROM[38478] <= 32'b00000000010000010000000100010011;
ROM[38479] <= 32'b00000001010000000000001110010011;
ROM[38480] <= 32'b00000000010000111000001110010011;
ROM[38481] <= 32'b01000000011100010000001110110011;
ROM[38482] <= 32'b00000000011100000000001000110011;
ROM[38483] <= 32'b00000000001000000000000110110011;
ROM[38484] <= 32'b11110011000011011010000011101111;
ROM[38485] <= 32'b11111111110000010000000100010011;
ROM[38486] <= 32'b00000000000000010010001110000011;
ROM[38487] <= 32'b00000000110100101000010000110011;
ROM[38488] <= 32'b00000000011101000010101000100011;
ROM[38489] <= 32'b00000000000000000000001110010011;
ROM[38490] <= 32'b00000000011100010010000000100011;
ROM[38491] <= 32'b00000000010000010000000100010011;
ROM[38492] <= 32'b11111111110000010000000100010011;
ROM[38493] <= 32'b00000000000000010010001110000011;
ROM[38494] <= 32'b00000000011100011010000000100011;
ROM[38495] <= 32'b00000000000000011010001110000011;
ROM[38496] <= 32'b00000000011100010010000000100011;
ROM[38497] <= 32'b00000000010000010000000100010011;
ROM[38498] <= 32'b00000000110100101000010000110011;
ROM[38499] <= 32'b00000000010001000010001110000011;
ROM[38500] <= 32'b00000000011100010010000000100011;
ROM[38501] <= 32'b00000000010000010000000100010011;
ROM[38502] <= 32'b11111111110000010000000100010011;
ROM[38503] <= 32'b00000000000000010010001110000011;
ROM[38504] <= 32'b11111111110000010000000100010011;
ROM[38505] <= 32'b00000000000000010010010000000011;
ROM[38506] <= 32'b00000000011101000010001110110011;
ROM[38507] <= 32'b00000000011100010010000000100011;
ROM[38508] <= 32'b00000000010000010000000100010011;
ROM[38509] <= 32'b11111111110000010000000100010011;
ROM[38510] <= 32'b00000000000000010010001110000011;
ROM[38511] <= 32'b01000000011100000000001110110011;
ROM[38512] <= 32'b00000000000100111000001110010011;
ROM[38513] <= 32'b00000000011100010010000000100011;
ROM[38514] <= 32'b00000000010000010000000100010011;
ROM[38515] <= 32'b11111111110000010000000100010011;
ROM[38516] <= 32'b00000000000000010010001110000011;
ROM[38517] <= 32'b00000000000000111000101001100011;
ROM[38518] <= 32'b00000000000000100110001110110111;
ROM[38519] <= 32'b11001100100000111000001110010011;
ROM[38520] <= 32'b00000000111000111000001110110011;
ROM[38521] <= 32'b00000000000000111000000011100111;
ROM[38522] <= 32'b00000000110100101000010000110011;
ROM[38523] <= 32'b00000000100001000010001110000011;
ROM[38524] <= 32'b00000000011100010010000000100011;
ROM[38525] <= 32'b00000000010000010000000100010011;
ROM[38526] <= 32'b00000000000000100110001110110111;
ROM[38527] <= 32'b10100100010000111000001110010011;
ROM[38528] <= 32'b00000000111000111000001110110011;
ROM[38529] <= 32'b00000000011100010010000000100011;
ROM[38530] <= 32'b00000000010000010000000100010011;
ROM[38531] <= 32'b00000000001100010010000000100011;
ROM[38532] <= 32'b00000000010000010000000100010011;
ROM[38533] <= 32'b00000000010000010010000000100011;
ROM[38534] <= 32'b00000000010000010000000100010011;
ROM[38535] <= 32'b00000000010100010010000000100011;
ROM[38536] <= 32'b00000000010000010000000100010011;
ROM[38537] <= 32'b00000000011000010010000000100011;
ROM[38538] <= 32'b00000000010000010000000100010011;
ROM[38539] <= 32'b00000001010000000000001110010011;
ROM[38540] <= 32'b00000000010000111000001110010011;
ROM[38541] <= 32'b01000000011100010000001110110011;
ROM[38542] <= 32'b00000000011100000000001000110011;
ROM[38543] <= 32'b00000000001000000000000110110011;
ROM[38544] <= 32'b11100100000011011010000011101111;
ROM[38545] <= 32'b11111111110000010000000100010011;
ROM[38546] <= 32'b00000000000000010010001110000011;
ROM[38547] <= 32'b00000000011100011010010000100011;
ROM[38548] <= 32'b00000000000000000000001110010011;
ROM[38549] <= 32'b00000000011100010010000000100011;
ROM[38550] <= 32'b00000000010000010000000100010011;
ROM[38551] <= 32'b11111111110000010000000100010011;
ROM[38552] <= 32'b00000000000000010010001110000011;
ROM[38553] <= 32'b00000000011100011010001000100011;
ROM[38554] <= 32'b00000000010000011010001110000011;
ROM[38555] <= 32'b00000000011100010010000000100011;
ROM[38556] <= 32'b00000000010000010000000100010011;
ROM[38557] <= 32'b00000000110100101000010000110011;
ROM[38558] <= 32'b00000000100001000010001110000011;
ROM[38559] <= 32'b00000000011100010010000000100011;
ROM[38560] <= 32'b00000000010000010000000100010011;
ROM[38561] <= 32'b11111111110000010000000100010011;
ROM[38562] <= 32'b00000000000000010010001110000011;
ROM[38563] <= 32'b11111111110000010000000100010011;
ROM[38564] <= 32'b00000000000000010010010000000011;
ROM[38565] <= 32'b00000000011101000010001110110011;
ROM[38566] <= 32'b00000000011100010010000000100011;
ROM[38567] <= 32'b00000000010000010000000100010011;
ROM[38568] <= 32'b11111111110000010000000100010011;
ROM[38569] <= 32'b00000000000000010010001110000011;
ROM[38570] <= 32'b01000000011100000000001110110011;
ROM[38571] <= 32'b00000000000100111000001110010011;
ROM[38572] <= 32'b00000000011100010010000000100011;
ROM[38573] <= 32'b00000000010000010000000100010011;
ROM[38574] <= 32'b11111111110000010000000100010011;
ROM[38575] <= 32'b00000000000000010010001110000011;
ROM[38576] <= 32'b00000000000000111000101001100011;
ROM[38577] <= 32'b00000000000000100110001110110111;
ROM[38578] <= 32'b10111100110000111000001110010011;
ROM[38579] <= 32'b00000000111000111000001110110011;
ROM[38580] <= 32'b00000000000000111000000011100111;
ROM[38581] <= 32'b00000000000000000000001110010011;
ROM[38582] <= 32'b00000000011100010010000000100011;
ROM[38583] <= 32'b00000000010000010000000100010011;
ROM[38584] <= 32'b00000000100000011010001110000011;
ROM[38585] <= 32'b00000000011100010010000000100011;
ROM[38586] <= 32'b00000000010000010000000100010011;
ROM[38587] <= 32'b00000000010000011010001110000011;
ROM[38588] <= 32'b00000000011100010010000000100011;
ROM[38589] <= 32'b00000000010000010000000100010011;
ROM[38590] <= 32'b00000000010000000000001110010011;
ROM[38591] <= 32'b00000000011100010010000000100011;
ROM[38592] <= 32'b00000000010000010000000100010011;
ROM[38593] <= 32'b00000000000000100110001110110111;
ROM[38594] <= 32'b10110101000000111000001110010011;
ROM[38595] <= 32'b00000000111000111000001110110011;
ROM[38596] <= 32'b00000000011100010010000000100011;
ROM[38597] <= 32'b00000000010000010000000100010011;
ROM[38598] <= 32'b00000000001100010010000000100011;
ROM[38599] <= 32'b00000000010000010000000100010011;
ROM[38600] <= 32'b00000000010000010010000000100011;
ROM[38601] <= 32'b00000000010000010000000100010011;
ROM[38602] <= 32'b00000000010100010010000000100011;
ROM[38603] <= 32'b00000000010000010000000100010011;
ROM[38604] <= 32'b00000000011000010010000000100011;
ROM[38605] <= 32'b00000000010000010000000100010011;
ROM[38606] <= 32'b00000001010000000000001110010011;
ROM[38607] <= 32'b00000000100000111000001110010011;
ROM[38608] <= 32'b01000000011100010000001110110011;
ROM[38609] <= 32'b00000000011100000000001000110011;
ROM[38610] <= 32'b00000000001000000000000110110011;
ROM[38611] <= 32'b11001110000111101011000011101111;
ROM[38612] <= 32'b11111111110000010000000100010011;
ROM[38613] <= 32'b00000000000000010010001110000011;
ROM[38614] <= 32'b11111111110000010000000100010011;
ROM[38615] <= 32'b00000000000000010010010000000011;
ROM[38616] <= 32'b00000000011101000000001110110011;
ROM[38617] <= 32'b00000000011100010010000000100011;
ROM[38618] <= 32'b00000000010000010000000100010011;
ROM[38619] <= 32'b11111111110000010000000100010011;
ROM[38620] <= 32'b00000000000000010010001110000011;
ROM[38621] <= 32'b00000000000000111000001100010011;
ROM[38622] <= 32'b11111111110000010000000100010011;
ROM[38623] <= 32'b00000000000000010010001110000011;
ROM[38624] <= 32'b00000000110100110000010000110011;
ROM[38625] <= 32'b00000000011101000010000000100011;
ROM[38626] <= 32'b00000000010000011010001110000011;
ROM[38627] <= 32'b00000000011100010010000000100011;
ROM[38628] <= 32'b00000000010000010000000100010011;
ROM[38629] <= 32'b00000000000100000000001110010011;
ROM[38630] <= 32'b00000000011100010010000000100011;
ROM[38631] <= 32'b00000000010000010000000100010011;
ROM[38632] <= 32'b11111111110000010000000100010011;
ROM[38633] <= 32'b00000000000000010010001110000011;
ROM[38634] <= 32'b11111111110000010000000100010011;
ROM[38635] <= 32'b00000000000000010010010000000011;
ROM[38636] <= 32'b00000000011101000000001110110011;
ROM[38637] <= 32'b00000000011100010010000000100011;
ROM[38638] <= 32'b00000000010000010000000100010011;
ROM[38639] <= 32'b11111111110000010000000100010011;
ROM[38640] <= 32'b00000000000000010010001110000011;
ROM[38641] <= 32'b00000000011100011010001000100011;
ROM[38642] <= 32'b11101010000111111111000011101111;
ROM[38643] <= 32'b00000000100000011010001110000011;
ROM[38644] <= 32'b00000000011100010010000000100011;
ROM[38645] <= 32'b00000000010000010000000100010011;
ROM[38646] <= 32'b00000000110100101000010000110011;
ROM[38647] <= 32'b00000001010001000010001110000011;
ROM[38648] <= 32'b00000000011100010010000000100011;
ROM[38649] <= 32'b00000000010000010000000100010011;
ROM[38650] <= 32'b00000000000000011010001110000011;
ROM[38651] <= 32'b00000000011100010010000000100011;
ROM[38652] <= 32'b00000000010000010000000100010011;
ROM[38653] <= 32'b00000000010000000000001110010011;
ROM[38654] <= 32'b00000000011100010010000000100011;
ROM[38655] <= 32'b00000000010000010000000100010011;
ROM[38656] <= 32'b00000000000000100110001110110111;
ROM[38657] <= 32'b11000100110000111000001110010011;
ROM[38658] <= 32'b00000000111000111000001110110011;
ROM[38659] <= 32'b00000000011100010010000000100011;
ROM[38660] <= 32'b00000000010000010000000100010011;
ROM[38661] <= 32'b00000000001100010010000000100011;
ROM[38662] <= 32'b00000000010000010000000100010011;
ROM[38663] <= 32'b00000000010000010010000000100011;
ROM[38664] <= 32'b00000000010000010000000100010011;
ROM[38665] <= 32'b00000000010100010010000000100011;
ROM[38666] <= 32'b00000000010000010000000100010011;
ROM[38667] <= 32'b00000000011000010010000000100011;
ROM[38668] <= 32'b00000000010000010000000100010011;
ROM[38669] <= 32'b00000001010000000000001110010011;
ROM[38670] <= 32'b00000000100000111000001110010011;
ROM[38671] <= 32'b01000000011100010000001110110011;
ROM[38672] <= 32'b00000000011100000000001000110011;
ROM[38673] <= 32'b00000000001000000000000110110011;
ROM[38674] <= 32'b10111110010111101011000011101111;
ROM[38675] <= 32'b11111111110000010000000100010011;
ROM[38676] <= 32'b00000000000000010010001110000011;
ROM[38677] <= 32'b11111111110000010000000100010011;
ROM[38678] <= 32'b00000000000000010010010000000011;
ROM[38679] <= 32'b00000000011101000000001110110011;
ROM[38680] <= 32'b00000000011100010010000000100011;
ROM[38681] <= 32'b00000000010000010000000100010011;
ROM[38682] <= 32'b11111111110000010000000100010011;
ROM[38683] <= 32'b00000000000000010010001110000011;
ROM[38684] <= 32'b00000000000000111000001100010011;
ROM[38685] <= 32'b11111111110000010000000100010011;
ROM[38686] <= 32'b00000000000000010010001110000011;
ROM[38687] <= 32'b00000000110100110000010000110011;
ROM[38688] <= 32'b00000000011101000010000000100011;
ROM[38689] <= 32'b00000000000000011010001110000011;
ROM[38690] <= 32'b00000000011100010010000000100011;
ROM[38691] <= 32'b00000000010000010000000100010011;
ROM[38692] <= 32'b00000000000100000000001110010011;
ROM[38693] <= 32'b00000000011100010010000000100011;
ROM[38694] <= 32'b00000000010000010000000100010011;
ROM[38695] <= 32'b11111111110000010000000100010011;
ROM[38696] <= 32'b00000000000000010010001110000011;
ROM[38697] <= 32'b11111111110000010000000100010011;
ROM[38698] <= 32'b00000000000000010010010000000011;
ROM[38699] <= 32'b00000000011101000000001110110011;
ROM[38700] <= 32'b00000000011100010010000000100011;
ROM[38701] <= 32'b00000000010000010000000100010011;
ROM[38702] <= 32'b11111111110000010000000100010011;
ROM[38703] <= 32'b00000000000000010010001110000011;
ROM[38704] <= 32'b00000000011100011010000000100011;
ROM[38705] <= 32'b11001011100111111111000011101111;
ROM[38706] <= 32'b00000000000100000000001110010011;
ROM[38707] <= 32'b00000000011100010010000000100011;
ROM[38708] <= 32'b00000000010000010000000100010011;
ROM[38709] <= 32'b11111111110000010000000100010011;
ROM[38710] <= 32'b00000000000000010010001110000011;
ROM[38711] <= 32'b01000000011100000000001110110011;
ROM[38712] <= 32'b00000000011100010010000000100011;
ROM[38713] <= 32'b00000000010000010000000100010011;
ROM[38714] <= 32'b00000000000000100110001110110111;
ROM[38715] <= 32'b11010011010000111000001110010011;
ROM[38716] <= 32'b00000000111000111000001110110011;
ROM[38717] <= 32'b00000000011100010010000000100011;
ROM[38718] <= 32'b00000000010000010000000100010011;
ROM[38719] <= 32'b00000000001100010010000000100011;
ROM[38720] <= 32'b00000000010000010000000100010011;
ROM[38721] <= 32'b00000000010000010010000000100011;
ROM[38722] <= 32'b00000000010000010000000100010011;
ROM[38723] <= 32'b00000000010100010010000000100011;
ROM[38724] <= 32'b00000000010000010000000100010011;
ROM[38725] <= 32'b00000000011000010010000000100011;
ROM[38726] <= 32'b00000000010000010000000100010011;
ROM[38727] <= 32'b00000001010000000000001110010011;
ROM[38728] <= 32'b00000000010000111000001110010011;
ROM[38729] <= 32'b01000000011100010000001110110011;
ROM[38730] <= 32'b00000000011100000000001000110011;
ROM[38731] <= 32'b00000000001000000000000110110011;
ROM[38732] <= 32'b10110010000011111000000011101111;
ROM[38733] <= 32'b11111111110000010000000100010011;
ROM[38734] <= 32'b00000000000000010010001110000011;
ROM[38735] <= 32'b00000000011101100010000000100011;
ROM[38736] <= 32'b00000000000000000000001110010011;
ROM[38737] <= 32'b00000000011100010010000000100011;
ROM[38738] <= 32'b00000000010000010000000100010011;
ROM[38739] <= 32'b00000000110100101000010000110011;
ROM[38740] <= 32'b00000000100001000010001110000011;
ROM[38741] <= 32'b00000000011100010010000000100011;
ROM[38742] <= 32'b00000000010000010000000100010011;
ROM[38743] <= 32'b00000000010000000000001110010011;
ROM[38744] <= 32'b00000000011100010010000000100011;
ROM[38745] <= 32'b00000000010000010000000100010011;
ROM[38746] <= 32'b00000000000000100110001110110111;
ROM[38747] <= 32'b11011011010000111000001110010011;
ROM[38748] <= 32'b00000000111000111000001110110011;
ROM[38749] <= 32'b00000000011100010010000000100011;
ROM[38750] <= 32'b00000000010000010000000100010011;
ROM[38751] <= 32'b00000000001100010010000000100011;
ROM[38752] <= 32'b00000000010000010000000100010011;
ROM[38753] <= 32'b00000000010000010010000000100011;
ROM[38754] <= 32'b00000000010000010000000100010011;
ROM[38755] <= 32'b00000000010100010010000000100011;
ROM[38756] <= 32'b00000000010000010000000100010011;
ROM[38757] <= 32'b00000000011000010010000000100011;
ROM[38758] <= 32'b00000000010000010000000100010011;
ROM[38759] <= 32'b00000001010000000000001110010011;
ROM[38760] <= 32'b00000000100000111000001110010011;
ROM[38761] <= 32'b01000000011100010000001110110011;
ROM[38762] <= 32'b00000000011100000000001000110011;
ROM[38763] <= 32'b00000000001000000000000110110011;
ROM[38764] <= 32'b10100111110111101011000011101111;
ROM[38765] <= 32'b00000000000100000000001110010011;
ROM[38766] <= 32'b00000000011100010010000000100011;
ROM[38767] <= 32'b00000000010000010000000100010011;
ROM[38768] <= 32'b11111111110000010000000100010011;
ROM[38769] <= 32'b00000000000000010010001110000011;
ROM[38770] <= 32'b11111111110000010000000100010011;
ROM[38771] <= 32'b00000000000000010010010000000011;
ROM[38772] <= 32'b00000000011101000000001110110011;
ROM[38773] <= 32'b00000000011100010010000000100011;
ROM[38774] <= 32'b00000000010000010000000100010011;
ROM[38775] <= 32'b00000000110100101000010000110011;
ROM[38776] <= 32'b00000000010001000010001110000011;
ROM[38777] <= 32'b00000000011100010010000000100011;
ROM[38778] <= 32'b00000000010000010000000100010011;
ROM[38779] <= 32'b00000000010000000000001110010011;
ROM[38780] <= 32'b00000000011100010010000000100011;
ROM[38781] <= 32'b00000000010000010000000100010011;
ROM[38782] <= 32'b00000000000000100110001110110111;
ROM[38783] <= 32'b11100100010000111000001110010011;
ROM[38784] <= 32'b00000000111000111000001110110011;
ROM[38785] <= 32'b00000000011100010010000000100011;
ROM[38786] <= 32'b00000000010000010000000100010011;
ROM[38787] <= 32'b00000000001100010010000000100011;
ROM[38788] <= 32'b00000000010000010000000100010011;
ROM[38789] <= 32'b00000000010000010010000000100011;
ROM[38790] <= 32'b00000000010000010000000100010011;
ROM[38791] <= 32'b00000000010100010010000000100011;
ROM[38792] <= 32'b00000000010000010000000100010011;
ROM[38793] <= 32'b00000000011000010010000000100011;
ROM[38794] <= 32'b00000000010000010000000100010011;
ROM[38795] <= 32'b00000001010000000000001110010011;
ROM[38796] <= 32'b00000000100000111000001110010011;
ROM[38797] <= 32'b01000000011100010000001110110011;
ROM[38798] <= 32'b00000000011100000000001000110011;
ROM[38799] <= 32'b00000000001000000000000110110011;
ROM[38800] <= 32'b10011110110111101011000011101111;
ROM[38801] <= 32'b00000000000100000000001110010011;
ROM[38802] <= 32'b00000000011100010010000000100011;
ROM[38803] <= 32'b00000000010000010000000100010011;
ROM[38804] <= 32'b11111111110000010000000100010011;
ROM[38805] <= 32'b00000000000000010010001110000011;
ROM[38806] <= 32'b11111111110000010000000100010011;
ROM[38807] <= 32'b00000000000000010010010000000011;
ROM[38808] <= 32'b01000000011101000000001110110011;
ROM[38809] <= 32'b00000000011100010010000000100011;
ROM[38810] <= 32'b00000000010000010000000100010011;
ROM[38811] <= 32'b00000000110100101000010000110011;
ROM[38812] <= 32'b00000000100001000010001110000011;
ROM[38813] <= 32'b00000000011100010010000000100011;
ROM[38814] <= 32'b00000000010000010000000100010011;
ROM[38815] <= 32'b00000000010000000000001110010011;
ROM[38816] <= 32'b00000000011100010010000000100011;
ROM[38817] <= 32'b00000000010000010000000100010011;
ROM[38818] <= 32'b00000000000000100110001110110111;
ROM[38819] <= 32'b11101101010000111000001110010011;
ROM[38820] <= 32'b00000000111000111000001110110011;
ROM[38821] <= 32'b00000000011100010010000000100011;
ROM[38822] <= 32'b00000000010000010000000100010011;
ROM[38823] <= 32'b00000000001100010010000000100011;
ROM[38824] <= 32'b00000000010000010000000100010011;
ROM[38825] <= 32'b00000000010000010010000000100011;
ROM[38826] <= 32'b00000000010000010000000100010011;
ROM[38827] <= 32'b00000000010100010010000000100011;
ROM[38828] <= 32'b00000000010000010000000100010011;
ROM[38829] <= 32'b00000000011000010010000000100011;
ROM[38830] <= 32'b00000000010000010000000100010011;
ROM[38831] <= 32'b00000001010000000000001110010011;
ROM[38832] <= 32'b00000000100000111000001110010011;
ROM[38833] <= 32'b01000000011100010000001110110011;
ROM[38834] <= 32'b00000000011100000000001000110011;
ROM[38835] <= 32'b00000000001000000000000110110011;
ROM[38836] <= 32'b10010101110111101011000011101111;
ROM[38837] <= 32'b00000000000100000000001110010011;
ROM[38838] <= 32'b00000000011100010010000000100011;
ROM[38839] <= 32'b00000000010000010000000100010011;
ROM[38840] <= 32'b11111111110000010000000100010011;
ROM[38841] <= 32'b00000000000000010010001110000011;
ROM[38842] <= 32'b11111111110000010000000100010011;
ROM[38843] <= 32'b00000000000000010010010000000011;
ROM[38844] <= 32'b00000000011101000000001110110011;
ROM[38845] <= 32'b00000000011100010010000000100011;
ROM[38846] <= 32'b00000000010000010000000100010011;
ROM[38847] <= 32'b00000000000000100110001110110111;
ROM[38848] <= 32'b11110100100000111000001110010011;
ROM[38849] <= 32'b00000000111000111000001110110011;
ROM[38850] <= 32'b00000000011100010010000000100011;
ROM[38851] <= 32'b00000000010000010000000100010011;
ROM[38852] <= 32'b00000000001100010010000000100011;
ROM[38853] <= 32'b00000000010000010000000100010011;
ROM[38854] <= 32'b00000000010000010010000000100011;
ROM[38855] <= 32'b00000000010000010000000100010011;
ROM[38856] <= 32'b00000000010100010010000000100011;
ROM[38857] <= 32'b00000000010000010000000100010011;
ROM[38858] <= 32'b00000000011000010010000000100011;
ROM[38859] <= 32'b00000000010000010000000100010011;
ROM[38860] <= 32'b00000001010000000000001110010011;
ROM[38861] <= 32'b00000001000000111000001110010011;
ROM[38862] <= 32'b01000000011100010000001110110011;
ROM[38863] <= 32'b00000000011100000000001000110011;
ROM[38864] <= 32'b00000000001000000000000110110011;
ROM[38865] <= 32'b11100000010011111000000011101111;
ROM[38866] <= 32'b11111111110000010000000100010011;
ROM[38867] <= 32'b00000000000000010010001110000011;
ROM[38868] <= 32'b00000000011101100010000000100011;
ROM[38869] <= 32'b00000000000000000000001110010011;
ROM[38870] <= 32'b00000000011100010010000000100011;
ROM[38871] <= 32'b00000000010000010000000100010011;
ROM[38872] <= 32'b00000001010000000000001110010011;
ROM[38873] <= 32'b01000000011100011000001110110011;
ROM[38874] <= 32'b00000000000000111010000010000011;
ROM[38875] <= 32'b11111111110000010000000100010011;
ROM[38876] <= 32'b00000000000000010010001110000011;
ROM[38877] <= 32'b00000000011100100010000000100011;
ROM[38878] <= 32'b00000000010000100000000100010011;
ROM[38879] <= 32'b00000001010000000000001110010011;
ROM[38880] <= 32'b01000000011100011000001110110011;
ROM[38881] <= 32'b00000000010000111010000110000011;
ROM[38882] <= 32'b00000000100000111010001000000011;
ROM[38883] <= 32'b00000000110000111010001010000011;
ROM[38884] <= 32'b00000001000000111010001100000011;
ROM[38885] <= 32'b00000000000000001000000011100111;
ROM[38886] <= 32'b00000000000000100010001110000011;
ROM[38887] <= 32'b00000000011100010010000000100011;
ROM[38888] <= 32'b00000000010000010000000100010011;
ROM[38889] <= 32'b11111111110000010000000100010011;
ROM[38890] <= 32'b00000000000000010010001110000011;
ROM[38891] <= 32'b00000000000000111000001010010011;
ROM[38892] <= 32'b00000000110100101000010000110011;
ROM[38893] <= 32'b00000000010001000010001110000011;
ROM[38894] <= 32'b00000000011100010010000000100011;
ROM[38895] <= 32'b00000000010000010000000100010011;
ROM[38896] <= 32'b00000001010000000000001110010011;
ROM[38897] <= 32'b01000000011100011000001110110011;
ROM[38898] <= 32'b00000000000000111010000010000011;
ROM[38899] <= 32'b11111111110000010000000100010011;
ROM[38900] <= 32'b00000000000000010010001110000011;
ROM[38901] <= 32'b00000000011100100010000000100011;
ROM[38902] <= 32'b00000000010000100000000100010011;
ROM[38903] <= 32'b00000001010000000000001110010011;
ROM[38904] <= 32'b01000000011100011000001110110011;
ROM[38905] <= 32'b00000000010000111010000110000011;
ROM[38906] <= 32'b00000000100000111010001000000011;
ROM[38907] <= 32'b00000000110000111010001010000011;
ROM[38908] <= 32'b00000001000000111010001100000011;
ROM[38909] <= 32'b00000000000000001000000011100111;
ROM[38910] <= 32'b00000000000000100010001110000011;
ROM[38911] <= 32'b00000000011100010010000000100011;
ROM[38912] <= 32'b00000000010000010000000100010011;
ROM[38913] <= 32'b11111111110000010000000100010011;
ROM[38914] <= 32'b00000000000000010010001110000011;
ROM[38915] <= 32'b00000000000000111000001010010011;
ROM[38916] <= 32'b00000000110100101000010000110011;
ROM[38917] <= 32'b00000000100001000010001110000011;
ROM[38918] <= 32'b00000000011100010010000000100011;
ROM[38919] <= 32'b00000000010000010000000100010011;
ROM[38920] <= 32'b00000001010000000000001110010011;
ROM[38921] <= 32'b01000000011100011000001110110011;
ROM[38922] <= 32'b00000000000000111010000010000011;
ROM[38923] <= 32'b11111111110000010000000100010011;
ROM[38924] <= 32'b00000000000000010010001110000011;
ROM[38925] <= 32'b00000000011100100010000000100011;
ROM[38926] <= 32'b00000000010000100000000100010011;
ROM[38927] <= 32'b00000001010000000000001110010011;
ROM[38928] <= 32'b01000000011100011000001110110011;
ROM[38929] <= 32'b00000000010000111010000110000011;
ROM[38930] <= 32'b00000000100000111010001000000011;
ROM[38931] <= 32'b00000000110000111010001010000011;
ROM[38932] <= 32'b00000001000000111010001100000011;
ROM[38933] <= 32'b00000000000000001000000011100111;
ROM[38934] <= 32'b00000000000000100010001110000011;
ROM[38935] <= 32'b00000000011100010010000000100011;
ROM[38936] <= 32'b00000000010000010000000100010011;
ROM[38937] <= 32'b11111111110000010000000100010011;
ROM[38938] <= 32'b00000000000000010010001110000011;
ROM[38939] <= 32'b00000000000000111000001010010011;
ROM[38940] <= 32'b00000000110100101000010000110011;
ROM[38941] <= 32'b00000000110001000010001110000011;
ROM[38942] <= 32'b00000000011100010010000000100011;
ROM[38943] <= 32'b00000000010000010000000100010011;
ROM[38944] <= 32'b00000001010000000000001110010011;
ROM[38945] <= 32'b01000000011100011000001110110011;
ROM[38946] <= 32'b00000000000000111010000010000011;
ROM[38947] <= 32'b11111111110000010000000100010011;
ROM[38948] <= 32'b00000000000000010010001110000011;
ROM[38949] <= 32'b00000000011100100010000000100011;
ROM[38950] <= 32'b00000000010000100000000100010011;
ROM[38951] <= 32'b00000001010000000000001110010011;
ROM[38952] <= 32'b01000000011100011000001110110011;
ROM[38953] <= 32'b00000000010000111010000110000011;
ROM[38954] <= 32'b00000000100000111010001000000011;
ROM[38955] <= 32'b00000000110000111010001010000011;
ROM[38956] <= 32'b00000001000000111010001100000011;
ROM[38957] <= 32'b00000000000000001000000011100111;
ROM[38958] <= 32'b00000000000000100010001110000011;
ROM[38959] <= 32'b00000000011100010010000000100011;
ROM[38960] <= 32'b00000000010000010000000100010011;
ROM[38961] <= 32'b11111111110000010000000100010011;
ROM[38962] <= 32'b00000000000000010010001110000011;
ROM[38963] <= 32'b00000000000000111000001010010011;
ROM[38964] <= 32'b00000000110100101000010000110011;
ROM[38965] <= 32'b00000001000001000010001110000011;
ROM[38966] <= 32'b00000000011100010010000000100011;
ROM[38967] <= 32'b00000000010000010000000100010011;
ROM[38968] <= 32'b00000001010000000000001110010011;
ROM[38969] <= 32'b01000000011100011000001110110011;
ROM[38970] <= 32'b00000000000000111010000010000011;
ROM[38971] <= 32'b11111111110000010000000100010011;
ROM[38972] <= 32'b00000000000000010010001110000011;
ROM[38973] <= 32'b00000000011100100010000000100011;
ROM[38974] <= 32'b00000000010000100000000100010011;
ROM[38975] <= 32'b00000001010000000000001110010011;
ROM[38976] <= 32'b01000000011100011000001110110011;
ROM[38977] <= 32'b00000000010000111010000110000011;
ROM[38978] <= 32'b00000000100000111010001000000011;
ROM[38979] <= 32'b00000000110000111010001010000011;
ROM[38980] <= 32'b00000001000000111010001100000011;
ROM[38981] <= 32'b00000000000000001000000011100111;
ROM[38982] <= 32'b00000000000000010010000000100011;
ROM[38983] <= 32'b00000000010000010000000100010011;
ROM[38984] <= 32'b00000000000000100010001110000011;
ROM[38985] <= 32'b00000000011100010010000000100011;
ROM[38986] <= 32'b00000000010000010000000100010011;
ROM[38987] <= 32'b11111111110000010000000100010011;
ROM[38988] <= 32'b00000000000000010010001110000011;
ROM[38989] <= 32'b00000000000000111000001010010011;
ROM[38990] <= 32'b00000000110100101000010000110011;
ROM[38991] <= 32'b00000001010001000010001110000011;
ROM[38992] <= 32'b00000000011100010010000000100011;
ROM[38993] <= 32'b00000000010000010000000100010011;
ROM[38994] <= 32'b00000000010000100010001110000011;
ROM[38995] <= 32'b00000000011100010010000000100011;
ROM[38996] <= 32'b00000000010000010000000100010011;
ROM[38997] <= 32'b00000000010000000000001110010011;
ROM[38998] <= 32'b00000000011100010010000000100011;
ROM[38999] <= 32'b00000000010000010000000100010011;
ROM[39000] <= 32'b00000000000000100110001110110111;
ROM[39001] <= 32'b00011010110000111000001110010011;
ROM[39002] <= 32'b00000000111000111000001110110011;
ROM[39003] <= 32'b00000000011100010010000000100011;
ROM[39004] <= 32'b00000000010000010000000100010011;
ROM[39005] <= 32'b00000000001100010010000000100011;
ROM[39006] <= 32'b00000000010000010000000100010011;
ROM[39007] <= 32'b00000000010000010010000000100011;
ROM[39008] <= 32'b00000000010000010000000100010011;
ROM[39009] <= 32'b00000000010100010010000000100011;
ROM[39010] <= 32'b00000000010000010000000100010011;
ROM[39011] <= 32'b00000000011000010010000000100011;
ROM[39012] <= 32'b00000000010000010000000100010011;
ROM[39013] <= 32'b00000001010000000000001110010011;
ROM[39014] <= 32'b00000000100000111000001110010011;
ROM[39015] <= 32'b01000000011100010000001110110011;
ROM[39016] <= 32'b00000000011100000000001000110011;
ROM[39017] <= 32'b00000000001000000000000110110011;
ROM[39018] <= 32'b11101000010011101011000011101111;
ROM[39019] <= 32'b11111111110000010000000100010011;
ROM[39020] <= 32'b00000000000000010010001110000011;
ROM[39021] <= 32'b11111111110000010000000100010011;
ROM[39022] <= 32'b00000000000000010010010000000011;
ROM[39023] <= 32'b00000000011101000000001110110011;
ROM[39024] <= 32'b00000000011100010010000000100011;
ROM[39025] <= 32'b00000000010000010000000100010011;
ROM[39026] <= 32'b11111111110000010000000100010011;
ROM[39027] <= 32'b00000000000000010010001110000011;
ROM[39028] <= 32'b00000000000000111000001100010011;
ROM[39029] <= 32'b00000000110100110000010000110011;
ROM[39030] <= 32'b00000000000001000010001110000011;
ROM[39031] <= 32'b00000000011100010010000000100011;
ROM[39032] <= 32'b00000000010000010000000100010011;
ROM[39033] <= 32'b11111111110000010000000100010011;
ROM[39034] <= 32'b00000000000000010010001110000011;
ROM[39035] <= 32'b00000000011100011010000000100011;
ROM[39036] <= 32'b00000000110000100010001110000011;
ROM[39037] <= 32'b00000000011100010010000000100011;
ROM[39038] <= 32'b00000000010000010000000100010011;
ROM[39039] <= 32'b00000000000000011010001110000011;
ROM[39040] <= 32'b00000000011100010010000000100011;
ROM[39041] <= 32'b00000000010000010000000100010011;
ROM[39042] <= 32'b00000000100000100010001110000011;
ROM[39043] <= 32'b00000000011100010010000000100011;
ROM[39044] <= 32'b00000000010000010000000100010011;
ROM[39045] <= 32'b00000000010000000000001110010011;
ROM[39046] <= 32'b00000000011100010010000000100011;
ROM[39047] <= 32'b00000000010000010000000100010011;
ROM[39048] <= 32'b00000000000000100110001110110111;
ROM[39049] <= 32'b00100110110000111000001110010011;
ROM[39050] <= 32'b00000000111000111000001110110011;
ROM[39051] <= 32'b00000000011100010010000000100011;
ROM[39052] <= 32'b00000000010000010000000100010011;
ROM[39053] <= 32'b00000000001100010010000000100011;
ROM[39054] <= 32'b00000000010000010000000100010011;
ROM[39055] <= 32'b00000000010000010010000000100011;
ROM[39056] <= 32'b00000000010000010000000100010011;
ROM[39057] <= 32'b00000000010100010010000000100011;
ROM[39058] <= 32'b00000000010000010000000100010011;
ROM[39059] <= 32'b00000000011000010010000000100011;
ROM[39060] <= 32'b00000000010000010000000100010011;
ROM[39061] <= 32'b00000001010000000000001110010011;
ROM[39062] <= 32'b00000000100000111000001110010011;
ROM[39063] <= 32'b01000000011100010000001110110011;
ROM[39064] <= 32'b00000000011100000000001000110011;
ROM[39065] <= 32'b00000000001000000000000110110011;
ROM[39066] <= 32'b11011100010011101011000011101111;
ROM[39067] <= 32'b11111111110000010000000100010011;
ROM[39068] <= 32'b00000000000000010010001110000011;
ROM[39069] <= 32'b11111111110000010000000100010011;
ROM[39070] <= 32'b00000000000000010010010000000011;
ROM[39071] <= 32'b00000000011101000000001110110011;
ROM[39072] <= 32'b00000000011100010010000000100011;
ROM[39073] <= 32'b00000000010000010000000100010011;
ROM[39074] <= 32'b11111111110000010000000100010011;
ROM[39075] <= 32'b00000000000000010010001110000011;
ROM[39076] <= 32'b00000000000000111000001100010011;
ROM[39077] <= 32'b11111111110000010000000100010011;
ROM[39078] <= 32'b00000000000000010010001110000011;
ROM[39079] <= 32'b00000000110100110000010000110011;
ROM[39080] <= 32'b00000000011101000010000000100011;
ROM[39081] <= 32'b00000000000000000000001110010011;
ROM[39082] <= 32'b00000000011100010010000000100011;
ROM[39083] <= 32'b00000000010000010000000100010011;
ROM[39084] <= 32'b00000001010000000000001110010011;
ROM[39085] <= 32'b01000000011100011000001110110011;
ROM[39086] <= 32'b00000000000000111010000010000011;
ROM[39087] <= 32'b11111111110000010000000100010011;
ROM[39088] <= 32'b00000000000000010010001110000011;
ROM[39089] <= 32'b00000000011100100010000000100011;
ROM[39090] <= 32'b00000000010000100000000100010011;
ROM[39091] <= 32'b00000001010000000000001110010011;
ROM[39092] <= 32'b01000000011100011000001110110011;
ROM[39093] <= 32'b00000000010000111010000110000011;
ROM[39094] <= 32'b00000000100000111010001000000011;
ROM[39095] <= 32'b00000000110000111010001010000011;
ROM[39096] <= 32'b00000001000000111010001100000011;
ROM[39097] <= 32'b00000000000000001000000011100111;
ROM[39098] <= 32'b00000000000000010010000000100011;
ROM[39099] <= 32'b00000000010000010000000100010011;
ROM[39100] <= 32'b00000000000000100010001110000011;
ROM[39101] <= 32'b00000000011100010010000000100011;
ROM[39102] <= 32'b00000000010000010000000100010011;
ROM[39103] <= 32'b11111111110000010000000100010011;
ROM[39104] <= 32'b00000000000000010010001110000011;
ROM[39105] <= 32'b00000000000000111000001010010011;
ROM[39106] <= 32'b00000000110100101000010000110011;
ROM[39107] <= 32'b00000001010001000010001110000011;
ROM[39108] <= 32'b00000000011100010010000000100011;
ROM[39109] <= 32'b00000000010000010000000100010011;
ROM[39110] <= 32'b00000000010000100010001110000011;
ROM[39111] <= 32'b00000000011100010010000000100011;
ROM[39112] <= 32'b00000000010000010000000100010011;
ROM[39113] <= 32'b00000000010000000000001110010011;
ROM[39114] <= 32'b00000000011100010010000000100011;
ROM[39115] <= 32'b00000000010000010000000100010011;
ROM[39116] <= 32'b00000000000000100110001110110111;
ROM[39117] <= 32'b00110111110000111000001110010011;
ROM[39118] <= 32'b00000000111000111000001110110011;
ROM[39119] <= 32'b00000000011100010010000000100011;
ROM[39120] <= 32'b00000000010000010000000100010011;
ROM[39121] <= 32'b00000000001100010010000000100011;
ROM[39122] <= 32'b00000000010000010000000100010011;
ROM[39123] <= 32'b00000000010000010010000000100011;
ROM[39124] <= 32'b00000000010000010000000100010011;
ROM[39125] <= 32'b00000000010100010010000000100011;
ROM[39126] <= 32'b00000000010000010000000100010011;
ROM[39127] <= 32'b00000000011000010010000000100011;
ROM[39128] <= 32'b00000000010000010000000100010011;
ROM[39129] <= 32'b00000001010000000000001110010011;
ROM[39130] <= 32'b00000000100000111000001110010011;
ROM[39131] <= 32'b01000000011100010000001110110011;
ROM[39132] <= 32'b00000000011100000000001000110011;
ROM[39133] <= 32'b00000000001000000000000110110011;
ROM[39134] <= 32'b11001011010011101011000011101111;
ROM[39135] <= 32'b11111111110000010000000100010011;
ROM[39136] <= 32'b00000000000000010010001110000011;
ROM[39137] <= 32'b11111111110000010000000100010011;
ROM[39138] <= 32'b00000000000000010010010000000011;
ROM[39139] <= 32'b00000000011101000000001110110011;
ROM[39140] <= 32'b00000000011100010010000000100011;
ROM[39141] <= 32'b00000000010000010000000100010011;
ROM[39142] <= 32'b11111111110000010000000100010011;
ROM[39143] <= 32'b00000000000000010010001110000011;
ROM[39144] <= 32'b00000000000000111000001100010011;
ROM[39145] <= 32'b00000000110100110000010000110011;
ROM[39146] <= 32'b00000000000001000010001110000011;
ROM[39147] <= 32'b00000000011100010010000000100011;
ROM[39148] <= 32'b00000000010000010000000100010011;
ROM[39149] <= 32'b11111111110000010000000100010011;
ROM[39150] <= 32'b00000000000000010010001110000011;
ROM[39151] <= 32'b00000000011100011010000000100011;
ROM[39152] <= 32'b00000000000000011010001110000011;
ROM[39153] <= 32'b00000000011100010010000000100011;
ROM[39154] <= 32'b00000000010000010000000100010011;
ROM[39155] <= 32'b00000000100000100010001110000011;
ROM[39156] <= 32'b00000000011100010010000000100011;
ROM[39157] <= 32'b00000000010000010000000100010011;
ROM[39158] <= 32'b00000000010000000000001110010011;
ROM[39159] <= 32'b00000000011100010010000000100011;
ROM[39160] <= 32'b00000000010000010000000100010011;
ROM[39161] <= 32'b00000000000000100110001110110111;
ROM[39162] <= 32'b01000011000000111000001110010011;
ROM[39163] <= 32'b00000000111000111000001110110011;
ROM[39164] <= 32'b00000000011100010010000000100011;
ROM[39165] <= 32'b00000000010000010000000100010011;
ROM[39166] <= 32'b00000000001100010010000000100011;
ROM[39167] <= 32'b00000000010000010000000100010011;
ROM[39168] <= 32'b00000000010000010010000000100011;
ROM[39169] <= 32'b00000000010000010000000100010011;
ROM[39170] <= 32'b00000000010100010010000000100011;
ROM[39171] <= 32'b00000000010000010000000100010011;
ROM[39172] <= 32'b00000000011000010010000000100011;
ROM[39173] <= 32'b00000000010000010000000100010011;
ROM[39174] <= 32'b00000001010000000000001110010011;
ROM[39175] <= 32'b00000000100000111000001110010011;
ROM[39176] <= 32'b01000000011100010000001110110011;
ROM[39177] <= 32'b00000000011100000000001000110011;
ROM[39178] <= 32'b00000000001000000000000110110011;
ROM[39179] <= 32'b11000000000011101011000011101111;
ROM[39180] <= 32'b11111111110000010000000100010011;
ROM[39181] <= 32'b00000000000000010010001110000011;
ROM[39182] <= 32'b11111111110000010000000100010011;
ROM[39183] <= 32'b00000000000000010010010000000011;
ROM[39184] <= 32'b00000000011101000000001110110011;
ROM[39185] <= 32'b00000000011100010010000000100011;
ROM[39186] <= 32'b00000000010000010000000100010011;
ROM[39187] <= 32'b11111111110000010000000100010011;
ROM[39188] <= 32'b00000000000000010010001110000011;
ROM[39189] <= 32'b00000000000000111000001100010011;
ROM[39190] <= 32'b00000000110100110000010000110011;
ROM[39191] <= 32'b00000000000001000010001110000011;
ROM[39192] <= 32'b00000000011100010010000000100011;
ROM[39193] <= 32'b00000000010000010000000100010011;
ROM[39194] <= 32'b11111111110000010000000100010011;
ROM[39195] <= 32'b00000000000000010010001110000011;
ROM[39196] <= 32'b00000000000000111000101001100011;
ROM[39197] <= 32'b00000000000000100110001110110111;
ROM[39198] <= 32'b01001100110000111000001110010011;
ROM[39199] <= 32'b00000000111000111000001110110011;
ROM[39200] <= 32'b00000000000000111000000011100111;
ROM[39201] <= 32'b00000000000000000000001110010011;
ROM[39202] <= 32'b00000000011100010010000000100011;
ROM[39203] <= 32'b00000000010000010000000100010011;
ROM[39204] <= 32'b00000001010000000000001110010011;
ROM[39205] <= 32'b01000000011100011000001110110011;
ROM[39206] <= 32'b00000000000000111010000010000011;
ROM[39207] <= 32'b11111111110000010000000100010011;
ROM[39208] <= 32'b00000000000000010010001110000011;
ROM[39209] <= 32'b00000000011100100010000000100011;
ROM[39210] <= 32'b00000000010000100000000100010011;
ROM[39211] <= 32'b00000001010000000000001110010011;
ROM[39212] <= 32'b01000000011100011000001110110011;
ROM[39213] <= 32'b00000000010000111010000110000011;
ROM[39214] <= 32'b00000000100000111010001000000011;
ROM[39215] <= 32'b00000000110000111010001010000011;
ROM[39216] <= 32'b00000001000000111010001100000011;
ROM[39217] <= 32'b00000000000000001000000011100111;
ROM[39218] <= 32'b00000101110000000000000011101111;
ROM[39219] <= 32'b00000000000100000000001110010011;
ROM[39220] <= 32'b00000000011100010010000000100011;
ROM[39221] <= 32'b00000000010000010000000100010011;
ROM[39222] <= 32'b11111111110000010000000100010011;
ROM[39223] <= 32'b00000000000000010010001110000011;
ROM[39224] <= 32'b01000000011100000000001110110011;
ROM[39225] <= 32'b00000000011100010010000000100011;
ROM[39226] <= 32'b00000000010000010000000100010011;
ROM[39227] <= 32'b00000001010000000000001110010011;
ROM[39228] <= 32'b01000000011100011000001110110011;
ROM[39229] <= 32'b00000000000000111010000010000011;
ROM[39230] <= 32'b11111111110000010000000100010011;
ROM[39231] <= 32'b00000000000000010010001110000011;
ROM[39232] <= 32'b00000000011100100010000000100011;
ROM[39233] <= 32'b00000000010000100000000100010011;
ROM[39234] <= 32'b00000001010000000000001110010011;
ROM[39235] <= 32'b01000000011100011000001110110011;
ROM[39236] <= 32'b00000000010000111010000110000011;
ROM[39237] <= 32'b00000000100000111010001000000011;
ROM[39238] <= 32'b00000000110000111010001010000011;
ROM[39239] <= 32'b00000001000000111010001100000011;
ROM[39240] <= 32'b00000000000000001000000011100111;
ROM[39241] <= 32'b00000000000000100010001110000011;
ROM[39242] <= 32'b00000000011100010010000000100011;
ROM[39243] <= 32'b00000000010000010000000100010011;
ROM[39244] <= 32'b11111111110000010000000100010011;
ROM[39245] <= 32'b00000000000000010010001110000011;
ROM[39246] <= 32'b00000000000000111000001010010011;
ROM[39247] <= 32'b00000000010000100010001110000011;
ROM[39248] <= 32'b00000000011100010010000000100011;
ROM[39249] <= 32'b00000000010000010000000100010011;
ROM[39250] <= 32'b00000000110100101000010000110011;
ROM[39251] <= 32'b00000000110001000010001110000011;
ROM[39252] <= 32'b00000000011100010010000000100011;
ROM[39253] <= 32'b00000000010000010000000100010011;
ROM[39254] <= 32'b11111111110000010000000100010011;
ROM[39255] <= 32'b00000000000000010010001110000011;
ROM[39256] <= 32'b11111111110000010000000100010011;
ROM[39257] <= 32'b00000000000000010010010000000011;
ROM[39258] <= 32'b00000000011101000010010010110011;
ROM[39259] <= 32'b00000000100000111010010100110011;
ROM[39260] <= 32'b00000000101001001000001110110011;
ROM[39261] <= 32'b00000000000100111000001110010011;
ROM[39262] <= 32'b00000000000100111111001110010011;
ROM[39263] <= 32'b00000000011100010010000000100011;
ROM[39264] <= 32'b00000000010000010000000100010011;
ROM[39265] <= 32'b11111111110000010000000100010011;
ROM[39266] <= 32'b00000000000000010010001110000011;
ROM[39267] <= 32'b00000000000000111000101001100011;
ROM[39268] <= 32'b00000000000000100110001110110111;
ROM[39269] <= 32'b01011010010000111000001110010011;
ROM[39270] <= 32'b00000000111000111000001110110011;
ROM[39271] <= 32'b00000000000000111000000011100111;
ROM[39272] <= 32'b00001100010000000000000011101111;
ROM[39273] <= 32'b00000000100000100010001110000011;
ROM[39274] <= 32'b00000000011100010010000000100011;
ROM[39275] <= 32'b00000000010000010000000100010011;
ROM[39276] <= 32'b00000000110100101000010000110011;
ROM[39277] <= 32'b00000001000001000010001110000011;
ROM[39278] <= 32'b00000000011100010010000000100011;
ROM[39279] <= 32'b00000000010000010000000100010011;
ROM[39280] <= 32'b11111111110000010000000100010011;
ROM[39281] <= 32'b00000000000000010010001110000011;
ROM[39282] <= 32'b11111111110000010000000100010011;
ROM[39283] <= 32'b00000000000000010010010000000011;
ROM[39284] <= 32'b00000000011101000010010010110011;
ROM[39285] <= 32'b00000000100000111010010100110011;
ROM[39286] <= 32'b00000000101001001000001110110011;
ROM[39287] <= 32'b00000000000100111000001110010011;
ROM[39288] <= 32'b00000000000100111111001110010011;
ROM[39289] <= 32'b00000000011100010010000000100011;
ROM[39290] <= 32'b00000000010000010000000100010011;
ROM[39291] <= 32'b11111111110000010000000100010011;
ROM[39292] <= 32'b00000000000000010010001110000011;
ROM[39293] <= 32'b00000000000000111000101001100011;
ROM[39294] <= 32'b00000000000000100110001110110111;
ROM[39295] <= 32'b01100000110000111000001110010011;
ROM[39296] <= 32'b00000000111000111000001110110011;
ROM[39297] <= 32'b00000000000000111000000011100111;
ROM[39298] <= 32'b00000101110000000000000011101111;
ROM[39299] <= 32'b00000000000100000000001110010011;
ROM[39300] <= 32'b00000000011100010010000000100011;
ROM[39301] <= 32'b00000000010000010000000100010011;
ROM[39302] <= 32'b11111111110000010000000100010011;
ROM[39303] <= 32'b00000000000000010010001110000011;
ROM[39304] <= 32'b01000000011100000000001110110011;
ROM[39305] <= 32'b00000000011100010010000000100011;
ROM[39306] <= 32'b00000000010000010000000100010011;
ROM[39307] <= 32'b00000001010000000000001110010011;
ROM[39308] <= 32'b01000000011100011000001110110011;
ROM[39309] <= 32'b00000000000000111010000010000011;
ROM[39310] <= 32'b11111111110000010000000100010011;
ROM[39311] <= 32'b00000000000000010010001110000011;
ROM[39312] <= 32'b00000000011100100010000000100011;
ROM[39313] <= 32'b00000000010000100000000100010011;
ROM[39314] <= 32'b00000001010000000000001110010011;
ROM[39315] <= 32'b01000000011100011000001110110011;
ROM[39316] <= 32'b00000000010000111010000110000011;
ROM[39317] <= 32'b00000000100000111010001000000011;
ROM[39318] <= 32'b00000000110000111010001010000011;
ROM[39319] <= 32'b00000001000000111010001100000011;
ROM[39320] <= 32'b00000000000000001000000011100111;
ROM[39321] <= 32'b00000000000000000000001110010011;
ROM[39322] <= 32'b00000000011100010010000000100011;
ROM[39323] <= 32'b00000000010000010000000100010011;
ROM[39324] <= 32'b00000001010000000000001110010011;
ROM[39325] <= 32'b01000000011100011000001110110011;
ROM[39326] <= 32'b00000000000000111010000010000011;
ROM[39327] <= 32'b11111111110000010000000100010011;
ROM[39328] <= 32'b00000000000000010010001110000011;
ROM[39329] <= 32'b00000000011100100010000000100011;
ROM[39330] <= 32'b00000000010000100000000100010011;
ROM[39331] <= 32'b00000001010000000000001110010011;
ROM[39332] <= 32'b01000000011100011000001110110011;
ROM[39333] <= 32'b00000000010000111010000110000011;
ROM[39334] <= 32'b00000000100000111010001000000011;
ROM[39335] <= 32'b00000000110000111010001010000011;
ROM[39336] <= 32'b00000001000000111010001100000011;
ROM[39337] <= 32'b00000000000000001000000011100111;
ROM[39338] <= 32'b00000000000000100010001110000011;
ROM[39339] <= 32'b00000000011100010010000000100011;
ROM[39340] <= 32'b00000000010000010000000100010011;
ROM[39341] <= 32'b11111111110000010000000100010011;
ROM[39342] <= 32'b00000000000000010010001110000011;
ROM[39343] <= 32'b00000000000000111000001010010011;
ROM[39344] <= 32'b00000001011000000000001110010011;
ROM[39345] <= 32'b00000000011100010010000000100011;
ROM[39346] <= 32'b00000000010000010000000100010011;
ROM[39347] <= 32'b00000001010100000000001110010011;
ROM[39348] <= 32'b00000000011100010010000000100011;
ROM[39349] <= 32'b00000000010000010000000100010011;
ROM[39350] <= 32'b00000000000000100110001110110111;
ROM[39351] <= 32'b01110010010000111000001110010011;
ROM[39352] <= 32'b00000000111000111000001110110011;
ROM[39353] <= 32'b00000000011100010010000000100011;
ROM[39354] <= 32'b00000000010000010000000100010011;
ROM[39355] <= 32'b00000000001100010010000000100011;
ROM[39356] <= 32'b00000000010000010000000100010011;
ROM[39357] <= 32'b00000000010000010010000000100011;
ROM[39358] <= 32'b00000000010000010000000100010011;
ROM[39359] <= 32'b00000000010100010010000000100011;
ROM[39360] <= 32'b00000000010000010000000100010011;
ROM[39361] <= 32'b00000000011000010010000000100011;
ROM[39362] <= 32'b00000000010000010000000100010011;
ROM[39363] <= 32'b00000001010000000000001110010011;
ROM[39364] <= 32'b00000000100000111000001110010011;
ROM[39365] <= 32'b01000000011100010000001110110011;
ROM[39366] <= 32'b00000000011100000000001000110011;
ROM[39367] <= 32'b00000000001000000000000110110011;
ROM[39368] <= 32'b11001110000011101111000011101111;
ROM[39369] <= 32'b11111111110000010000000100010011;
ROM[39370] <= 32'b00000000000000010010001110000011;
ROM[39371] <= 32'b00000000011101100010000000100011;
ROM[39372] <= 32'b00000000110100101000010000110011;
ROM[39373] <= 32'b00000000000001000010001110000011;
ROM[39374] <= 32'b00000000011100010010000000100011;
ROM[39375] <= 32'b00000000010000010000000100010011;
ROM[39376] <= 32'b00000000000000100110001110110111;
ROM[39377] <= 32'b01111000110000111000001110010011;
ROM[39378] <= 32'b00000000111000111000001110110011;
ROM[39379] <= 32'b00000000011100010010000000100011;
ROM[39380] <= 32'b00000000010000010000000100010011;
ROM[39381] <= 32'b00000000001100010010000000100011;
ROM[39382] <= 32'b00000000010000010000000100010011;
ROM[39383] <= 32'b00000000010000010010000000100011;
ROM[39384] <= 32'b00000000010000010000000100010011;
ROM[39385] <= 32'b00000000010100010010000000100011;
ROM[39386] <= 32'b00000000010000010000000100010011;
ROM[39387] <= 32'b00000000011000010010000000100011;
ROM[39388] <= 32'b00000000010000010000000100010011;
ROM[39389] <= 32'b00000001010000000000001110010011;
ROM[39390] <= 32'b00000000010000111000001110010011;
ROM[39391] <= 32'b01000000011100010000001110110011;
ROM[39392] <= 32'b00000000011100000000001000110011;
ROM[39393] <= 32'b00000000001000000000000110110011;
ROM[39394] <= 32'b10111001110011111101000011101111;
ROM[39395] <= 32'b00000000000000100110001110110111;
ROM[39396] <= 32'b01111101100000111000001110010011;
ROM[39397] <= 32'b00000000111000111000001110110011;
ROM[39398] <= 32'b00000000011100010010000000100011;
ROM[39399] <= 32'b00000000010000010000000100010011;
ROM[39400] <= 32'b00000000001100010010000000100011;
ROM[39401] <= 32'b00000000010000010000000100010011;
ROM[39402] <= 32'b00000000010000010010000000100011;
ROM[39403] <= 32'b00000000010000010000000100010011;
ROM[39404] <= 32'b00000000010100010010000000100011;
ROM[39405] <= 32'b00000000010000010000000100010011;
ROM[39406] <= 32'b00000000011000010010000000100011;
ROM[39407] <= 32'b00000000010000010000000100010011;
ROM[39408] <= 32'b00000001010000000000001110010011;
ROM[39409] <= 32'b00000000010000111000001110010011;
ROM[39410] <= 32'b01000000011100010000001110110011;
ROM[39411] <= 32'b00000000011100000000001000110011;
ROM[39412] <= 32'b00000000001000000000000110110011;
ROM[39413] <= 32'b10011010110111110000000011101111;
ROM[39414] <= 32'b11111111110000010000000100010011;
ROM[39415] <= 32'b00000000000000010010001110000011;
ROM[39416] <= 32'b00000000011101100010000000100011;
ROM[39417] <= 32'b00000001011000000000001110010011;
ROM[39418] <= 32'b00000000011100010010000000100011;
ROM[39419] <= 32'b00000000010000010000000100010011;
ROM[39420] <= 32'b00000010101000000000001110010011;
ROM[39421] <= 32'b00000000011100010010000000100011;
ROM[39422] <= 32'b00000000010000010000000100010011;
ROM[39423] <= 32'b00000000000000100111001110110111;
ROM[39424] <= 32'b10000100100000111000001110010011;
ROM[39425] <= 32'b00000000111000111000001110110011;
ROM[39426] <= 32'b00000000011100010010000000100011;
ROM[39427] <= 32'b00000000010000010000000100010011;
ROM[39428] <= 32'b00000000001100010010000000100011;
ROM[39429] <= 32'b00000000010000010000000100010011;
ROM[39430] <= 32'b00000000010000010010000000100011;
ROM[39431] <= 32'b00000000010000010000000100010011;
ROM[39432] <= 32'b00000000010100010010000000100011;
ROM[39433] <= 32'b00000000010000010000000100010011;
ROM[39434] <= 32'b00000000011000010010000000100011;
ROM[39435] <= 32'b00000000010000010000000100010011;
ROM[39436] <= 32'b00000001010000000000001110010011;
ROM[39437] <= 32'b00000000100000111000001110010011;
ROM[39438] <= 32'b01000000011100010000001110110011;
ROM[39439] <= 32'b00000000011100000000001000110011;
ROM[39440] <= 32'b00000000001000000000000110110011;
ROM[39441] <= 32'b10111011110011101111000011101111;
ROM[39442] <= 32'b11111111110000010000000100010011;
ROM[39443] <= 32'b00000000000000010010001110000011;
ROM[39444] <= 32'b00000000011101100010000000100011;
ROM[39445] <= 32'b00000000010000100010001110000011;
ROM[39446] <= 32'b00000000011100010010000000100011;
ROM[39447] <= 32'b00000000010000010000000100010011;
ROM[39448] <= 32'b00000000000000100111001110110111;
ROM[39449] <= 32'b10001010110000111000001110010011;
ROM[39450] <= 32'b00000000111000111000001110110011;
ROM[39451] <= 32'b00000000011100010010000000100011;
ROM[39452] <= 32'b00000000010000010000000100010011;
ROM[39453] <= 32'b00000000001100010010000000100011;
ROM[39454] <= 32'b00000000010000010000000100010011;
ROM[39455] <= 32'b00000000010000010010000000100011;
ROM[39456] <= 32'b00000000010000010000000100010011;
ROM[39457] <= 32'b00000000010100010010000000100011;
ROM[39458] <= 32'b00000000010000010000000100010011;
ROM[39459] <= 32'b00000000011000010010000000100011;
ROM[39460] <= 32'b00000000010000010000000100010011;
ROM[39461] <= 32'b00000001010000000000001110010011;
ROM[39462] <= 32'b00000000010000111000001110010011;
ROM[39463] <= 32'b01000000011100010000001110110011;
ROM[39464] <= 32'b00000000011100000000001000110011;
ROM[39465] <= 32'b00000000001000000000000110110011;
ROM[39466] <= 32'b10001101100111110000000011101111;
ROM[39467] <= 32'b11111111110000010000000100010011;
ROM[39468] <= 32'b00000000000000010010001110000011;
ROM[39469] <= 32'b00000000011101100010000000100011;
ROM[39470] <= 32'b00000001011000000000001110010011;
ROM[39471] <= 32'b00000000011100010010000000100011;
ROM[39472] <= 32'b00000000010000010000000100010011;
ROM[39473] <= 32'b00000010111000000000001110010011;
ROM[39474] <= 32'b00000000011100010010000000100011;
ROM[39475] <= 32'b00000000010000010000000100010011;
ROM[39476] <= 32'b00000000000000100111001110110111;
ROM[39477] <= 32'b10010001110000111000001110010011;
ROM[39478] <= 32'b00000000111000111000001110110011;
ROM[39479] <= 32'b00000000011100010010000000100011;
ROM[39480] <= 32'b00000000010000010000000100010011;
ROM[39481] <= 32'b00000000001100010010000000100011;
ROM[39482] <= 32'b00000000010000010000000100010011;
ROM[39483] <= 32'b00000000010000010010000000100011;
ROM[39484] <= 32'b00000000010000010000000100010011;
ROM[39485] <= 32'b00000000010100010010000000100011;
ROM[39486] <= 32'b00000000010000010000000100010011;
ROM[39487] <= 32'b00000000011000010010000000100011;
ROM[39488] <= 32'b00000000010000010000000100010011;
ROM[39489] <= 32'b00000001010000000000001110010011;
ROM[39490] <= 32'b00000000100000111000001110010011;
ROM[39491] <= 32'b01000000011100010000001110110011;
ROM[39492] <= 32'b00000000011100000000001000110011;
ROM[39493] <= 32'b00000000001000000000000110110011;
ROM[39494] <= 32'b10101110100011101111000011101111;
ROM[39495] <= 32'b11111111110000010000000100010011;
ROM[39496] <= 32'b00000000000000010010001110000011;
ROM[39497] <= 32'b00000000011101100010000000100011;
ROM[39498] <= 32'b00000000100000100010001110000011;
ROM[39499] <= 32'b00000000011100010010000000100011;
ROM[39500] <= 32'b00000000010000010000000100010011;
ROM[39501] <= 32'b00000000000000100111001110110111;
ROM[39502] <= 32'b10011000000000111000001110010011;
ROM[39503] <= 32'b00000000111000111000001110110011;
ROM[39504] <= 32'b00000000011100010010000000100011;
ROM[39505] <= 32'b00000000010000010000000100010011;
ROM[39506] <= 32'b00000000001100010010000000100011;
ROM[39507] <= 32'b00000000010000010000000100010011;
ROM[39508] <= 32'b00000000010000010010000000100011;
ROM[39509] <= 32'b00000000010000010000000100010011;
ROM[39510] <= 32'b00000000010100010010000000100011;
ROM[39511] <= 32'b00000000010000010000000100010011;
ROM[39512] <= 32'b00000000011000010010000000100011;
ROM[39513] <= 32'b00000000010000010000000100010011;
ROM[39514] <= 32'b00000001010000000000001110010011;
ROM[39515] <= 32'b00000000010000111000001110010011;
ROM[39516] <= 32'b01000000011100010000001110110011;
ROM[39517] <= 32'b00000000011100000000001000110011;
ROM[39518] <= 32'b00000000001000000000000110110011;
ROM[39519] <= 32'b10000000010111110000000011101111;
ROM[39520] <= 32'b11111111110000010000000100010011;
ROM[39521] <= 32'b00000000000000010010001110000011;
ROM[39522] <= 32'b00000000011101100010000000100011;
ROM[39523] <= 32'b00000000000000000000001110010011;
ROM[39524] <= 32'b00000000011100010010000000100011;
ROM[39525] <= 32'b00000000010000010000000100010011;
ROM[39526] <= 32'b00000001010000000000001110010011;
ROM[39527] <= 32'b01000000011100011000001110110011;
ROM[39528] <= 32'b00000000000000111010000010000011;
ROM[39529] <= 32'b11111111110000010000000100010011;
ROM[39530] <= 32'b00000000000000010010001110000011;
ROM[39531] <= 32'b00000000011100100010000000100011;
ROM[39532] <= 32'b00000000010000100000000100010011;
ROM[39533] <= 32'b00000001010000000000001110010011;
ROM[39534] <= 32'b01000000011100011000001110110011;
ROM[39535] <= 32'b00000000010000111010000110000011;
ROM[39536] <= 32'b00000000100000111010001000000011;
ROM[39537] <= 32'b00000000110000111010001010000011;
ROM[39538] <= 32'b00000001000000111010001100000011;
ROM[39539] <= 32'b00000000000000001000000011100111;
ROM[39540] <= 32'b00000000000000100010001110000011;
ROM[39541] <= 32'b00000000011100010010000000100011;
ROM[39542] <= 32'b00000000010000010000000100010011;
ROM[39543] <= 32'b11111111110000010000000100010011;
ROM[39544] <= 32'b00000000000000010010001110000011;
ROM[39545] <= 32'b00000000000000111000001010010011;
ROM[39546] <= 32'b00000000000100000000001110010011;
ROM[39547] <= 32'b00000000011100010010000000100011;
ROM[39548] <= 32'b00000000010000010000000100010011;
ROM[39549] <= 32'b11111111110000010000000100010011;
ROM[39550] <= 32'b00000000000000010010001110000011;
ROM[39551] <= 32'b01000000011100000000001110110011;
ROM[39552] <= 32'b00000000011100010010000000100011;
ROM[39553] <= 32'b00000000010000010000000100010011;
ROM[39554] <= 32'b00000000000000100111001110110111;
ROM[39555] <= 32'b10100101010000111000001110010011;
ROM[39556] <= 32'b00000000111000111000001110110011;
ROM[39557] <= 32'b00000000011100010010000000100011;
ROM[39558] <= 32'b00000000010000010000000100010011;
ROM[39559] <= 32'b00000000001100010010000000100011;
ROM[39560] <= 32'b00000000010000010000000100010011;
ROM[39561] <= 32'b00000000010000010010000000100011;
ROM[39562] <= 32'b00000000010000010000000100010011;
ROM[39563] <= 32'b00000000010100010010000000100011;
ROM[39564] <= 32'b00000000010000010000000100010011;
ROM[39565] <= 32'b00000000011000010010000000100011;
ROM[39566] <= 32'b00000000010000010000000100010011;
ROM[39567] <= 32'b00000001010000000000001110010011;
ROM[39568] <= 32'b00000000010000111000001110010011;
ROM[39569] <= 32'b01000000011100010000001110110011;
ROM[39570] <= 32'b00000000011100000000001000110011;
ROM[39571] <= 32'b00000000001000000000000110110011;
ROM[39572] <= 32'b11100000000011110111000011101111;
ROM[39573] <= 32'b11111111110000010000000100010011;
ROM[39574] <= 32'b00000000000000010010001110000011;
ROM[39575] <= 32'b00000000011101100010000000100011;
ROM[39576] <= 32'b00000000010000100010001110000011;
ROM[39577] <= 32'b00000000011100010010000000100011;
ROM[39578] <= 32'b00000000010000010000000100010011;
ROM[39579] <= 32'b00000000010000000000001110010011;
ROM[39580] <= 32'b00000000011100010010000000100011;
ROM[39581] <= 32'b00000000010000010000000100010011;
ROM[39582] <= 32'b00000000000000100111001110110111;
ROM[39583] <= 32'b10101100010000111000001110010011;
ROM[39584] <= 32'b00000000111000111000001110110011;
ROM[39585] <= 32'b00000000011100010010000000100011;
ROM[39586] <= 32'b00000000010000010000000100010011;
ROM[39587] <= 32'b00000000001100010010000000100011;
ROM[39588] <= 32'b00000000010000010000000100010011;
ROM[39589] <= 32'b00000000010000010010000000100011;
ROM[39590] <= 32'b00000000010000010000000100010011;
ROM[39591] <= 32'b00000000010100010010000000100011;
ROM[39592] <= 32'b00000000010000010000000100010011;
ROM[39593] <= 32'b00000000011000010010000000100011;
ROM[39594] <= 32'b00000000010000010000000100010011;
ROM[39595] <= 32'b00000001010000000000001110010011;
ROM[39596] <= 32'b00000000100000111000001110010011;
ROM[39597] <= 32'b01000000011100010000001110110011;
ROM[39598] <= 32'b00000000011100000000001000110011;
ROM[39599] <= 32'b00000000001000000000000110110011;
ROM[39600] <= 32'b11010110110111101010000011101111;
ROM[39601] <= 32'b00000000100000100010001110000011;
ROM[39602] <= 32'b00000000011100010010000000100011;
ROM[39603] <= 32'b00000000010000010000000100010011;
ROM[39604] <= 32'b00000000010000000000001110010011;
ROM[39605] <= 32'b00000000011100010010000000100011;
ROM[39606] <= 32'b00000000010000010000000100010011;
ROM[39607] <= 32'b00000000000000100111001110110111;
ROM[39608] <= 32'b10110010100000111000001110010011;
ROM[39609] <= 32'b00000000111000111000001110110011;
ROM[39610] <= 32'b00000000011100010010000000100011;
ROM[39611] <= 32'b00000000010000010000000100010011;
ROM[39612] <= 32'b00000000001100010010000000100011;
ROM[39613] <= 32'b00000000010000010000000100010011;
ROM[39614] <= 32'b00000000010000010010000000100011;
ROM[39615] <= 32'b00000000010000010000000100010011;
ROM[39616] <= 32'b00000000010100010010000000100011;
ROM[39617] <= 32'b00000000010000010000000100010011;
ROM[39618] <= 32'b00000000011000010010000000100011;
ROM[39619] <= 32'b00000000010000010000000100010011;
ROM[39620] <= 32'b00000001010000000000001110010011;
ROM[39621] <= 32'b00000000100000111000001110010011;
ROM[39622] <= 32'b01000000011100010000001110110011;
ROM[39623] <= 32'b00000000011100000000001000110011;
ROM[39624] <= 32'b00000000001000000000000110110011;
ROM[39625] <= 32'b11010000100111101010000011101111;
ROM[39626] <= 32'b00000000010000100010001110000011;
ROM[39627] <= 32'b00000000011100010010000000100011;
ROM[39628] <= 32'b00000000010000010000000100010011;
ROM[39629] <= 32'b00000000010000000000001110010011;
ROM[39630] <= 32'b00000000011100010010000000100011;
ROM[39631] <= 32'b00000000010000010000000100010011;
ROM[39632] <= 32'b00000000000000100111001110110111;
ROM[39633] <= 32'b10111000110000111000001110010011;
ROM[39634] <= 32'b00000000111000111000001110110011;
ROM[39635] <= 32'b00000000011100010010000000100011;
ROM[39636] <= 32'b00000000010000010000000100010011;
ROM[39637] <= 32'b00000000001100010010000000100011;
ROM[39638] <= 32'b00000000010000010000000100010011;
ROM[39639] <= 32'b00000000010000010010000000100011;
ROM[39640] <= 32'b00000000010000010000000100010011;
ROM[39641] <= 32'b00000000010100010010000000100011;
ROM[39642] <= 32'b00000000010000010000000100010011;
ROM[39643] <= 32'b00000000011000010010000000100011;
ROM[39644] <= 32'b00000000010000010000000100010011;
ROM[39645] <= 32'b00000001010000000000001110010011;
ROM[39646] <= 32'b00000000100000111000001110010011;
ROM[39647] <= 32'b01000000011100010000001110110011;
ROM[39648] <= 32'b00000000011100000000001000110011;
ROM[39649] <= 32'b00000000001000000000000110110011;
ROM[39650] <= 32'b11001010010111101010000011101111;
ROM[39651] <= 32'b00000000010000000000001110010011;
ROM[39652] <= 32'b00000000011100010010000000100011;
ROM[39653] <= 32'b00000000010000010000000100010011;
ROM[39654] <= 32'b11111111110000010000000100010011;
ROM[39655] <= 32'b00000000000000010010001110000011;
ROM[39656] <= 32'b11111111110000010000000100010011;
ROM[39657] <= 32'b00000000000000010010010000000011;
ROM[39658] <= 32'b00000000011101000000001110110011;
ROM[39659] <= 32'b00000000011100010010000000100011;
ROM[39660] <= 32'b00000000010000010000000100010011;
ROM[39661] <= 32'b00000000100000100010001110000011;
ROM[39662] <= 32'b00000000011100010010000000100011;
ROM[39663] <= 32'b00000000010000010000000100010011;
ROM[39664] <= 32'b00000000010000000000001110010011;
ROM[39665] <= 32'b00000000011100010010000000100011;
ROM[39666] <= 32'b00000000010000010000000100010011;
ROM[39667] <= 32'b00000000000000100111001110110111;
ROM[39668] <= 32'b11000001100000111000001110010011;
ROM[39669] <= 32'b00000000111000111000001110110011;
ROM[39670] <= 32'b00000000011100010010000000100011;
ROM[39671] <= 32'b00000000010000010000000100010011;
ROM[39672] <= 32'b00000000001100010010000000100011;
ROM[39673] <= 32'b00000000010000010000000100010011;
ROM[39674] <= 32'b00000000010000010010000000100011;
ROM[39675] <= 32'b00000000010000010000000100010011;
ROM[39676] <= 32'b00000000010100010010000000100011;
ROM[39677] <= 32'b00000000010000010000000100010011;
ROM[39678] <= 32'b00000000011000010010000000100011;
ROM[39679] <= 32'b00000000010000010000000100010011;
ROM[39680] <= 32'b00000001010000000000001110010011;
ROM[39681] <= 32'b00000000100000111000001110010011;
ROM[39682] <= 32'b01000000011100010000001110110011;
ROM[39683] <= 32'b00000000011100000000001000110011;
ROM[39684] <= 32'b00000000001000000000000110110011;
ROM[39685] <= 32'b11000001100111101010000011101111;
ROM[39686] <= 32'b00000000010000000000001110010011;
ROM[39687] <= 32'b00000000011100010010000000100011;
ROM[39688] <= 32'b00000000010000010000000100010011;
ROM[39689] <= 32'b11111111110000010000000100010011;
ROM[39690] <= 32'b00000000000000010010001110000011;
ROM[39691] <= 32'b11111111110000010000000100010011;
ROM[39692] <= 32'b00000000000000010010010000000011;
ROM[39693] <= 32'b00000000011101000000001110110011;
ROM[39694] <= 32'b00000000011100010010000000100011;
ROM[39695] <= 32'b00000000010000010000000100010011;
ROM[39696] <= 32'b00000000000000100111001110110111;
ROM[39697] <= 32'b11001000110000111000001110010011;
ROM[39698] <= 32'b00000000111000111000001110110011;
ROM[39699] <= 32'b00000000011100010010000000100011;
ROM[39700] <= 32'b00000000010000010000000100010011;
ROM[39701] <= 32'b00000000001100010010000000100011;
ROM[39702] <= 32'b00000000010000010000000100010011;
ROM[39703] <= 32'b00000000010000010010000000100011;
ROM[39704] <= 32'b00000000010000010000000100010011;
ROM[39705] <= 32'b00000000010100010010000000100011;
ROM[39706] <= 32'b00000000010000010000000100010011;
ROM[39707] <= 32'b00000000011000010010000000100011;
ROM[39708] <= 32'b00000000010000010000000100010011;
ROM[39709] <= 32'b00000001010000000000001110010011;
ROM[39710] <= 32'b00000001000000111000001110010011;
ROM[39711] <= 32'b01000000011100010000001110110011;
ROM[39712] <= 32'b00000000011100000000001000110011;
ROM[39713] <= 32'b00000000001000000000000110110011;
ROM[39714] <= 32'b11110101110011111000000011101111;
ROM[39715] <= 32'b11111111110000010000000100010011;
ROM[39716] <= 32'b00000000000000010010001110000011;
ROM[39717] <= 32'b00000000011101100010000000100011;
ROM[39718] <= 32'b00000000010100010010000000100011;
ROM[39719] <= 32'b00000000010000010000000100010011;
ROM[39720] <= 32'b00000000010000100010001110000011;
ROM[39721] <= 32'b00000000011100010010000000100011;
ROM[39722] <= 32'b00000000010000010000000100010011;
ROM[39723] <= 32'b00000000100000100010001110000011;
ROM[39724] <= 32'b00000000011100010010000000100011;
ROM[39725] <= 32'b00000000010000010000000100010011;
ROM[39726] <= 32'b00000000000100000000001110010011;
ROM[39727] <= 32'b00000000011100010010000000100011;
ROM[39728] <= 32'b00000000010000010000000100010011;
ROM[39729] <= 32'b11111111110000010000000100010011;
ROM[39730] <= 32'b00000000000000010010001110000011;
ROM[39731] <= 32'b01000000011100000000001110110011;
ROM[39732] <= 32'b00000000011100010010000000100011;
ROM[39733] <= 32'b00000000010000010000000100010011;
ROM[39734] <= 32'b00000000000000100111001110110111;
ROM[39735] <= 32'b11010010010000111000001110010011;
ROM[39736] <= 32'b00000000111000111000001110110011;
ROM[39737] <= 32'b00000000011100010010000000100011;
ROM[39738] <= 32'b00000000010000010000000100010011;
ROM[39739] <= 32'b00000000001100010010000000100011;
ROM[39740] <= 32'b00000000010000010000000100010011;
ROM[39741] <= 32'b00000000010000010010000000100011;
ROM[39742] <= 32'b00000000010000010000000100010011;
ROM[39743] <= 32'b00000000010100010010000000100011;
ROM[39744] <= 32'b00000000010000010000000100010011;
ROM[39745] <= 32'b00000000011000010010000000100011;
ROM[39746] <= 32'b00000000010000010000000100010011;
ROM[39747] <= 32'b00000001010000000000001110010011;
ROM[39748] <= 32'b00000001000000111000001110010011;
ROM[39749] <= 32'b01000000011100010000001110110011;
ROM[39750] <= 32'b00000000011100000000001000110011;
ROM[39751] <= 32'b00000000001000000000000110110011;
ROM[39752] <= 32'b10111111100011111111000011101111;
ROM[39753] <= 32'b11111111110000010000000100010011;
ROM[39754] <= 32'b00000000000000010010001110000011;
ROM[39755] <= 32'b00000000011101100010000000100011;
ROM[39756] <= 32'b00000000000000000000001110010011;
ROM[39757] <= 32'b00000000011100010010000000100011;
ROM[39758] <= 32'b00000000010000010000000100010011;
ROM[39759] <= 32'b00000001010000000000001110010011;
ROM[39760] <= 32'b01000000011100011000001110110011;
ROM[39761] <= 32'b00000000000000111010000010000011;
ROM[39762] <= 32'b11111111110000010000000100010011;
ROM[39763] <= 32'b00000000000000010010001110000011;
ROM[39764] <= 32'b00000000011100100010000000100011;
ROM[39765] <= 32'b00000000010000100000000100010011;
ROM[39766] <= 32'b00000001010000000000001110010011;
ROM[39767] <= 32'b01000000011100011000001110110011;
ROM[39768] <= 32'b00000000010000111010000110000011;
ROM[39769] <= 32'b00000000100000111010001000000011;
ROM[39770] <= 32'b00000000110000111010001010000011;
ROM[39771] <= 32'b00000001000000111010001100000011;
ROM[39772] <= 32'b00000000000000001000000011100111;
ROM[39773] <= 32'b00000000000000100010001110000011;
ROM[39774] <= 32'b00000000011100010010000000100011;
ROM[39775] <= 32'b00000000010000010000000100010011;
ROM[39776] <= 32'b11111111110000010000000100010011;
ROM[39777] <= 32'b00000000000000010010001110000011;
ROM[39778] <= 32'b00000000000000111000001010010011;
ROM[39779] <= 32'b00000000000000000000001110010011;
ROM[39780] <= 32'b00000000011100010010000000100011;
ROM[39781] <= 32'b00000000010000010000000100010011;
ROM[39782] <= 32'b00000000000000100111001110110111;
ROM[39783] <= 32'b11011110010000111000001110010011;
ROM[39784] <= 32'b00000000111000111000001110110011;
ROM[39785] <= 32'b00000000011100010010000000100011;
ROM[39786] <= 32'b00000000010000010000000100010011;
ROM[39787] <= 32'b00000000001100010010000000100011;
ROM[39788] <= 32'b00000000010000010000000100010011;
ROM[39789] <= 32'b00000000010000010010000000100011;
ROM[39790] <= 32'b00000000010000010000000100010011;
ROM[39791] <= 32'b00000000010100010010000000100011;
ROM[39792] <= 32'b00000000010000010000000100010011;
ROM[39793] <= 32'b00000000011000010010000000100011;
ROM[39794] <= 32'b00000000010000010000000100010011;
ROM[39795] <= 32'b00000001010000000000001110010011;
ROM[39796] <= 32'b00000000010000111000001110010011;
ROM[39797] <= 32'b01000000011100010000001110110011;
ROM[39798] <= 32'b00000000011100000000001000110011;
ROM[39799] <= 32'b00000000001000000000000110110011;
ROM[39800] <= 32'b10100111000011110111000011101111;
ROM[39801] <= 32'b11111111110000010000000100010011;
ROM[39802] <= 32'b00000000000000010010001110000011;
ROM[39803] <= 32'b00000000011101100010000000100011;
ROM[39804] <= 32'b00000000010000100010001110000011;
ROM[39805] <= 32'b00000000011100010010000000100011;
ROM[39806] <= 32'b00000000010000010000000100010011;
ROM[39807] <= 32'b00000000010000000000001110010011;
ROM[39808] <= 32'b00000000011100010010000000100011;
ROM[39809] <= 32'b00000000010000010000000100010011;
ROM[39810] <= 32'b00000000000000100111001110110111;
ROM[39811] <= 32'b11100101010000111000001110010011;
ROM[39812] <= 32'b00000000111000111000001110110011;
ROM[39813] <= 32'b00000000011100010010000000100011;
ROM[39814] <= 32'b00000000010000010000000100010011;
ROM[39815] <= 32'b00000000001100010010000000100011;
ROM[39816] <= 32'b00000000010000010000000100010011;
ROM[39817] <= 32'b00000000010000010010000000100011;
ROM[39818] <= 32'b00000000010000010000000100010011;
ROM[39819] <= 32'b00000000010100010010000000100011;
ROM[39820] <= 32'b00000000010000010000000100010011;
ROM[39821] <= 32'b00000000011000010010000000100011;
ROM[39822] <= 32'b00000000010000010000000100010011;
ROM[39823] <= 32'b00000001010000000000001110010011;
ROM[39824] <= 32'b00000000100000111000001110010011;
ROM[39825] <= 32'b01000000011100010000001110110011;
ROM[39826] <= 32'b00000000011100000000001000110011;
ROM[39827] <= 32'b00000000001000000000000110110011;
ROM[39828] <= 32'b10011101110111101010000011101111;
ROM[39829] <= 32'b00000000100000100010001110000011;
ROM[39830] <= 32'b00000000011100010010000000100011;
ROM[39831] <= 32'b00000000010000010000000100010011;
ROM[39832] <= 32'b00000000010000000000001110010011;
ROM[39833] <= 32'b00000000011100010010000000100011;
ROM[39834] <= 32'b00000000010000010000000100010011;
ROM[39835] <= 32'b00000000000000100111001110110111;
ROM[39836] <= 32'b11101011100000111000001110010011;
ROM[39837] <= 32'b00000000111000111000001110110011;
ROM[39838] <= 32'b00000000011100010010000000100011;
ROM[39839] <= 32'b00000000010000010000000100010011;
ROM[39840] <= 32'b00000000001100010010000000100011;
ROM[39841] <= 32'b00000000010000010000000100010011;
ROM[39842] <= 32'b00000000010000010010000000100011;
ROM[39843] <= 32'b00000000010000010000000100010011;
ROM[39844] <= 32'b00000000010100010010000000100011;
ROM[39845] <= 32'b00000000010000010000000100010011;
ROM[39846] <= 32'b00000000011000010010000000100011;
ROM[39847] <= 32'b00000000010000010000000100010011;
ROM[39848] <= 32'b00000001010000000000001110010011;
ROM[39849] <= 32'b00000000100000111000001110010011;
ROM[39850] <= 32'b01000000011100010000001110110011;
ROM[39851] <= 32'b00000000011100000000001000110011;
ROM[39852] <= 32'b00000000001000000000000110110011;
ROM[39853] <= 32'b10010111100111101010000011101111;
ROM[39854] <= 32'b00000000010000100010001110000011;
ROM[39855] <= 32'b00000000011100010010000000100011;
ROM[39856] <= 32'b00000000010000010000000100010011;
ROM[39857] <= 32'b00000000010000000000001110010011;
ROM[39858] <= 32'b00000000011100010010000000100011;
ROM[39859] <= 32'b00000000010000010000000100010011;
ROM[39860] <= 32'b00000000000000100111001110110111;
ROM[39861] <= 32'b11110001110000111000001110010011;
ROM[39862] <= 32'b00000000111000111000001110110011;
ROM[39863] <= 32'b00000000011100010010000000100011;
ROM[39864] <= 32'b00000000010000010000000100010011;
ROM[39865] <= 32'b00000000001100010010000000100011;
ROM[39866] <= 32'b00000000010000010000000100010011;
ROM[39867] <= 32'b00000000010000010010000000100011;
ROM[39868] <= 32'b00000000010000010000000100010011;
ROM[39869] <= 32'b00000000010100010010000000100011;
ROM[39870] <= 32'b00000000010000010000000100010011;
ROM[39871] <= 32'b00000000011000010010000000100011;
ROM[39872] <= 32'b00000000010000010000000100010011;
ROM[39873] <= 32'b00000001010000000000001110010011;
ROM[39874] <= 32'b00000000100000111000001110010011;
ROM[39875] <= 32'b01000000011100010000001110110011;
ROM[39876] <= 32'b00000000011100000000001000110011;
ROM[39877] <= 32'b00000000001000000000000110110011;
ROM[39878] <= 32'b10010001010111101010000011101111;
ROM[39879] <= 32'b00000000010000000000001110010011;
ROM[39880] <= 32'b00000000011100010010000000100011;
ROM[39881] <= 32'b00000000010000010000000100010011;
ROM[39882] <= 32'b11111111110000010000000100010011;
ROM[39883] <= 32'b00000000000000010010001110000011;
ROM[39884] <= 32'b11111111110000010000000100010011;
ROM[39885] <= 32'b00000000000000010010010000000011;
ROM[39886] <= 32'b00000000011101000000001110110011;
ROM[39887] <= 32'b00000000011100010010000000100011;
ROM[39888] <= 32'b00000000010000010000000100010011;
ROM[39889] <= 32'b00000000100000100010001110000011;
ROM[39890] <= 32'b00000000011100010010000000100011;
ROM[39891] <= 32'b00000000010000010000000100010011;
ROM[39892] <= 32'b00000000010000000000001110010011;
ROM[39893] <= 32'b00000000011100010010000000100011;
ROM[39894] <= 32'b00000000010000010000000100010011;
ROM[39895] <= 32'b00000000000000100111001110110111;
ROM[39896] <= 32'b11111010100000111000001110010011;
ROM[39897] <= 32'b00000000111000111000001110110011;
ROM[39898] <= 32'b00000000011100010010000000100011;
ROM[39899] <= 32'b00000000010000010000000100010011;
ROM[39900] <= 32'b00000000001100010010000000100011;
ROM[39901] <= 32'b00000000010000010000000100010011;
ROM[39902] <= 32'b00000000010000010010000000100011;
ROM[39903] <= 32'b00000000010000010000000100010011;
ROM[39904] <= 32'b00000000010100010010000000100011;
ROM[39905] <= 32'b00000000010000010000000100010011;
ROM[39906] <= 32'b00000000011000010010000000100011;
ROM[39907] <= 32'b00000000010000010000000100010011;
ROM[39908] <= 32'b00000001010000000000001110010011;
ROM[39909] <= 32'b00000000100000111000001110010011;
ROM[39910] <= 32'b01000000011100010000001110110011;
ROM[39911] <= 32'b00000000011100000000001000110011;
ROM[39912] <= 32'b00000000001000000000000110110011;
ROM[39913] <= 32'b10001000100111101010000011101111;
ROM[39914] <= 32'b00000000010000000000001110010011;
ROM[39915] <= 32'b00000000011100010010000000100011;
ROM[39916] <= 32'b00000000010000010000000100010011;
ROM[39917] <= 32'b11111111110000010000000100010011;
ROM[39918] <= 32'b00000000000000010010001110000011;
ROM[39919] <= 32'b11111111110000010000000100010011;
ROM[39920] <= 32'b00000000000000010010010000000011;
ROM[39921] <= 32'b00000000011101000000001110110011;
ROM[39922] <= 32'b00000000011100010010000000100011;
ROM[39923] <= 32'b00000000010000010000000100010011;
ROM[39924] <= 32'b00000000000000100111001110110111;
ROM[39925] <= 32'b00000001110000111000001110010011;
ROM[39926] <= 32'b00000000111000111000001110110011;
ROM[39927] <= 32'b00000000011100010010000000100011;
ROM[39928] <= 32'b00000000010000010000000100010011;
ROM[39929] <= 32'b00000000001100010010000000100011;
ROM[39930] <= 32'b00000000010000010000000100010011;
ROM[39931] <= 32'b00000000010000010010000000100011;
ROM[39932] <= 32'b00000000010000010000000100010011;
ROM[39933] <= 32'b00000000010100010010000000100011;
ROM[39934] <= 32'b00000000010000010000000100010011;
ROM[39935] <= 32'b00000000011000010010000000100011;
ROM[39936] <= 32'b00000000010000010000000100010011;
ROM[39937] <= 32'b00000001010000000000001110010011;
ROM[39938] <= 32'b00000001000000111000001110010011;
ROM[39939] <= 32'b01000000011100010000001110110011;
ROM[39940] <= 32'b00000000011100000000001000110011;
ROM[39941] <= 32'b00000000001000000000000110110011;
ROM[39942] <= 32'b10111100110011111000000011101111;
ROM[39943] <= 32'b11111111110000010000000100010011;
ROM[39944] <= 32'b00000000000000010010001110000011;
ROM[39945] <= 32'b00000000011101100010000000100011;
ROM[39946] <= 32'b00000000010100010010000000100011;
ROM[39947] <= 32'b00000000010000010000000100010011;
ROM[39948] <= 32'b00000000010000100010001110000011;
ROM[39949] <= 32'b00000000011100010010000000100011;
ROM[39950] <= 32'b00000000010000010000000100010011;
ROM[39951] <= 32'b00000000100000100010001110000011;
ROM[39952] <= 32'b00000000011100010010000000100011;
ROM[39953] <= 32'b00000000010000010000000100010011;
ROM[39954] <= 32'b00000000000000000000001110010011;
ROM[39955] <= 32'b00000000011100010010000000100011;
ROM[39956] <= 32'b00000000010000010000000100010011;
ROM[39957] <= 32'b00000000000000100111001110110111;
ROM[39958] <= 32'b00001010000000111000001110010011;
ROM[39959] <= 32'b00000000111000111000001110110011;
ROM[39960] <= 32'b00000000011100010010000000100011;
ROM[39961] <= 32'b00000000010000010000000100010011;
ROM[39962] <= 32'b00000000001100010010000000100011;
ROM[39963] <= 32'b00000000010000010000000100010011;
ROM[39964] <= 32'b00000000010000010010000000100011;
ROM[39965] <= 32'b00000000010000010000000100010011;
ROM[39966] <= 32'b00000000010100010010000000100011;
ROM[39967] <= 32'b00000000010000010000000100010011;
ROM[39968] <= 32'b00000000011000010010000000100011;
ROM[39969] <= 32'b00000000010000010000000100010011;
ROM[39970] <= 32'b00000001010000000000001110010011;
ROM[39971] <= 32'b00000001000000111000001110010011;
ROM[39972] <= 32'b01000000011100010000001110110011;
ROM[39973] <= 32'b00000000011100000000001000110011;
ROM[39974] <= 32'b00000000001000000000000110110011;
ROM[39975] <= 32'b10000111110011111111000011101111;
ROM[39976] <= 32'b11111111110000010000000100010011;
ROM[39977] <= 32'b00000000000000010010001110000011;
ROM[39978] <= 32'b00000000011101100010000000100011;
ROM[39979] <= 32'b00000000000000000000001110010011;
ROM[39980] <= 32'b00000000011100010010000000100011;
ROM[39981] <= 32'b00000000010000010000000100010011;
ROM[39982] <= 32'b00000001010000000000001110010011;
ROM[39983] <= 32'b01000000011100011000001110110011;
ROM[39984] <= 32'b00000000000000111010000010000011;
ROM[39985] <= 32'b11111111110000010000000100010011;
ROM[39986] <= 32'b00000000000000010010001110000011;
ROM[39987] <= 32'b00000000011100100010000000100011;
ROM[39988] <= 32'b00000000010000100000000100010011;
ROM[39989] <= 32'b00000001010000000000001110010011;
ROM[39990] <= 32'b01000000011100011000001110110011;
ROM[39991] <= 32'b00000000010000111010000110000011;
ROM[39992] <= 32'b00000000100000111010001000000011;
ROM[39993] <= 32'b00000000110000111010001010000011;
ROM[39994] <= 32'b00000001000000111010001100000011;
ROM[39995] <= 32'b00000000000000001000000011100111;
ROM[39996] <= 32'b00000000000000010010000000100011;
ROM[39997] <= 32'b00000000010000010000000100010011;
ROM[39998] <= 32'b00000000000000010010000000100011;
ROM[39999] <= 32'b00000000010000010000000100010011;
ROM[40000] <= 32'b00000000000000100010001110000011;
ROM[40001] <= 32'b00000000011100010010000000100011;
ROM[40002] <= 32'b00000000010000010000000100010011;
ROM[40003] <= 32'b11111111110000010000000100010011;
ROM[40004] <= 32'b00000000000000010010001110000011;
ROM[40005] <= 32'b00000000000000111000001010010011;
ROM[40006] <= 32'b00000001011000000000001110010011;
ROM[40007] <= 32'b00000000011100010010000000100011;
ROM[40008] <= 32'b00000000010000010000000100010011;
ROM[40009] <= 32'b00000000000000000000001110010011;
ROM[40010] <= 32'b00000000011100010010000000100011;
ROM[40011] <= 32'b00000000010000010000000100010011;
ROM[40012] <= 32'b00000000000000100111001110110111;
ROM[40013] <= 32'b00010111110000111000001110010011;
ROM[40014] <= 32'b00000000111000111000001110110011;
ROM[40015] <= 32'b00000000011100010010000000100011;
ROM[40016] <= 32'b00000000010000010000000100010011;
ROM[40017] <= 32'b00000000001100010010000000100011;
ROM[40018] <= 32'b00000000010000010000000100010011;
ROM[40019] <= 32'b00000000010000010010000000100011;
ROM[40020] <= 32'b00000000010000010000000100010011;
ROM[40021] <= 32'b00000000010100010010000000100011;
ROM[40022] <= 32'b00000000010000010000000100010011;
ROM[40023] <= 32'b00000000011000010010000000100011;
ROM[40024] <= 32'b00000000010000010000000100010011;
ROM[40025] <= 32'b00000001010000000000001110010011;
ROM[40026] <= 32'b00000000100000111000001110010011;
ROM[40027] <= 32'b01000000011100010000001110110011;
ROM[40028] <= 32'b00000000011100000000001000110011;
ROM[40029] <= 32'b00000000001000000000000110110011;
ROM[40030] <= 32'b10101000100111101110000011101111;
ROM[40031] <= 32'b11111111110000010000000100010011;
ROM[40032] <= 32'b00000000000000010010001110000011;
ROM[40033] <= 32'b00000000011101100010000000100011;
ROM[40034] <= 32'b00000000011100000000001110010011;
ROM[40035] <= 32'b00000000011100010010000000100011;
ROM[40036] <= 32'b00000000010000010000000100010011;
ROM[40037] <= 32'b00000000000000100111001110110111;
ROM[40038] <= 32'b00011110000000111000001110010011;
ROM[40039] <= 32'b00000000111000111000001110110011;
ROM[40040] <= 32'b00000000011100010010000000100011;
ROM[40041] <= 32'b00000000010000010000000100010011;
ROM[40042] <= 32'b00000000001100010010000000100011;
ROM[40043] <= 32'b00000000010000010000000100010011;
ROM[40044] <= 32'b00000000010000010010000000100011;
ROM[40045] <= 32'b00000000010000010000000100010011;
ROM[40046] <= 32'b00000000010100010010000000100011;
ROM[40047] <= 32'b00000000010000010000000100010011;
ROM[40048] <= 32'b00000000011000010010000000100011;
ROM[40049] <= 32'b00000000010000010000000100010011;
ROM[40050] <= 32'b00000001010000000000001110010011;
ROM[40051] <= 32'b00000000010000111000001110010011;
ROM[40052] <= 32'b01000000011100010000001110110011;
ROM[40053] <= 32'b00000000011100000000001000110011;
ROM[40054] <= 32'b00000000001000000000000110110011;
ROM[40055] <= 32'b01010110000000000010000011101111;
ROM[40056] <= 32'b00000100110000000000001110010011;
ROM[40057] <= 32'b00000000011100010010000000100011;
ROM[40058] <= 32'b00000000010000010000000100010011;
ROM[40059] <= 32'b00000000000000100111001110110111;
ROM[40060] <= 32'b00100011100000111000001110010011;
ROM[40061] <= 32'b00000000111000111000001110110011;
ROM[40062] <= 32'b00000000011100010010000000100011;
ROM[40063] <= 32'b00000000010000010000000100010011;
ROM[40064] <= 32'b00000000001100010010000000100011;
ROM[40065] <= 32'b00000000010000010000000100010011;
ROM[40066] <= 32'b00000000010000010010000000100011;
ROM[40067] <= 32'b00000000010000010000000100010011;
ROM[40068] <= 32'b00000000010100010010000000100011;
ROM[40069] <= 32'b00000000010000010000000100010011;
ROM[40070] <= 32'b00000000011000010010000000100011;
ROM[40071] <= 32'b00000000010000010000000100010011;
ROM[40072] <= 32'b00000001010000000000001110010011;
ROM[40073] <= 32'b00000000100000111000001110010011;
ROM[40074] <= 32'b01000000011100010000001110110011;
ROM[40075] <= 32'b00000000011100000000001000110011;
ROM[40076] <= 32'b00000000001000000000000110110011;
ROM[40077] <= 32'b00010111100100000010000011101111;
ROM[40078] <= 32'b00000110010100000000001110010011;
ROM[40079] <= 32'b00000000011100010010000000100011;
ROM[40080] <= 32'b00000000010000010000000100010011;
ROM[40081] <= 32'b00000000000000100111001110110111;
ROM[40082] <= 32'b00101001000000111000001110010011;
ROM[40083] <= 32'b00000000111000111000001110110011;
ROM[40084] <= 32'b00000000011100010010000000100011;
ROM[40085] <= 32'b00000000010000010000000100010011;
ROM[40086] <= 32'b00000000001100010010000000100011;
ROM[40087] <= 32'b00000000010000010000000100010011;
ROM[40088] <= 32'b00000000010000010010000000100011;
ROM[40089] <= 32'b00000000010000010000000100010011;
ROM[40090] <= 32'b00000000010100010010000000100011;
ROM[40091] <= 32'b00000000010000010000000100010011;
ROM[40092] <= 32'b00000000011000010010000000100011;
ROM[40093] <= 32'b00000000010000010000000100010011;
ROM[40094] <= 32'b00000001010000000000001110010011;
ROM[40095] <= 32'b00000000100000111000001110010011;
ROM[40096] <= 32'b01000000011100010000001110110011;
ROM[40097] <= 32'b00000000011100000000001000110011;
ROM[40098] <= 32'b00000000001000000000000110110011;
ROM[40099] <= 32'b00010010000100000010000011101111;
ROM[40100] <= 32'b00000111011000000000001110010011;
ROM[40101] <= 32'b00000000011100010010000000100011;
ROM[40102] <= 32'b00000000010000010000000100010011;
ROM[40103] <= 32'b00000000000000100111001110110111;
ROM[40104] <= 32'b00101110100000111000001110010011;
ROM[40105] <= 32'b00000000111000111000001110110011;
ROM[40106] <= 32'b00000000011100010010000000100011;
ROM[40107] <= 32'b00000000010000010000000100010011;
ROM[40108] <= 32'b00000000001100010010000000100011;
ROM[40109] <= 32'b00000000010000010000000100010011;
ROM[40110] <= 32'b00000000010000010010000000100011;
ROM[40111] <= 32'b00000000010000010000000100010011;
ROM[40112] <= 32'b00000000010100010010000000100011;
ROM[40113] <= 32'b00000000010000010000000100010011;
ROM[40114] <= 32'b00000000011000010010000000100011;
ROM[40115] <= 32'b00000000010000010000000100010011;
ROM[40116] <= 32'b00000001010000000000001110010011;
ROM[40117] <= 32'b00000000100000111000001110010011;
ROM[40118] <= 32'b01000000011100010000001110110011;
ROM[40119] <= 32'b00000000011100000000001000110011;
ROM[40120] <= 32'b00000000001000000000000110110011;
ROM[40121] <= 32'b00001100100100000010000011101111;
ROM[40122] <= 32'b00000110010100000000001110010011;
ROM[40123] <= 32'b00000000011100010010000000100011;
ROM[40124] <= 32'b00000000010000010000000100010011;
ROM[40125] <= 32'b00000000000000100111001110110111;
ROM[40126] <= 32'b00110100000000111000001110010011;
ROM[40127] <= 32'b00000000111000111000001110110011;
ROM[40128] <= 32'b00000000011100010010000000100011;
ROM[40129] <= 32'b00000000010000010000000100010011;
ROM[40130] <= 32'b00000000001100010010000000100011;
ROM[40131] <= 32'b00000000010000010000000100010011;
ROM[40132] <= 32'b00000000010000010010000000100011;
ROM[40133] <= 32'b00000000010000010000000100010011;
ROM[40134] <= 32'b00000000010100010010000000100011;
ROM[40135] <= 32'b00000000010000010000000100010011;
ROM[40136] <= 32'b00000000011000010010000000100011;
ROM[40137] <= 32'b00000000010000010000000100010011;
ROM[40138] <= 32'b00000001010000000000001110010011;
ROM[40139] <= 32'b00000000100000111000001110010011;
ROM[40140] <= 32'b01000000011100010000001110110011;
ROM[40141] <= 32'b00000000011100000000001000110011;
ROM[40142] <= 32'b00000000001000000000000110110011;
ROM[40143] <= 32'b00000111000100000010000011101111;
ROM[40144] <= 32'b00000110110000000000001110010011;
ROM[40145] <= 32'b00000000011100010010000000100011;
ROM[40146] <= 32'b00000000010000010000000100010011;
ROM[40147] <= 32'b00000000000000100111001110110111;
ROM[40148] <= 32'b00111001100000111000001110010011;
ROM[40149] <= 32'b00000000111000111000001110110011;
ROM[40150] <= 32'b00000000011100010010000000100011;
ROM[40151] <= 32'b00000000010000010000000100010011;
ROM[40152] <= 32'b00000000001100010010000000100011;
ROM[40153] <= 32'b00000000010000010000000100010011;
ROM[40154] <= 32'b00000000010000010010000000100011;
ROM[40155] <= 32'b00000000010000010000000100010011;
ROM[40156] <= 32'b00000000010100010010000000100011;
ROM[40157] <= 32'b00000000010000010000000100010011;
ROM[40158] <= 32'b00000000011000010010000000100011;
ROM[40159] <= 32'b00000000010000010000000100010011;
ROM[40160] <= 32'b00000001010000000000001110010011;
ROM[40161] <= 32'b00000000100000111000001110010011;
ROM[40162] <= 32'b01000000011100010000001110110011;
ROM[40163] <= 32'b00000000011100000000001000110011;
ROM[40164] <= 32'b00000000001000000000000110110011;
ROM[40165] <= 32'b00000001100100000010000011101111;
ROM[40166] <= 32'b00000011101000000000001110010011;
ROM[40167] <= 32'b00000000011100010010000000100011;
ROM[40168] <= 32'b00000000010000010000000100010011;
ROM[40169] <= 32'b00000000000000100111001110110111;
ROM[40170] <= 32'b00111111000000111000001110010011;
ROM[40171] <= 32'b00000000111000111000001110110011;
ROM[40172] <= 32'b00000000011100010010000000100011;
ROM[40173] <= 32'b00000000010000010000000100010011;
ROM[40174] <= 32'b00000000001100010010000000100011;
ROM[40175] <= 32'b00000000010000010000000100010011;
ROM[40176] <= 32'b00000000010000010010000000100011;
ROM[40177] <= 32'b00000000010000010000000100010011;
ROM[40178] <= 32'b00000000010100010010000000100011;
ROM[40179] <= 32'b00000000010000010000000100010011;
ROM[40180] <= 32'b00000000011000010010000000100011;
ROM[40181] <= 32'b00000000010000010000000100010011;
ROM[40182] <= 32'b00000001010000000000001110010011;
ROM[40183] <= 32'b00000000100000111000001110010011;
ROM[40184] <= 32'b01000000011100010000001110110011;
ROM[40185] <= 32'b00000000011100000000001000110011;
ROM[40186] <= 32'b00000000001000000000000110110011;
ROM[40187] <= 32'b01111100000000000010000011101111;
ROM[40188] <= 32'b00000010000000000000001110010011;
ROM[40189] <= 32'b00000000011100010010000000100011;
ROM[40190] <= 32'b00000000010000010000000100010011;
ROM[40191] <= 32'b00000000000000100111001110110111;
ROM[40192] <= 32'b01000100100000111000001110010011;
ROM[40193] <= 32'b00000000111000111000001110110011;
ROM[40194] <= 32'b00000000011100010010000000100011;
ROM[40195] <= 32'b00000000010000010000000100010011;
ROM[40196] <= 32'b00000000001100010010000000100011;
ROM[40197] <= 32'b00000000010000010000000100010011;
ROM[40198] <= 32'b00000000010000010010000000100011;
ROM[40199] <= 32'b00000000010000010000000100010011;
ROM[40200] <= 32'b00000000010100010010000000100011;
ROM[40201] <= 32'b00000000010000010000000100010011;
ROM[40202] <= 32'b00000000011000010010000000100011;
ROM[40203] <= 32'b00000000010000010000000100010011;
ROM[40204] <= 32'b00000001010000000000001110010011;
ROM[40205] <= 32'b00000000100000111000001110010011;
ROM[40206] <= 32'b01000000011100010000001110110011;
ROM[40207] <= 32'b00000000011100000000001000110011;
ROM[40208] <= 32'b00000000001000000000000110110011;
ROM[40209] <= 32'b01110110100000000010000011101111;
ROM[40210] <= 32'b11111111110000010000000100010011;
ROM[40211] <= 32'b00000000000000010010001110000011;
ROM[40212] <= 32'b00000000011100011010001000100011;
ROM[40213] <= 32'b00000000010000011010001110000011;
ROM[40214] <= 32'b00000000011100010010000000100011;
ROM[40215] <= 32'b00000000010000010000000100010011;
ROM[40216] <= 32'b00000000000000100111001110110111;
ROM[40217] <= 32'b01001010110000111000001110010011;
ROM[40218] <= 32'b00000000111000111000001110110011;
ROM[40219] <= 32'b00000000011100010010000000100011;
ROM[40220] <= 32'b00000000010000010000000100010011;
ROM[40221] <= 32'b00000000001100010010000000100011;
ROM[40222] <= 32'b00000000010000010000000100010011;
ROM[40223] <= 32'b00000000010000010010000000100011;
ROM[40224] <= 32'b00000000010000010000000100010011;
ROM[40225] <= 32'b00000000010100010010000000100011;
ROM[40226] <= 32'b00000000010000010000000100010011;
ROM[40227] <= 32'b00000000011000010010000000100011;
ROM[40228] <= 32'b00000000010000010000000100010011;
ROM[40229] <= 32'b00000001010000000000001110010011;
ROM[40230] <= 32'b00000000010000111000001110010011;
ROM[40231] <= 32'b01000000011100010000001110110011;
ROM[40232] <= 32'b00000000011100000000001000110011;
ROM[40233] <= 32'b00000000001000000000000110110011;
ROM[40234] <= 32'b10101100000111101111000011101111;
ROM[40235] <= 32'b11111111110000010000000100010011;
ROM[40236] <= 32'b00000000000000010010001110000011;
ROM[40237] <= 32'b00000000011101100010000000100011;
ROM[40238] <= 32'b00000000010000011010001110000011;
ROM[40239] <= 32'b00000000011100010010000000100011;
ROM[40240] <= 32'b00000000010000010000000100010011;
ROM[40241] <= 32'b00000000000000100111001110110111;
ROM[40242] <= 32'b01010001000000111000001110010011;
ROM[40243] <= 32'b00000000111000111000001110110011;
ROM[40244] <= 32'b00000000011100010010000000100011;
ROM[40245] <= 32'b00000000010000010000000100010011;
ROM[40246] <= 32'b00000000001100010010000000100011;
ROM[40247] <= 32'b00000000010000010000000100010011;
ROM[40248] <= 32'b00000000010000010010000000100011;
ROM[40249] <= 32'b00000000010000010000000100010011;
ROM[40250] <= 32'b00000000010100010010000000100011;
ROM[40251] <= 32'b00000000010000010000000100010011;
ROM[40252] <= 32'b00000000011000010010000000100011;
ROM[40253] <= 32'b00000000010000010000000100010011;
ROM[40254] <= 32'b00000001010000000000001110010011;
ROM[40255] <= 32'b00000000010000111000001110010011;
ROM[40256] <= 32'b01000000011100010000001110110011;
ROM[40257] <= 32'b00000000011100000000001000110011;
ROM[40258] <= 32'b00000000001000000000000110110011;
ROM[40259] <= 32'b00000000010100000011000011101111;
ROM[40260] <= 32'b11111111110000010000000100010011;
ROM[40261] <= 32'b00000000000000010010001110000011;
ROM[40262] <= 32'b00000000011101100010000000100011;
ROM[40263] <= 32'b00000000110100101000010000110011;
ROM[40264] <= 32'b00000000000001000010001110000011;
ROM[40265] <= 32'b00000000011100010010000000100011;
ROM[40266] <= 32'b00000000010000010000000100010011;
ROM[40267] <= 32'b00000000000000100111001110110111;
ROM[40268] <= 32'b01010111100000111000001110010011;
ROM[40269] <= 32'b00000000111000111000001110110011;
ROM[40270] <= 32'b00000000011100010010000000100011;
ROM[40271] <= 32'b00000000010000010000000100010011;
ROM[40272] <= 32'b00000000001100010010000000100011;
ROM[40273] <= 32'b00000000010000010000000100010011;
ROM[40274] <= 32'b00000000010000010010000000100011;
ROM[40275] <= 32'b00000000010000010000000100010011;
ROM[40276] <= 32'b00000000010100010010000000100011;
ROM[40277] <= 32'b00000000010000010000000100010011;
ROM[40278] <= 32'b00000000011000010010000000100011;
ROM[40279] <= 32'b00000000010000010000000100010011;
ROM[40280] <= 32'b00000001010000000000001110010011;
ROM[40281] <= 32'b00000000010000111000001110010011;
ROM[40282] <= 32'b01000000011100010000001110110011;
ROM[40283] <= 32'b00000000011100000000001000110011;
ROM[40284] <= 32'b00000000001000000000000110110011;
ROM[40285] <= 32'b11100111000011111100000011101111;
ROM[40286] <= 32'b00000000000000100111001110110111;
ROM[40287] <= 32'b01011100010000111000001110010011;
ROM[40288] <= 32'b00000000111000111000001110110011;
ROM[40289] <= 32'b00000000011100010010000000100011;
ROM[40290] <= 32'b00000000010000010000000100010011;
ROM[40291] <= 32'b00000000001100010010000000100011;
ROM[40292] <= 32'b00000000010000010000000100010011;
ROM[40293] <= 32'b00000000010000010010000000100011;
ROM[40294] <= 32'b00000000010000010000000100010011;
ROM[40295] <= 32'b00000000010100010010000000100011;
ROM[40296] <= 32'b00000000010000010000000100010011;
ROM[40297] <= 32'b00000000011000010010000000100011;
ROM[40298] <= 32'b00000000010000010000000100010011;
ROM[40299] <= 32'b00000001010000000000001110010011;
ROM[40300] <= 32'b00000000010000111000001110010011;
ROM[40301] <= 32'b01000000011100010000001110110011;
ROM[40302] <= 32'b00000000011100000000001000110011;
ROM[40303] <= 32'b00000000001000000000000110110011;
ROM[40304] <= 32'b10111100000111101111000011101111;
ROM[40305] <= 32'b11111111110000010000000100010011;
ROM[40306] <= 32'b00000000000000010010001110000011;
ROM[40307] <= 32'b00000000011101100010000000100011;
ROM[40308] <= 32'b00000001011000000000001110010011;
ROM[40309] <= 32'b00000000011100010010000000100011;
ROM[40310] <= 32'b00000000010000010000000100010011;
ROM[40311] <= 32'b00000001100100000000001110010011;
ROM[40312] <= 32'b00000000011100010010000000100011;
ROM[40313] <= 32'b00000000010000010000000100010011;
ROM[40314] <= 32'b00000000000000100111001110110111;
ROM[40315] <= 32'b01100011010000111000001110010011;
ROM[40316] <= 32'b00000000111000111000001110110011;
ROM[40317] <= 32'b00000000011100010010000000100011;
ROM[40318] <= 32'b00000000010000010000000100010011;
ROM[40319] <= 32'b00000000001100010010000000100011;
ROM[40320] <= 32'b00000000010000010000000100010011;
ROM[40321] <= 32'b00000000010000010010000000100011;
ROM[40322] <= 32'b00000000010000010000000100010011;
ROM[40323] <= 32'b00000000010100010010000000100011;
ROM[40324] <= 32'b00000000010000010000000100010011;
ROM[40325] <= 32'b00000000011000010010000000100011;
ROM[40326] <= 32'b00000000010000010000000100010011;
ROM[40327] <= 32'b00000001010000000000001110010011;
ROM[40328] <= 32'b00000000100000111000001110010011;
ROM[40329] <= 32'b01000000011100010000001110110011;
ROM[40330] <= 32'b00000000011100000000001000110011;
ROM[40331] <= 32'b00000000001000000000000110110011;
ROM[40332] <= 32'b11011101000011101110000011101111;
ROM[40333] <= 32'b11111111110000010000000100010011;
ROM[40334] <= 32'b00000000000000010010001110000011;
ROM[40335] <= 32'b00000000011101100010000000100011;
ROM[40336] <= 32'b00000000011100000000001110010011;
ROM[40337] <= 32'b00000000011100010010000000100011;
ROM[40338] <= 32'b00000000010000010000000100010011;
ROM[40339] <= 32'b00000000000000100111001110110111;
ROM[40340] <= 32'b01101001100000111000001110010011;
ROM[40341] <= 32'b00000000111000111000001110110011;
ROM[40342] <= 32'b00000000011100010010000000100011;
ROM[40343] <= 32'b00000000010000010000000100010011;
ROM[40344] <= 32'b00000000001100010010000000100011;
ROM[40345] <= 32'b00000000010000010000000100010011;
ROM[40346] <= 32'b00000000010000010010000000100011;
ROM[40347] <= 32'b00000000010000010000000100010011;
ROM[40348] <= 32'b00000000010100010010000000100011;
ROM[40349] <= 32'b00000000010000010000000100010011;
ROM[40350] <= 32'b00000000011000010010000000100011;
ROM[40351] <= 32'b00000000010000010000000100010011;
ROM[40352] <= 32'b00000001010000000000001110010011;
ROM[40353] <= 32'b00000000010000111000001110010011;
ROM[40354] <= 32'b01000000011100010000001110110011;
ROM[40355] <= 32'b00000000011100000000001000110011;
ROM[40356] <= 32'b00000000001000000000000110110011;
ROM[40357] <= 32'b00001010100000000010000011101111;
ROM[40358] <= 32'b00000101001100000000001110010011;
ROM[40359] <= 32'b00000000011100010010000000100011;
ROM[40360] <= 32'b00000000010000010000000100010011;
ROM[40361] <= 32'b00000000000000100111001110110111;
ROM[40362] <= 32'b01101111000000111000001110010011;
ROM[40363] <= 32'b00000000111000111000001110110011;
ROM[40364] <= 32'b00000000011100010010000000100011;
ROM[40365] <= 32'b00000000010000010000000100010011;
ROM[40366] <= 32'b00000000001100010010000000100011;
ROM[40367] <= 32'b00000000010000010000000100010011;
ROM[40368] <= 32'b00000000010000010010000000100011;
ROM[40369] <= 32'b00000000010000010000000100010011;
ROM[40370] <= 32'b00000000010100010010000000100011;
ROM[40371] <= 32'b00000000010000010000000100010011;
ROM[40372] <= 32'b00000000011000010010000000100011;
ROM[40373] <= 32'b00000000010000010000000100010011;
ROM[40374] <= 32'b00000001010000000000001110010011;
ROM[40375] <= 32'b00000000100000111000001110010011;
ROM[40376] <= 32'b01000000011100010000001110110011;
ROM[40377] <= 32'b00000000011100000000001000110011;
ROM[40378] <= 32'b00000000001000000000000110110011;
ROM[40379] <= 32'b01001100000000000010000011101111;
ROM[40380] <= 32'b00000110001100000000001110010011;
ROM[40381] <= 32'b00000000011100010010000000100011;
ROM[40382] <= 32'b00000000010000010000000100010011;
ROM[40383] <= 32'b00000000000000100111001110110111;
ROM[40384] <= 32'b01110100100000111000001110010011;
ROM[40385] <= 32'b00000000111000111000001110110011;
ROM[40386] <= 32'b00000000011100010010000000100011;
ROM[40387] <= 32'b00000000010000010000000100010011;
ROM[40388] <= 32'b00000000001100010010000000100011;
ROM[40389] <= 32'b00000000010000010000000100010011;
ROM[40390] <= 32'b00000000010000010010000000100011;
ROM[40391] <= 32'b00000000010000010000000100010011;
ROM[40392] <= 32'b00000000010100010010000000100011;
ROM[40393] <= 32'b00000000010000010000000100010011;
ROM[40394] <= 32'b00000000011000010010000000100011;
ROM[40395] <= 32'b00000000010000010000000100010011;
ROM[40396] <= 32'b00000001010000000000001110010011;
ROM[40397] <= 32'b00000000100000111000001110010011;
ROM[40398] <= 32'b01000000011100010000001110110011;
ROM[40399] <= 32'b00000000011100000000001000110011;
ROM[40400] <= 32'b00000000001000000000000110110011;
ROM[40401] <= 32'b01000110100000000010000011101111;
ROM[40402] <= 32'b00000110111100000000001110010011;
ROM[40403] <= 32'b00000000011100010010000000100011;
ROM[40404] <= 32'b00000000010000010000000100010011;
ROM[40405] <= 32'b00000000000000100111001110110111;
ROM[40406] <= 32'b01111010000000111000001110010011;
ROM[40407] <= 32'b00000000111000111000001110110011;
ROM[40408] <= 32'b00000000011100010010000000100011;
ROM[40409] <= 32'b00000000010000010000000100010011;
ROM[40410] <= 32'b00000000001100010010000000100011;
ROM[40411] <= 32'b00000000010000010000000100010011;
ROM[40412] <= 32'b00000000010000010010000000100011;
ROM[40413] <= 32'b00000000010000010000000100010011;
ROM[40414] <= 32'b00000000010100010010000000100011;
ROM[40415] <= 32'b00000000010000010000000100010011;
ROM[40416] <= 32'b00000000011000010010000000100011;
ROM[40417] <= 32'b00000000010000010000000100010011;
ROM[40418] <= 32'b00000001010000000000001110010011;
ROM[40419] <= 32'b00000000100000111000001110010011;
ROM[40420] <= 32'b01000000011100010000001110110011;
ROM[40421] <= 32'b00000000011100000000001000110011;
ROM[40422] <= 32'b00000000001000000000000110110011;
ROM[40423] <= 32'b01000001000000000010000011101111;
ROM[40424] <= 32'b00000111001000000000001110010011;
ROM[40425] <= 32'b00000000011100010010000000100011;
ROM[40426] <= 32'b00000000010000010000000100010011;
ROM[40427] <= 32'b00000000000000100111001110110111;
ROM[40428] <= 32'b01111111100000111000001110010011;
ROM[40429] <= 32'b00000000111000111000001110110011;
ROM[40430] <= 32'b00000000011100010010000000100011;
ROM[40431] <= 32'b00000000010000010000000100010011;
ROM[40432] <= 32'b00000000001100010010000000100011;
ROM[40433] <= 32'b00000000010000010000000100010011;
ROM[40434] <= 32'b00000000010000010010000000100011;
ROM[40435] <= 32'b00000000010000010000000100010011;
ROM[40436] <= 32'b00000000010100010010000000100011;
ROM[40437] <= 32'b00000000010000010000000100010011;
ROM[40438] <= 32'b00000000011000010010000000100011;
ROM[40439] <= 32'b00000000010000010000000100010011;
ROM[40440] <= 32'b00000001010000000000001110010011;
ROM[40441] <= 32'b00000000100000111000001110010011;
ROM[40442] <= 32'b01000000011100010000001110110011;
ROM[40443] <= 32'b00000000011100000000001000110011;
ROM[40444] <= 32'b00000000001000000000000110110011;
ROM[40445] <= 32'b00111011100000000010000011101111;
ROM[40446] <= 32'b00000110010100000000001110010011;
ROM[40447] <= 32'b00000000011100010010000000100011;
ROM[40448] <= 32'b00000000010000010000000100010011;
ROM[40449] <= 32'b00000000000000101000001110110111;
ROM[40450] <= 32'b10000101000000111000001110010011;
ROM[40451] <= 32'b00000000111000111000001110110011;
ROM[40452] <= 32'b00000000011100010010000000100011;
ROM[40453] <= 32'b00000000010000010000000100010011;
ROM[40454] <= 32'b00000000001100010010000000100011;
ROM[40455] <= 32'b00000000010000010000000100010011;
ROM[40456] <= 32'b00000000010000010010000000100011;
ROM[40457] <= 32'b00000000010000010000000100010011;
ROM[40458] <= 32'b00000000010100010010000000100011;
ROM[40459] <= 32'b00000000010000010000000100010011;
ROM[40460] <= 32'b00000000011000010010000000100011;
ROM[40461] <= 32'b00000000010000010000000100010011;
ROM[40462] <= 32'b00000001010000000000001110010011;
ROM[40463] <= 32'b00000000100000111000001110010011;
ROM[40464] <= 32'b01000000011100010000001110110011;
ROM[40465] <= 32'b00000000011100000000001000110011;
ROM[40466] <= 32'b00000000001000000000000110110011;
ROM[40467] <= 32'b00110110000000000010000011101111;
ROM[40468] <= 32'b00000011101000000000001110010011;
ROM[40469] <= 32'b00000000011100010010000000100011;
ROM[40470] <= 32'b00000000010000010000000100010011;
ROM[40471] <= 32'b00000000000000101000001110110111;
ROM[40472] <= 32'b10001010100000111000001110010011;
ROM[40473] <= 32'b00000000111000111000001110110011;
ROM[40474] <= 32'b00000000011100010010000000100011;
ROM[40475] <= 32'b00000000010000010000000100010011;
ROM[40476] <= 32'b00000000001100010010000000100011;
ROM[40477] <= 32'b00000000010000010000000100010011;
ROM[40478] <= 32'b00000000010000010010000000100011;
ROM[40479] <= 32'b00000000010000010000000100010011;
ROM[40480] <= 32'b00000000010100010010000000100011;
ROM[40481] <= 32'b00000000010000010000000100010011;
ROM[40482] <= 32'b00000000011000010010000000100011;
ROM[40483] <= 32'b00000000010000010000000100010011;
ROM[40484] <= 32'b00000001010000000000001110010011;
ROM[40485] <= 32'b00000000100000111000001110010011;
ROM[40486] <= 32'b01000000011100010000001110110011;
ROM[40487] <= 32'b00000000011100000000001000110011;
ROM[40488] <= 32'b00000000001000000000000110110011;
ROM[40489] <= 32'b00110000100000000010000011101111;
ROM[40490] <= 32'b00000010000000000000001110010011;
ROM[40491] <= 32'b00000000011100010010000000100011;
ROM[40492] <= 32'b00000000010000010000000100010011;
ROM[40493] <= 32'b00000000000000101000001110110111;
ROM[40494] <= 32'b10010000000000111000001110010011;
ROM[40495] <= 32'b00000000111000111000001110110011;
ROM[40496] <= 32'b00000000011100010010000000100011;
ROM[40497] <= 32'b00000000010000010000000100010011;
ROM[40498] <= 32'b00000000001100010010000000100011;
ROM[40499] <= 32'b00000000010000010000000100010011;
ROM[40500] <= 32'b00000000010000010010000000100011;
ROM[40501] <= 32'b00000000010000010000000100010011;
ROM[40502] <= 32'b00000000010100010010000000100011;
ROM[40503] <= 32'b00000000010000010000000100010011;
ROM[40504] <= 32'b00000000011000010010000000100011;
ROM[40505] <= 32'b00000000010000010000000100010011;
ROM[40506] <= 32'b00000001010000000000001110010011;
ROM[40507] <= 32'b00000000100000111000001110010011;
ROM[40508] <= 32'b01000000011100010000001110110011;
ROM[40509] <= 32'b00000000011100000000001000110011;
ROM[40510] <= 32'b00000000001000000000000110110011;
ROM[40511] <= 32'b00101011000000000010000011101111;
ROM[40512] <= 32'b11111111110000010000000100010011;
ROM[40513] <= 32'b00000000000000010010001110000011;
ROM[40514] <= 32'b00000000011100011010001000100011;
ROM[40515] <= 32'b00000000010000011010001110000011;
ROM[40516] <= 32'b00000000011100010010000000100011;
ROM[40517] <= 32'b00000000010000010000000100010011;
ROM[40518] <= 32'b00000000000000101000001110110111;
ROM[40519] <= 32'b10010110010000111000001110010011;
ROM[40520] <= 32'b00000000111000111000001110110011;
ROM[40521] <= 32'b00000000011100010010000000100011;
ROM[40522] <= 32'b00000000010000010000000100010011;
ROM[40523] <= 32'b00000000001100010010000000100011;
ROM[40524] <= 32'b00000000010000010000000100010011;
ROM[40525] <= 32'b00000000010000010010000000100011;
ROM[40526] <= 32'b00000000010000010000000100010011;
ROM[40527] <= 32'b00000000010100010010000000100011;
ROM[40528] <= 32'b00000000010000010000000100010011;
ROM[40529] <= 32'b00000000011000010010000000100011;
ROM[40530] <= 32'b00000000010000010000000100010011;
ROM[40531] <= 32'b00000001010000000000001110010011;
ROM[40532] <= 32'b00000000010000111000001110010011;
ROM[40533] <= 32'b01000000011100010000001110110011;
ROM[40534] <= 32'b00000000011100000000001000110011;
ROM[40535] <= 32'b00000000001000000000000110110011;
ROM[40536] <= 32'b11100000100011101111000011101111;
ROM[40537] <= 32'b11111111110000010000000100010011;
ROM[40538] <= 32'b00000000000000010010001110000011;
ROM[40539] <= 32'b00000000011101100010000000100011;
ROM[40540] <= 32'b00000000010000011010001110000011;
ROM[40541] <= 32'b00000000011100010010000000100011;
ROM[40542] <= 32'b00000000010000010000000100010011;
ROM[40543] <= 32'b00000000000000101000001110110111;
ROM[40544] <= 32'b10011100100000111000001110010011;
ROM[40545] <= 32'b00000000111000111000001110110011;
ROM[40546] <= 32'b00000000011100010010000000100011;
ROM[40547] <= 32'b00000000010000010000000100010011;
ROM[40548] <= 32'b00000000001100010010000000100011;
ROM[40549] <= 32'b00000000010000010000000100010011;
ROM[40550] <= 32'b00000000010000010010000000100011;
ROM[40551] <= 32'b00000000010000010000000100010011;
ROM[40552] <= 32'b00000000010100010010000000100011;
ROM[40553] <= 32'b00000000010000010000000100010011;
ROM[40554] <= 32'b00000000011000010010000000100011;
ROM[40555] <= 32'b00000000010000010000000100010011;
ROM[40556] <= 32'b00000001010000000000001110010011;
ROM[40557] <= 32'b00000000010000111000001110010011;
ROM[40558] <= 32'b01000000011100010000001110110011;
ROM[40559] <= 32'b00000000011100000000001000110011;
ROM[40560] <= 32'b00000000001000000000000110110011;
ROM[40561] <= 32'b00110100110000000011000011101111;
ROM[40562] <= 32'b11111111110000010000000100010011;
ROM[40563] <= 32'b00000000000000010010001110000011;
ROM[40564] <= 32'b00000000011101100010000000100011;
ROM[40565] <= 32'b00000000110100101000010000110011;
ROM[40566] <= 32'b00000000000001000010001110000011;
ROM[40567] <= 32'b00000000011100010010000000100011;
ROM[40568] <= 32'b00000000010000010000000100010011;
ROM[40569] <= 32'b00000000000000101000001110110111;
ROM[40570] <= 32'b10100011000000111000001110010011;
ROM[40571] <= 32'b00000000111000111000001110110011;
ROM[40572] <= 32'b00000000011100010010000000100011;
ROM[40573] <= 32'b00000000010000010000000100010011;
ROM[40574] <= 32'b00000000001100010010000000100011;
ROM[40575] <= 32'b00000000010000010000000100010011;
ROM[40576] <= 32'b00000000010000010010000000100011;
ROM[40577] <= 32'b00000000010000010000000100010011;
ROM[40578] <= 32'b00000000010100010010000000100011;
ROM[40579] <= 32'b00000000010000010000000100010011;
ROM[40580] <= 32'b00000000011000010010000000100011;
ROM[40581] <= 32'b00000000010000010000000100010011;
ROM[40582] <= 32'b00000001010000000000001110010011;
ROM[40583] <= 32'b00000000010000111000001110010011;
ROM[40584] <= 32'b01000000011100010000001110110011;
ROM[40585] <= 32'b00000000011100000000001000110011;
ROM[40586] <= 32'b00000000001000000000000110110011;
ROM[40587] <= 32'b10010101100011111100000011101111;
ROM[40588] <= 32'b00000000000000101000001110110111;
ROM[40589] <= 32'b10100111110000111000001110010011;
ROM[40590] <= 32'b00000000111000111000001110110011;
ROM[40591] <= 32'b00000000011100010010000000100011;
ROM[40592] <= 32'b00000000010000010000000100010011;
ROM[40593] <= 32'b00000000001100010010000000100011;
ROM[40594] <= 32'b00000000010000010000000100010011;
ROM[40595] <= 32'b00000000010000010010000000100011;
ROM[40596] <= 32'b00000000010000010000000100010011;
ROM[40597] <= 32'b00000000010100010010000000100011;
ROM[40598] <= 32'b00000000010000010000000100010011;
ROM[40599] <= 32'b00000000011000010010000000100011;
ROM[40600] <= 32'b00000000010000010000000100010011;
ROM[40601] <= 32'b00000001010000000000001110010011;
ROM[40602] <= 32'b00000000010000111000001110010011;
ROM[40603] <= 32'b01000000011100010000001110110011;
ROM[40604] <= 32'b00000000011100000000001000110011;
ROM[40605] <= 32'b00000000001000000000000110110011;
ROM[40606] <= 32'b11110000100011101111000011101111;
ROM[40607] <= 32'b11111111110000010000000100010011;
ROM[40608] <= 32'b00000000000000010010001110000011;
ROM[40609] <= 32'b00000000011101100010000000100011;
ROM[40610] <= 32'b00000001011000000000001110010011;
ROM[40611] <= 32'b00000000011100010010000000100011;
ROM[40612] <= 32'b00000000010000010000000100010011;
ROM[40613] <= 32'b00000011010000000000001110010011;
ROM[40614] <= 32'b00000000011100010010000000100011;
ROM[40615] <= 32'b00000000010000010000000100010011;
ROM[40616] <= 32'b00000000000000101000001110110111;
ROM[40617] <= 32'b10101110110000111000001110010011;
ROM[40618] <= 32'b00000000111000111000001110110011;
ROM[40619] <= 32'b00000000011100010010000000100011;
ROM[40620] <= 32'b00000000010000010000000100010011;
ROM[40621] <= 32'b00000000001100010010000000100011;
ROM[40622] <= 32'b00000000010000010000000100010011;
ROM[40623] <= 32'b00000000010000010010000000100011;
ROM[40624] <= 32'b00000000010000010000000100010011;
ROM[40625] <= 32'b00000000010100010010000000100011;
ROM[40626] <= 32'b00000000010000010000000100010011;
ROM[40627] <= 32'b00000000011000010010000000100011;
ROM[40628] <= 32'b00000000010000010000000100010011;
ROM[40629] <= 32'b00000001010000000000001110010011;
ROM[40630] <= 32'b00000000100000111000001110010011;
ROM[40631] <= 32'b01000000011100010000001110110011;
ROM[40632] <= 32'b00000000011100000000001000110011;
ROM[40633] <= 32'b00000000001000000000000110110011;
ROM[40634] <= 32'b10010001100011101110000011101111;
ROM[40635] <= 32'b11111111110000010000000100010011;
ROM[40636] <= 32'b00000000000000010010001110000011;
ROM[40637] <= 32'b00000000011101100010000000100011;
ROM[40638] <= 32'b00000000100000000000001110010011;
ROM[40639] <= 32'b00000000011100010010000000100011;
ROM[40640] <= 32'b00000000010000010000000100010011;
ROM[40641] <= 32'b00000000000000101000001110110111;
ROM[40642] <= 32'b10110101000000111000001110010011;
ROM[40643] <= 32'b00000000111000111000001110110011;
ROM[40644] <= 32'b00000000011100010010000000100011;
ROM[40645] <= 32'b00000000010000010000000100010011;
ROM[40646] <= 32'b00000000001100010010000000100011;
ROM[40647] <= 32'b00000000010000010000000100010011;
ROM[40648] <= 32'b00000000010000010010000000100011;
ROM[40649] <= 32'b00000000010000010000000100010011;
ROM[40650] <= 32'b00000000010100010010000000100011;
ROM[40651] <= 32'b00000000010000010000000100010011;
ROM[40652] <= 32'b00000000011000010010000000100011;
ROM[40653] <= 32'b00000000010000010000000100010011;
ROM[40654] <= 32'b00000001010000000000001110010011;
ROM[40655] <= 32'b00000000010000111000001110010011;
ROM[40656] <= 32'b01000000011100010000001110110011;
ROM[40657] <= 32'b00000000011100000000001000110011;
ROM[40658] <= 32'b00000000001000000000000110110011;
ROM[40659] <= 32'b00111111000100000001000011101111;
ROM[40660] <= 32'b00000100110000000000001110010011;
ROM[40661] <= 32'b00000000011100010010000000100011;
ROM[40662] <= 32'b00000000010000010000000100010011;
ROM[40663] <= 32'b00000000000000101000001110110111;
ROM[40664] <= 32'b10111010100000111000001110010011;
ROM[40665] <= 32'b00000000111000111000001110110011;
ROM[40666] <= 32'b00000000011100010010000000100011;
ROM[40667] <= 32'b00000000010000010000000100010011;
ROM[40668] <= 32'b00000000001100010010000000100011;
ROM[40669] <= 32'b00000000010000010000000100010011;
ROM[40670] <= 32'b00000000010000010010000000100011;
ROM[40671] <= 32'b00000000010000010000000100010011;
ROM[40672] <= 32'b00000000010100010010000000100011;
ROM[40673] <= 32'b00000000010000010000000100010011;
ROM[40674] <= 32'b00000000011000010010000000100011;
ROM[40675] <= 32'b00000000010000010000000100010011;
ROM[40676] <= 32'b00000001010000000000001110010011;
ROM[40677] <= 32'b00000000100000111000001110010011;
ROM[40678] <= 32'b01000000011100010000001110110011;
ROM[40679] <= 32'b00000000011100000000001000110011;
ROM[40680] <= 32'b00000000001000000000000110110011;
ROM[40681] <= 32'b00000000100000000010000011101111;
ROM[40682] <= 32'b00000110010100000000001110010011;
ROM[40683] <= 32'b00000000011100010010000000100011;
ROM[40684] <= 32'b00000000010000010000000100010011;
ROM[40685] <= 32'b00000000000000101000001110110111;
ROM[40686] <= 32'b11000000000000111000001110010011;
ROM[40687] <= 32'b00000000111000111000001110110011;
ROM[40688] <= 32'b00000000011100010010000000100011;
ROM[40689] <= 32'b00000000010000010000000100010011;
ROM[40690] <= 32'b00000000001100010010000000100011;
ROM[40691] <= 32'b00000000010000010000000100010011;
ROM[40692] <= 32'b00000000010000010010000000100011;
ROM[40693] <= 32'b00000000010000010000000100010011;
ROM[40694] <= 32'b00000000010100010010000000100011;
ROM[40695] <= 32'b00000000010000010000000100010011;
ROM[40696] <= 32'b00000000011000010010000000100011;
ROM[40697] <= 32'b00000000010000010000000100010011;
ROM[40698] <= 32'b00000001010000000000001110010011;
ROM[40699] <= 32'b00000000100000111000001110010011;
ROM[40700] <= 32'b01000000011100010000001110110011;
ROM[40701] <= 32'b00000000011100000000001000110011;
ROM[40702] <= 32'b00000000001000000000000110110011;
ROM[40703] <= 32'b01111011000100000001000011101111;
ROM[40704] <= 32'b00000110111000000000001110010011;
ROM[40705] <= 32'b00000000011100010010000000100011;
ROM[40706] <= 32'b00000000010000010000000100010011;
ROM[40707] <= 32'b00000000000000101000001110110111;
ROM[40708] <= 32'b11000101100000111000001110010011;
ROM[40709] <= 32'b00000000111000111000001110110011;
ROM[40710] <= 32'b00000000011100010010000000100011;
ROM[40711] <= 32'b00000000010000010000000100010011;
ROM[40712] <= 32'b00000000001100010010000000100011;
ROM[40713] <= 32'b00000000010000010000000100010011;
ROM[40714] <= 32'b00000000010000010010000000100011;
ROM[40715] <= 32'b00000000010000010000000100010011;
ROM[40716] <= 32'b00000000010100010010000000100011;
ROM[40717] <= 32'b00000000010000010000000100010011;
ROM[40718] <= 32'b00000000011000010010000000100011;
ROM[40719] <= 32'b00000000010000010000000100010011;
ROM[40720] <= 32'b00000001010000000000001110010011;
ROM[40721] <= 32'b00000000100000111000001110010011;
ROM[40722] <= 32'b01000000011100010000001110110011;
ROM[40723] <= 32'b00000000011100000000001000110011;
ROM[40724] <= 32'b00000000001000000000000110110011;
ROM[40725] <= 32'b01110101100100000001000011101111;
ROM[40726] <= 32'b00000110011100000000001110010011;
ROM[40727] <= 32'b00000000011100010010000000100011;
ROM[40728] <= 32'b00000000010000010000000100010011;
ROM[40729] <= 32'b00000000000000101000001110110111;
ROM[40730] <= 32'b11001011000000111000001110010011;
ROM[40731] <= 32'b00000000111000111000001110110011;
ROM[40732] <= 32'b00000000011100010010000000100011;
ROM[40733] <= 32'b00000000010000010000000100010011;
ROM[40734] <= 32'b00000000001100010010000000100011;
ROM[40735] <= 32'b00000000010000010000000100010011;
ROM[40736] <= 32'b00000000010000010010000000100011;
ROM[40737] <= 32'b00000000010000010000000100010011;
ROM[40738] <= 32'b00000000010100010010000000100011;
ROM[40739] <= 32'b00000000010000010000000100010011;
ROM[40740] <= 32'b00000000011000010010000000100011;
ROM[40741] <= 32'b00000000010000010000000100010011;
ROM[40742] <= 32'b00000001010000000000001110010011;
ROM[40743] <= 32'b00000000100000111000001110010011;
ROM[40744] <= 32'b01000000011100010000001110110011;
ROM[40745] <= 32'b00000000011100000000001000110011;
ROM[40746] <= 32'b00000000001000000000000110110011;
ROM[40747] <= 32'b01110000000100000001000011101111;
ROM[40748] <= 32'b00000111010000000000001110010011;
ROM[40749] <= 32'b00000000011100010010000000100011;
ROM[40750] <= 32'b00000000010000010000000100010011;
ROM[40751] <= 32'b00000000000000101000001110110111;
ROM[40752] <= 32'b11010000100000111000001110010011;
ROM[40753] <= 32'b00000000111000111000001110110011;
ROM[40754] <= 32'b00000000011100010010000000100011;
ROM[40755] <= 32'b00000000010000010000000100010011;
ROM[40756] <= 32'b00000000001100010010000000100011;
ROM[40757] <= 32'b00000000010000010000000100010011;
ROM[40758] <= 32'b00000000010000010010000000100011;
ROM[40759] <= 32'b00000000010000010000000100010011;
ROM[40760] <= 32'b00000000010100010010000000100011;
ROM[40761] <= 32'b00000000010000010000000100010011;
ROM[40762] <= 32'b00000000011000010010000000100011;
ROM[40763] <= 32'b00000000010000010000000100010011;
ROM[40764] <= 32'b00000001010000000000001110010011;
ROM[40765] <= 32'b00000000100000111000001110010011;
ROM[40766] <= 32'b01000000011100010000001110110011;
ROM[40767] <= 32'b00000000011100000000001000110011;
ROM[40768] <= 32'b00000000001000000000000110110011;
ROM[40769] <= 32'b01101010100100000001000011101111;
ROM[40770] <= 32'b00000110100000000000001110010011;
ROM[40771] <= 32'b00000000011100010010000000100011;
ROM[40772] <= 32'b00000000010000010000000100010011;
ROM[40773] <= 32'b00000000000000101000001110110111;
ROM[40774] <= 32'b11010110000000111000001110010011;
ROM[40775] <= 32'b00000000111000111000001110110011;
ROM[40776] <= 32'b00000000011100010010000000100011;
ROM[40777] <= 32'b00000000010000010000000100010011;
ROM[40778] <= 32'b00000000001100010010000000100011;
ROM[40779] <= 32'b00000000010000010000000100010011;
ROM[40780] <= 32'b00000000010000010010000000100011;
ROM[40781] <= 32'b00000000010000010000000100010011;
ROM[40782] <= 32'b00000000010100010010000000100011;
ROM[40783] <= 32'b00000000010000010000000100010011;
ROM[40784] <= 32'b00000000011000010010000000100011;
ROM[40785] <= 32'b00000000010000010000000100010011;
ROM[40786] <= 32'b00000001010000000000001110010011;
ROM[40787] <= 32'b00000000100000111000001110010011;
ROM[40788] <= 32'b01000000011100010000001110110011;
ROM[40789] <= 32'b00000000011100000000001000110011;
ROM[40790] <= 32'b00000000001000000000000110110011;
ROM[40791] <= 32'b01100101000100000001000011101111;
ROM[40792] <= 32'b00000011101000000000001110010011;
ROM[40793] <= 32'b00000000011100010010000000100011;
ROM[40794] <= 32'b00000000010000010000000100010011;
ROM[40795] <= 32'b00000000000000101000001110110111;
ROM[40796] <= 32'b11011011100000111000001110010011;
ROM[40797] <= 32'b00000000111000111000001110110011;
ROM[40798] <= 32'b00000000011100010010000000100011;
ROM[40799] <= 32'b00000000010000010000000100010011;
ROM[40800] <= 32'b00000000001100010010000000100011;
ROM[40801] <= 32'b00000000010000010000000100010011;
ROM[40802] <= 32'b00000000010000010010000000100011;
ROM[40803] <= 32'b00000000010000010000000100010011;
ROM[40804] <= 32'b00000000010100010010000000100011;
ROM[40805] <= 32'b00000000010000010000000100010011;
ROM[40806] <= 32'b00000000011000010010000000100011;
ROM[40807] <= 32'b00000000010000010000000100010011;
ROM[40808] <= 32'b00000001010000000000001110010011;
ROM[40809] <= 32'b00000000100000111000001110010011;
ROM[40810] <= 32'b01000000011100010000001110110011;
ROM[40811] <= 32'b00000000011100000000001000110011;
ROM[40812] <= 32'b00000000001000000000000110110011;
ROM[40813] <= 32'b01011111100100000001000011101111;
ROM[40814] <= 32'b00000010000000000000001110010011;
ROM[40815] <= 32'b00000000011100010010000000100011;
ROM[40816] <= 32'b00000000010000010000000100010011;
ROM[40817] <= 32'b00000000000000101000001110110111;
ROM[40818] <= 32'b11100001000000111000001110010011;
ROM[40819] <= 32'b00000000111000111000001110110011;
ROM[40820] <= 32'b00000000011100010010000000100011;
ROM[40821] <= 32'b00000000010000010000000100010011;
ROM[40822] <= 32'b00000000001100010010000000100011;
ROM[40823] <= 32'b00000000010000010000000100010011;
ROM[40824] <= 32'b00000000010000010010000000100011;
ROM[40825] <= 32'b00000000010000010000000100010011;
ROM[40826] <= 32'b00000000010100010010000000100011;
ROM[40827] <= 32'b00000000010000010000000100010011;
ROM[40828] <= 32'b00000000011000010010000000100011;
ROM[40829] <= 32'b00000000010000010000000100010011;
ROM[40830] <= 32'b00000001010000000000001110010011;
ROM[40831] <= 32'b00000000100000111000001110010011;
ROM[40832] <= 32'b01000000011100010000001110110011;
ROM[40833] <= 32'b00000000011100000000001000110011;
ROM[40834] <= 32'b00000000001000000000000110110011;
ROM[40835] <= 32'b01011010000100000001000011101111;
ROM[40836] <= 32'b11111111110000010000000100010011;
ROM[40837] <= 32'b00000000000000010010001110000011;
ROM[40838] <= 32'b00000000011100011010001000100011;
ROM[40839] <= 32'b00000000010000011010001110000011;
ROM[40840] <= 32'b00000000011100010010000000100011;
ROM[40841] <= 32'b00000000010000010000000100010011;
ROM[40842] <= 32'b00000000000000101000001110110111;
ROM[40843] <= 32'b11100111010000111000001110010011;
ROM[40844] <= 32'b00000000111000111000001110110011;
ROM[40845] <= 32'b00000000011100010010000000100011;
ROM[40846] <= 32'b00000000010000010000000100010011;
ROM[40847] <= 32'b00000000001100010010000000100011;
ROM[40848] <= 32'b00000000010000010000000100010011;
ROM[40849] <= 32'b00000000010000010010000000100011;
ROM[40850] <= 32'b00000000010000010000000100010011;
ROM[40851] <= 32'b00000000010100010010000000100011;
ROM[40852] <= 32'b00000000010000010000000100010011;
ROM[40853] <= 32'b00000000011000010010000000100011;
ROM[40854] <= 32'b00000000010000010000000100010011;
ROM[40855] <= 32'b00000001010000000000001110010011;
ROM[40856] <= 32'b00000000010000111000001110010011;
ROM[40857] <= 32'b01000000011100010000001110110011;
ROM[40858] <= 32'b00000000011100000000001000110011;
ROM[40859] <= 32'b00000000001000000000000110110011;
ROM[40860] <= 32'b10001111100011101111000011101111;
ROM[40861] <= 32'b11111111110000010000000100010011;
ROM[40862] <= 32'b00000000000000010010001110000011;
ROM[40863] <= 32'b00000000011101100010000000100011;
ROM[40864] <= 32'b00000000010000011010001110000011;
ROM[40865] <= 32'b00000000011100010010000000100011;
ROM[40866] <= 32'b00000000010000010000000100010011;
ROM[40867] <= 32'b00000000000000101000001110110111;
ROM[40868] <= 32'b11101101100000111000001110010011;
ROM[40869] <= 32'b00000000111000111000001110110011;
ROM[40870] <= 32'b00000000011100010010000000100011;
ROM[40871] <= 32'b00000000010000010000000100010011;
ROM[40872] <= 32'b00000000001100010010000000100011;
ROM[40873] <= 32'b00000000010000010000000100010011;
ROM[40874] <= 32'b00000000010000010010000000100011;
ROM[40875] <= 32'b00000000010000010000000100010011;
ROM[40876] <= 32'b00000000010100010010000000100011;
ROM[40877] <= 32'b00000000010000010000000100010011;
ROM[40878] <= 32'b00000000011000010010000000100011;
ROM[40879] <= 32'b00000000010000010000000100010011;
ROM[40880] <= 32'b00000001010000000000001110010011;
ROM[40881] <= 32'b00000000010000111000001110010011;
ROM[40882] <= 32'b01000000011100010000001110110011;
ROM[40883] <= 32'b00000000011100000000001000110011;
ROM[40884] <= 32'b00000000001000000000000110110011;
ROM[40885] <= 32'b01100011110100000010000011101111;
ROM[40886] <= 32'b11111111110000010000000100010011;
ROM[40887] <= 32'b00000000000000010010001110000011;
ROM[40888] <= 32'b00000000011101100010000000100011;
ROM[40889] <= 32'b00000000110100101000010000110011;
ROM[40890] <= 32'b00000000000001000010001110000011;
ROM[40891] <= 32'b00000000011100010010000000100011;
ROM[40892] <= 32'b00000000010000010000000100010011;
ROM[40893] <= 32'b00000000000000101000001110110111;
ROM[40894] <= 32'b11110100000000111000001110010011;
ROM[40895] <= 32'b00000000111000111000001110110011;
ROM[40896] <= 32'b00000000011100010010000000100011;
ROM[40897] <= 32'b00000000010000010000000100010011;
ROM[40898] <= 32'b00000000001100010010000000100011;
ROM[40899] <= 32'b00000000010000010000000100010011;
ROM[40900] <= 32'b00000000010000010010000000100011;
ROM[40901] <= 32'b00000000010000010000000100010011;
ROM[40902] <= 32'b00000000010100010010000000100011;
ROM[40903] <= 32'b00000000010000010000000100010011;
ROM[40904] <= 32'b00000000011000010010000000100011;
ROM[40905] <= 32'b00000000010000010000000100010011;
ROM[40906] <= 32'b00000001010000000000001110010011;
ROM[40907] <= 32'b00000000010000111000001110010011;
ROM[40908] <= 32'b01000000011100010000001110110011;
ROM[40909] <= 32'b00000000011100000000001000110011;
ROM[40910] <= 32'b00000000001000000000000110110011;
ROM[40911] <= 32'b10111000100111111011000011101111;
ROM[40912] <= 32'b11111111110000010000000100010011;
ROM[40913] <= 32'b00000000000000010010001110000011;
ROM[40914] <= 32'b00000000011100011010000000100011;
ROM[40915] <= 32'b00000000000000011010001110000011;
ROM[40916] <= 32'b00000000011100010010000000100011;
ROM[40917] <= 32'b00000000010000010000000100010011;
ROM[40918] <= 32'b00000000000000101000001110110111;
ROM[40919] <= 32'b11111010010000111000001110010011;
ROM[40920] <= 32'b00000000111000111000001110110011;
ROM[40921] <= 32'b00000000011100010010000000100011;
ROM[40922] <= 32'b00000000010000010000000100010011;
ROM[40923] <= 32'b00000000001100010010000000100011;
ROM[40924] <= 32'b00000000010000010000000100010011;
ROM[40925] <= 32'b00000000010000010010000000100011;
ROM[40926] <= 32'b00000000010000010000000100010011;
ROM[40927] <= 32'b00000000010100010010000000100011;
ROM[40928] <= 32'b00000000010000010000000100010011;
ROM[40929] <= 32'b00000000011000010010000000100011;
ROM[40930] <= 32'b00000000010000010000000100010011;
ROM[40931] <= 32'b00000001010000000000001110010011;
ROM[40932] <= 32'b00000000010000111000001110010011;
ROM[40933] <= 32'b01000000011100010000001110110011;
ROM[40934] <= 32'b00000000011100000000001000110011;
ROM[40935] <= 32'b00000000001000000000000110110011;
ROM[40936] <= 32'b11110001110011111000000011101111;
ROM[40937] <= 32'b00000000000000101000001110110111;
ROM[40938] <= 32'b11111111000000111000001110010011;
ROM[40939] <= 32'b00000000111000111000001110110011;
ROM[40940] <= 32'b00000000011100010010000000100011;
ROM[40941] <= 32'b00000000010000010000000100010011;
ROM[40942] <= 32'b00000000001100010010000000100011;
ROM[40943] <= 32'b00000000010000010000000100010011;
ROM[40944] <= 32'b00000000010000010010000000100011;
ROM[40945] <= 32'b00000000010000010000000100010011;
ROM[40946] <= 32'b00000000010100010010000000100011;
ROM[40947] <= 32'b00000000010000010000000100010011;
ROM[40948] <= 32'b00000000011000010010000000100011;
ROM[40949] <= 32'b00000000010000010000000100010011;
ROM[40950] <= 32'b00000001010000000000001110010011;
ROM[40951] <= 32'b00000000010000111000001110010011;
ROM[40952] <= 32'b01000000011100010000001110110011;
ROM[40953] <= 32'b00000000011100000000001000110011;
ROM[40954] <= 32'b00000000001000000000000110110011;
ROM[40955] <= 32'b10011001010011101111000011101111;
ROM[40956] <= 32'b11111111110000010000000100010011;
ROM[40957] <= 32'b00000000000000010010001110000011;
ROM[40958] <= 32'b00000000011101100010000000100011;
ROM[40959] <= 32'b00000000110100101000010000110011;
ROM[40960] <= 32'b00000000000001000010001110000011;
ROM[40961] <= 32'b00000000011100010010000000100011;
ROM[40962] <= 32'b00000000010000010000000100010011;
ROM[40963] <= 32'b00000000000000101000001110110111;
ROM[40964] <= 32'b00000101100000111000001110010011;
ROM[40965] <= 32'b00000000111000111000001110110011;
ROM[40966] <= 32'b00000000011100010010000000100011;
ROM[40967] <= 32'b00000000010000010000000100010011;
ROM[40968] <= 32'b00000000001100010010000000100011;
ROM[40969] <= 32'b00000000010000010000000100010011;
ROM[40970] <= 32'b00000000010000010010000000100011;
ROM[40971] <= 32'b00000000010000010000000100010011;
ROM[40972] <= 32'b00000000010100010010000000100011;
ROM[40973] <= 32'b00000000010000010000000100010011;
ROM[40974] <= 32'b00000000011000010010000000100011;
ROM[40975] <= 32'b00000000010000010000000100010011;
ROM[40976] <= 32'b00000001010000000000001110010011;
ROM[40977] <= 32'b00000000010000111000001110010011;
ROM[40978] <= 32'b01000000011100010000001110110011;
ROM[40979] <= 32'b00000000011100000000001000110011;
ROM[40980] <= 32'b00000000001000000000000110110011;
ROM[40981] <= 32'b10111111000111111011000011101111;
ROM[40982] <= 32'b11111111110000010000000100010011;
ROM[40983] <= 32'b00000000000000010010001110000011;
ROM[40984] <= 32'b00000000000000111000101001100011;
ROM[40985] <= 32'b00000000000000101000001110110111;
ROM[40986] <= 32'b00001101100000111000001110010011;
ROM[40987] <= 32'b00000000111000111000001110110011;
ROM[40988] <= 32'b00000000000000111000000011100111;
ROM[40989] <= 32'b00000000010100010010000000100011;
ROM[40990] <= 32'b00000000010000010000000100010011;
ROM[40991] <= 32'b00000000000000101000001110110111;
ROM[40992] <= 32'b00001100100000111000001110010011;
ROM[40993] <= 32'b00000000111000111000001110110011;
ROM[40994] <= 32'b00000000011100010010000000100011;
ROM[40995] <= 32'b00000000010000010000000100010011;
ROM[40996] <= 32'b00000000001100010010000000100011;
ROM[40997] <= 32'b00000000010000010000000100010011;
ROM[40998] <= 32'b00000000010000010010000000100011;
ROM[40999] <= 32'b00000000010000010000000100010011;
ROM[41000] <= 32'b00000000010100010010000000100011;
ROM[41001] <= 32'b00000000010000010000000100010011;
ROM[41002] <= 32'b00000000011000010010000000100011;
ROM[41003] <= 32'b00000000010000010000000100010011;
ROM[41004] <= 32'b00000001010000000000001110010011;
ROM[41005] <= 32'b00000000010000111000001110010011;
ROM[41006] <= 32'b01000000011100010000001110110011;
ROM[41007] <= 32'b00000000011100000000001000110011;
ROM[41008] <= 32'b00000000001000000000000110110011;
ROM[41009] <= 32'b01101000000000000000000011101111;
ROM[41010] <= 32'b11111111110000010000000100010011;
ROM[41011] <= 32'b00000000000000010010001110000011;
ROM[41012] <= 32'b00000000011101100010000000100011;
ROM[41013] <= 32'b00000110010000000000000011101111;
ROM[41014] <= 32'b00000000010100010010000000100011;
ROM[41015] <= 32'b00000000010000010000000100010011;
ROM[41016] <= 32'b00000000000000101000001110110111;
ROM[41017] <= 32'b00010010110000111000001110010011;
ROM[41018] <= 32'b00000000111000111000001110110011;
ROM[41019] <= 32'b00000000011100010010000000100011;
ROM[41020] <= 32'b00000000010000010000000100010011;
ROM[41021] <= 32'b00000000001100010010000000100011;
ROM[41022] <= 32'b00000000010000010000000100010011;
ROM[41023] <= 32'b00000000010000010010000000100011;
ROM[41024] <= 32'b00000000010000010000000100010011;
ROM[41025] <= 32'b00000000010100010010000000100011;
ROM[41026] <= 32'b00000000010000010000000100010011;
ROM[41027] <= 32'b00000000011000010010000000100011;
ROM[41028] <= 32'b00000000010000010000000100010011;
ROM[41029] <= 32'b00000001010000000000001110010011;
ROM[41030] <= 32'b00000000010000111000001110010011;
ROM[41031] <= 32'b01000000011100010000001110110011;
ROM[41032] <= 32'b00000000011100000000001000110011;
ROM[41033] <= 32'b00000000001000000000000110110011;
ROM[41034] <= 32'b00000101010000000000000011101111;
ROM[41035] <= 32'b11111111110000010000000100010011;
ROM[41036] <= 32'b00000000000000010010001110000011;
ROM[41037] <= 32'b00000000011101100010000000100011;
ROM[41038] <= 32'b00000000000000000000001110010011;
ROM[41039] <= 32'b00000000011100010010000000100011;
ROM[41040] <= 32'b00000000010000010000000100010011;
ROM[41041] <= 32'b00000001010000000000001110010011;
ROM[41042] <= 32'b01000000011100011000001110110011;
ROM[41043] <= 32'b00000000000000111010000010000011;
ROM[41044] <= 32'b11111111110000010000000100010011;
ROM[41045] <= 32'b00000000000000010010001110000011;
ROM[41046] <= 32'b00000000011100100010000000100011;
ROM[41047] <= 32'b00000000010000100000000100010011;
ROM[41048] <= 32'b00000001010000000000001110010011;
ROM[41049] <= 32'b01000000011100011000001110110011;
ROM[41050] <= 32'b00000000010000111010000110000011;
ROM[41051] <= 32'b00000000100000111010001000000011;
ROM[41052] <= 32'b00000000110000111010001010000011;
ROM[41053] <= 32'b00000001000000111010001100000011;
ROM[41054] <= 32'b00000000000000001000000011100111;
ROM[41055] <= 32'b00000000000000010010000000100011;
ROM[41056] <= 32'b00000000010000010000000100010011;
ROM[41057] <= 32'b00000000000000100010001110000011;
ROM[41058] <= 32'b00000000011100010010000000100011;
ROM[41059] <= 32'b00000000010000010000000100010011;
ROM[41060] <= 32'b11111111110000010000000100010011;
ROM[41061] <= 32'b00000000000000010010001110000011;
ROM[41062] <= 32'b00000000000000111000001010010011;
ROM[41063] <= 32'b00000001011000000000001110010011;
ROM[41064] <= 32'b00000000011100010010000000100011;
ROM[41065] <= 32'b00000000010000010000000100010011;
ROM[41066] <= 32'b00000000110000000000001110010011;
ROM[41067] <= 32'b00000000011100010010000000100011;
ROM[41068] <= 32'b00000000010000010000000100010011;
ROM[41069] <= 32'b00000000000000101000001110110111;
ROM[41070] <= 32'b00100000000000111000001110010011;
ROM[41071] <= 32'b00000000111000111000001110110011;
ROM[41072] <= 32'b00000000011100010010000000100011;
ROM[41073] <= 32'b00000000010000010000000100010011;
ROM[41074] <= 32'b00000000001100010010000000100011;
ROM[41075] <= 32'b00000000010000010000000100010011;
ROM[41076] <= 32'b00000000010000010010000000100011;
ROM[41077] <= 32'b00000000010000010000000100010011;
ROM[41078] <= 32'b00000000010100010010000000100011;
ROM[41079] <= 32'b00000000010000010000000100010011;
ROM[41080] <= 32'b00000000011000010010000000100011;
ROM[41081] <= 32'b00000000010000010000000100010011;
ROM[41082] <= 32'b00000001010000000000001110010011;
ROM[41083] <= 32'b00000000100000111000001110010011;
ROM[41084] <= 32'b01000000011100010000001110110011;
ROM[41085] <= 32'b00000000011100000000001000110011;
ROM[41086] <= 32'b00000000001000000000000110110011;
ROM[41087] <= 32'b10100000010111101101000011101111;
ROM[41088] <= 32'b11111111110000010000000100010011;
ROM[41089] <= 32'b00000000000000010010001110000011;
ROM[41090] <= 32'b00000000011101100010000000100011;
ROM[41091] <= 32'b00000000101100000000001110010011;
ROM[41092] <= 32'b00000000011100010010000000100011;
ROM[41093] <= 32'b00000000010000010000000100010011;
ROM[41094] <= 32'b00000000000000101000001110110111;
ROM[41095] <= 32'b00100110010000111000001110010011;
ROM[41096] <= 32'b00000000111000111000001110110011;
ROM[41097] <= 32'b00000000011100010010000000100011;
ROM[41098] <= 32'b00000000010000010000000100010011;
ROM[41099] <= 32'b00000000001100010010000000100011;
ROM[41100] <= 32'b00000000010000010000000100010011;
ROM[41101] <= 32'b00000000010000010010000000100011;
ROM[41102] <= 32'b00000000010000010000000100010011;
ROM[41103] <= 32'b00000000010100010010000000100011;
ROM[41104] <= 32'b00000000010000010000000100010011;
ROM[41105] <= 32'b00000000011000010010000000100011;
ROM[41106] <= 32'b00000000010000010000000100010011;
ROM[41107] <= 32'b00000001010000000000001110010011;
ROM[41108] <= 32'b00000000010000111000001110010011;
ROM[41109] <= 32'b01000000011100010000001110110011;
ROM[41110] <= 32'b00000000011100000000001000110011;
ROM[41111] <= 32'b00000000001000000000000110110011;
ROM[41112] <= 32'b01001101110000000001000011101111;
ROM[41113] <= 32'b00000101101100000000001110010011;
ROM[41114] <= 32'b00000000011100010010000000100011;
ROM[41115] <= 32'b00000000010000010000000100010011;
ROM[41116] <= 32'b00000000000000101000001110110111;
ROM[41117] <= 32'b00101011110000111000001110010011;
ROM[41118] <= 32'b00000000111000111000001110110011;
ROM[41119] <= 32'b00000000011100010010000000100011;
ROM[41120] <= 32'b00000000010000010000000100010011;
ROM[41121] <= 32'b00000000001100010010000000100011;
ROM[41122] <= 32'b00000000010000010000000100010011;
ROM[41123] <= 32'b00000000010000010010000000100011;
ROM[41124] <= 32'b00000000010000010000000100010011;
ROM[41125] <= 32'b00000000010100010010000000100011;
ROM[41126] <= 32'b00000000010000010000000100010011;
ROM[41127] <= 32'b00000000011000010010000000100011;
ROM[41128] <= 32'b00000000010000010000000100010011;
ROM[41129] <= 32'b00000001010000000000001110010011;
ROM[41130] <= 32'b00000000100000111000001110010011;
ROM[41131] <= 32'b01000000011100010000001110110011;
ROM[41132] <= 32'b00000000011100000000001000110011;
ROM[41133] <= 32'b00000000001000000000000110110011;
ROM[41134] <= 32'b00001111010100000001000011101111;
ROM[41135] <= 32'b00000101000000000000001110010011;
ROM[41136] <= 32'b00000000011100010010000000100011;
ROM[41137] <= 32'b00000000010000010000000100010011;
ROM[41138] <= 32'b00000000000000101000001110110111;
ROM[41139] <= 32'b00110001010000111000001110010011;
ROM[41140] <= 32'b00000000111000111000001110110011;
ROM[41141] <= 32'b00000000011100010010000000100011;
ROM[41142] <= 32'b00000000010000010000000100010011;
ROM[41143] <= 32'b00000000001100010010000000100011;
ROM[41144] <= 32'b00000000010000010000000100010011;
ROM[41145] <= 32'b00000000010000010010000000100011;
ROM[41146] <= 32'b00000000010000010000000100010011;
ROM[41147] <= 32'b00000000010100010010000000100011;
ROM[41148] <= 32'b00000000010000010000000100010011;
ROM[41149] <= 32'b00000000011000010010000000100011;
ROM[41150] <= 32'b00000000010000010000000100010011;
ROM[41151] <= 32'b00000001010000000000001110010011;
ROM[41152] <= 32'b00000000100000111000001110010011;
ROM[41153] <= 32'b01000000011100010000001110110011;
ROM[41154] <= 32'b00000000011100000000001000110011;
ROM[41155] <= 32'b00000000001000000000000110110011;
ROM[41156] <= 32'b00001001110100000001000011101111;
ROM[41157] <= 32'b00000100000100000000001110010011;
ROM[41158] <= 32'b00000000011100010010000000100011;
ROM[41159] <= 32'b00000000010000010000000100010011;
ROM[41160] <= 32'b00000000000000101000001110110111;
ROM[41161] <= 32'b00110110110000111000001110010011;
ROM[41162] <= 32'b00000000111000111000001110110011;
ROM[41163] <= 32'b00000000011100010010000000100011;
ROM[41164] <= 32'b00000000010000010000000100010011;
ROM[41165] <= 32'b00000000001100010010000000100011;
ROM[41166] <= 32'b00000000010000010000000100010011;
ROM[41167] <= 32'b00000000010000010010000000100011;
ROM[41168] <= 32'b00000000010000010000000100010011;
ROM[41169] <= 32'b00000000010100010010000000100011;
ROM[41170] <= 32'b00000000010000010000000100010011;
ROM[41171] <= 32'b00000000011000010010000000100011;
ROM[41172] <= 32'b00000000010000010000000100010011;
ROM[41173] <= 32'b00000001010000000000001110010011;
ROM[41174] <= 32'b00000000100000111000001110010011;
ROM[41175] <= 32'b01000000011100010000001110110011;
ROM[41176] <= 32'b00000000011100000000001000110011;
ROM[41177] <= 32'b00000000001000000000000110110011;
ROM[41178] <= 32'b00000100010100000001000011101111;
ROM[41179] <= 32'b00000101010100000000001110010011;
ROM[41180] <= 32'b00000000011100010010000000100011;
ROM[41181] <= 32'b00000000010000010000000100010011;
ROM[41182] <= 32'b00000000000000101000001110110111;
ROM[41183] <= 32'b00111100010000111000001110010011;
ROM[41184] <= 32'b00000000111000111000001110110011;
ROM[41185] <= 32'b00000000011100010010000000100011;
ROM[41186] <= 32'b00000000010000010000000100010011;
ROM[41187] <= 32'b00000000001100010010000000100011;
ROM[41188] <= 32'b00000000010000010000000100010011;
ROM[41189] <= 32'b00000000010000010010000000100011;
ROM[41190] <= 32'b00000000010000010000000100010011;
ROM[41191] <= 32'b00000000010100010010000000100011;
ROM[41192] <= 32'b00000000010000010000000100010011;
ROM[41193] <= 32'b00000000011000010010000000100011;
ROM[41194] <= 32'b00000000010000010000000100010011;
ROM[41195] <= 32'b00000001010000000000001110010011;
ROM[41196] <= 32'b00000000100000111000001110010011;
ROM[41197] <= 32'b01000000011100010000001110110011;
ROM[41198] <= 32'b00000000011100000000001000110011;
ROM[41199] <= 32'b00000000001000000000000110110011;
ROM[41200] <= 32'b01111110110000000001000011101111;
ROM[41201] <= 32'b00000101001100000000001110010011;
ROM[41202] <= 32'b00000000011100010010000000100011;
ROM[41203] <= 32'b00000000010000010000000100010011;
ROM[41204] <= 32'b00000000000000101000001110110111;
ROM[41205] <= 32'b01000001110000111000001110010011;
ROM[41206] <= 32'b00000000111000111000001110110011;
ROM[41207] <= 32'b00000000011100010010000000100011;
ROM[41208] <= 32'b00000000010000010000000100010011;
ROM[41209] <= 32'b00000000001100010010000000100011;
ROM[41210] <= 32'b00000000010000010000000100010011;
ROM[41211] <= 32'b00000000010000010010000000100011;
ROM[41212] <= 32'b00000000010000010000000100010011;
ROM[41213] <= 32'b00000000010100010010000000100011;
ROM[41214] <= 32'b00000000010000010000000100010011;
ROM[41215] <= 32'b00000000011000010010000000100011;
ROM[41216] <= 32'b00000000010000010000000100010011;
ROM[41217] <= 32'b00000001010000000000001110010011;
ROM[41218] <= 32'b00000000100000111000001110010011;
ROM[41219] <= 32'b01000000011100010000001110110011;
ROM[41220] <= 32'b00000000011100000000001000110011;
ROM[41221] <= 32'b00000000001000000000000110110011;
ROM[41222] <= 32'b01111001010000000001000011101111;
ROM[41223] <= 32'b00000100010100000000001110010011;
ROM[41224] <= 32'b00000000011100010010000000100011;
ROM[41225] <= 32'b00000000010000010000000100010011;
ROM[41226] <= 32'b00000000000000101000001110110111;
ROM[41227] <= 32'b01000111010000111000001110010011;
ROM[41228] <= 32'b00000000111000111000001110110011;
ROM[41229] <= 32'b00000000011100010010000000100011;
ROM[41230] <= 32'b00000000010000010000000100010011;
ROM[41231] <= 32'b00000000001100010010000000100011;
ROM[41232] <= 32'b00000000010000010000000100010011;
ROM[41233] <= 32'b00000000010000010010000000100011;
ROM[41234] <= 32'b00000000010000010000000100010011;
ROM[41235] <= 32'b00000000010100010010000000100011;
ROM[41236] <= 32'b00000000010000010000000100010011;
ROM[41237] <= 32'b00000000011000010010000000100011;
ROM[41238] <= 32'b00000000010000010000000100010011;
ROM[41239] <= 32'b00000001010000000000001110010011;
ROM[41240] <= 32'b00000000100000111000001110010011;
ROM[41241] <= 32'b01000000011100010000001110110011;
ROM[41242] <= 32'b00000000011100000000001000110011;
ROM[41243] <= 32'b00000000001000000000000110110011;
ROM[41244] <= 32'b01110011110000000001000011101111;
ROM[41245] <= 32'b00000100010000000000001110010011;
ROM[41246] <= 32'b00000000011100010010000000100011;
ROM[41247] <= 32'b00000000010000010000000100010011;
ROM[41248] <= 32'b00000000000000101000001110110111;
ROM[41249] <= 32'b01001100110000111000001110010011;
ROM[41250] <= 32'b00000000111000111000001110110011;
ROM[41251] <= 32'b00000000011100010010000000100011;
ROM[41252] <= 32'b00000000010000010000000100010011;
ROM[41253] <= 32'b00000000001100010010000000100011;
ROM[41254] <= 32'b00000000010000010000000100010011;
ROM[41255] <= 32'b00000000010000010010000000100011;
ROM[41256] <= 32'b00000000010000010000000100010011;
ROM[41257] <= 32'b00000000010100010010000000100011;
ROM[41258] <= 32'b00000000010000010000000100010011;
ROM[41259] <= 32'b00000000011000010010000000100011;
ROM[41260] <= 32'b00000000010000010000000100010011;
ROM[41261] <= 32'b00000001010000000000001110010011;
ROM[41262] <= 32'b00000000100000111000001110010011;
ROM[41263] <= 32'b01000000011100010000001110110011;
ROM[41264] <= 32'b00000000011100000000001000110011;
ROM[41265] <= 32'b00000000001000000000000110110011;
ROM[41266] <= 32'b01101110010000000001000011101111;
ROM[41267] <= 32'b00000010101000000000001110010011;
ROM[41268] <= 32'b00000000011100010010000000100011;
ROM[41269] <= 32'b00000000010000010000000100010011;
ROM[41270] <= 32'b00000000000000101000001110110111;
ROM[41271] <= 32'b01010010010000111000001110010011;
ROM[41272] <= 32'b00000000111000111000001110110011;
ROM[41273] <= 32'b00000000011100010010000000100011;
ROM[41274] <= 32'b00000000010000010000000100010011;
ROM[41275] <= 32'b00000000001100010010000000100011;
ROM[41276] <= 32'b00000000010000010000000100010011;
ROM[41277] <= 32'b00000000010000010010000000100011;
ROM[41278] <= 32'b00000000010000010000000100010011;
ROM[41279] <= 32'b00000000010100010010000000100011;
ROM[41280] <= 32'b00000000010000010000000100010011;
ROM[41281] <= 32'b00000000011000010010000000100011;
ROM[41282] <= 32'b00000000010000010000000100010011;
ROM[41283] <= 32'b00000001010000000000001110010011;
ROM[41284] <= 32'b00000000100000111000001110010011;
ROM[41285] <= 32'b01000000011100010000001110110011;
ROM[41286] <= 32'b00000000011100000000001000110011;
ROM[41287] <= 32'b00000000001000000000000110110011;
ROM[41288] <= 32'b01101000110000000001000011101111;
ROM[41289] <= 32'b00000011010000000000001110010011;
ROM[41290] <= 32'b00000000011100010010000000100011;
ROM[41291] <= 32'b00000000010000010000000100010011;
ROM[41292] <= 32'b00000000000000101000001110110111;
ROM[41293] <= 32'b01010111110000111000001110010011;
ROM[41294] <= 32'b00000000111000111000001110110011;
ROM[41295] <= 32'b00000000011100010010000000100011;
ROM[41296] <= 32'b00000000010000010000000100010011;
ROM[41297] <= 32'b00000000001100010010000000100011;
ROM[41298] <= 32'b00000000010000010000000100010011;
ROM[41299] <= 32'b00000000010000010010000000100011;
ROM[41300] <= 32'b00000000010000010000000100010011;
ROM[41301] <= 32'b00000000010100010010000000100011;
ROM[41302] <= 32'b00000000010000010000000100010011;
ROM[41303] <= 32'b00000000011000010010000000100011;
ROM[41304] <= 32'b00000000010000010000000100010011;
ROM[41305] <= 32'b00000001010000000000001110010011;
ROM[41306] <= 32'b00000000100000111000001110010011;
ROM[41307] <= 32'b01000000011100010000001110110011;
ROM[41308] <= 32'b00000000011100000000001000110011;
ROM[41309] <= 32'b00000000001000000000000110110011;
ROM[41310] <= 32'b01100011010000000001000011101111;
ROM[41311] <= 32'b00000101110100000000001110010011;
ROM[41312] <= 32'b00000000011100010010000000100011;
ROM[41313] <= 32'b00000000010000010000000100010011;
ROM[41314] <= 32'b00000000000000101000001110110111;
ROM[41315] <= 32'b01011101010000111000001110010011;
ROM[41316] <= 32'b00000000111000111000001110110011;
ROM[41317] <= 32'b00000000011100010010000000100011;
ROM[41318] <= 32'b00000000010000010000000100010011;
ROM[41319] <= 32'b00000000001100010010000000100011;
ROM[41320] <= 32'b00000000010000010000000100010011;
ROM[41321] <= 32'b00000000010000010010000000100011;
ROM[41322] <= 32'b00000000010000010000000100010011;
ROM[41323] <= 32'b00000000010100010010000000100011;
ROM[41324] <= 32'b00000000010000010000000100010011;
ROM[41325] <= 32'b00000000011000010010000000100011;
ROM[41326] <= 32'b00000000010000010000000100010011;
ROM[41327] <= 32'b00000001010000000000001110010011;
ROM[41328] <= 32'b00000000100000111000001110010011;
ROM[41329] <= 32'b01000000011100010000001110110011;
ROM[41330] <= 32'b00000000011100000000001000110011;
ROM[41331] <= 32'b00000000001000000000000110110011;
ROM[41332] <= 32'b01011101110000000001000011101111;
ROM[41333] <= 32'b00000010000000000000001110010011;
ROM[41334] <= 32'b00000000011100010010000000100011;
ROM[41335] <= 32'b00000000010000010000000100010011;
ROM[41336] <= 32'b00000000000000101000001110110111;
ROM[41337] <= 32'b01100010110000111000001110010011;
ROM[41338] <= 32'b00000000111000111000001110110011;
ROM[41339] <= 32'b00000000011100010010000000100011;
ROM[41340] <= 32'b00000000010000010000000100010011;
ROM[41341] <= 32'b00000000001100010010000000100011;
ROM[41342] <= 32'b00000000010000010000000100010011;
ROM[41343] <= 32'b00000000010000010010000000100011;
ROM[41344] <= 32'b00000000010000010000000100010011;
ROM[41345] <= 32'b00000000010100010010000000100011;
ROM[41346] <= 32'b00000000010000010000000100010011;
ROM[41347] <= 32'b00000000011000010010000000100011;
ROM[41348] <= 32'b00000000010000010000000100010011;
ROM[41349] <= 32'b00000001010000000000001110010011;
ROM[41350] <= 32'b00000000100000111000001110010011;
ROM[41351] <= 32'b01000000011100010000001110110011;
ROM[41352] <= 32'b00000000011100000000001000110011;
ROM[41353] <= 32'b00000000001000000000000110110011;
ROM[41354] <= 32'b01011000010000000001000011101111;
ROM[41355] <= 32'b11111111110000010000000100010011;
ROM[41356] <= 32'b00000000000000010010001110000011;
ROM[41357] <= 32'b00000000011100011010000000100011;
ROM[41358] <= 32'b00000000000000011010001110000011;
ROM[41359] <= 32'b00000000011100010010000000100011;
ROM[41360] <= 32'b00000000010000010000000100010011;
ROM[41361] <= 32'b00000000000000101000001110110111;
ROM[41362] <= 32'b01101001000000111000001110010011;
ROM[41363] <= 32'b00000000111000111000001110110011;
ROM[41364] <= 32'b00000000011100010010000000100011;
ROM[41365] <= 32'b00000000010000010000000100010011;
ROM[41366] <= 32'b00000000001100010010000000100011;
ROM[41367] <= 32'b00000000010000010000000100010011;
ROM[41368] <= 32'b00000000010000010010000000100011;
ROM[41369] <= 32'b00000000010000010000000100010011;
ROM[41370] <= 32'b00000000010100010010000000100011;
ROM[41371] <= 32'b00000000010000010000000100010011;
ROM[41372] <= 32'b00000000011000010010000000100011;
ROM[41373] <= 32'b00000000010000010000000100010011;
ROM[41374] <= 32'b00000001010000000000001110010011;
ROM[41375] <= 32'b00000000010000111000001110010011;
ROM[41376] <= 32'b01000000011100010000001110110011;
ROM[41377] <= 32'b00000000011100000000001000110011;
ROM[41378] <= 32'b00000000001000000000000110110011;
ROM[41379] <= 32'b10001101110111101110000011101111;
ROM[41380] <= 32'b11111111110000010000000100010011;
ROM[41381] <= 32'b00000000000000010010001110000011;
ROM[41382] <= 32'b00000000011101100010000000100011;
ROM[41383] <= 32'b00000000000000011010001110000011;
ROM[41384] <= 32'b00000000011100010010000000100011;
ROM[41385] <= 32'b00000000010000010000000100010011;
ROM[41386] <= 32'b00000000000000101000001110110111;
ROM[41387] <= 32'b01101111010000111000001110010011;
ROM[41388] <= 32'b00000000111000111000001110110011;
ROM[41389] <= 32'b00000000011100010010000000100011;
ROM[41390] <= 32'b00000000010000010000000100010011;
ROM[41391] <= 32'b00000000001100010010000000100011;
ROM[41392] <= 32'b00000000010000010000000100010011;
ROM[41393] <= 32'b00000000010000010010000000100011;
ROM[41394] <= 32'b00000000010000010000000100010011;
ROM[41395] <= 32'b00000000010100010010000000100011;
ROM[41396] <= 32'b00000000010000010000000100010011;
ROM[41397] <= 32'b00000000011000010010000000100011;
ROM[41398] <= 32'b00000000010000010000000100010011;
ROM[41399] <= 32'b00000001010000000000001110010011;
ROM[41400] <= 32'b00000000010000111000001110010011;
ROM[41401] <= 32'b01000000011100010000001110110011;
ROM[41402] <= 32'b00000000011100000000001000110011;
ROM[41403] <= 32'b00000000001000000000000110110011;
ROM[41404] <= 32'b01100010000000000010000011101111;
ROM[41405] <= 32'b11111111110000010000000100010011;
ROM[41406] <= 32'b00000000000000010010001110000011;
ROM[41407] <= 32'b00000000011101100010000000100011;
ROM[41408] <= 32'b00000000000000000000001110010011;
ROM[41409] <= 32'b00000000011100010010000000100011;
ROM[41410] <= 32'b00000000010000010000000100010011;
ROM[41411] <= 32'b00000001010000000000001110010011;
ROM[41412] <= 32'b01000000011100011000001110110011;
ROM[41413] <= 32'b00000000000000111010000010000011;
ROM[41414] <= 32'b11111111110000010000000100010011;
ROM[41415] <= 32'b00000000000000010010001110000011;
ROM[41416] <= 32'b00000000011100100010000000100011;
ROM[41417] <= 32'b00000000010000100000000100010011;
ROM[41418] <= 32'b00000001010000000000001110010011;
ROM[41419] <= 32'b01000000011100011000001110110011;
ROM[41420] <= 32'b00000000010000111010000110000011;
ROM[41421] <= 32'b00000000100000111010001000000011;
ROM[41422] <= 32'b00000000110000111010001010000011;
ROM[41423] <= 32'b00000001000000111010001100000011;
ROM[41424] <= 32'b00000000000000001000000011100111;
ROM[41425] <= 32'b00000000000000010010000000100011;
ROM[41426] <= 32'b00000000010000010000000100010011;
ROM[41427] <= 32'b00000000000000100010001110000011;
ROM[41428] <= 32'b00000000011100010010000000100011;
ROM[41429] <= 32'b00000000010000010000000100010011;
ROM[41430] <= 32'b11111111110000010000000100010011;
ROM[41431] <= 32'b00000000000000010010001110000011;
ROM[41432] <= 32'b00000000000000111000001010010011;
ROM[41433] <= 32'b00000001011000000000001110010011;
ROM[41434] <= 32'b00000000011100010010000000100011;
ROM[41435] <= 32'b00000000010000010000000100010011;
ROM[41436] <= 32'b00000000110000000000001110010011;
ROM[41437] <= 32'b00000000011100010010000000100011;
ROM[41438] <= 32'b00000000010000010000000100010011;
ROM[41439] <= 32'b00000000000000101000001110110111;
ROM[41440] <= 32'b01111100100000111000001110010011;
ROM[41441] <= 32'b00000000111000111000001110110011;
ROM[41442] <= 32'b00000000011100010010000000100011;
ROM[41443] <= 32'b00000000010000010000000100010011;
ROM[41444] <= 32'b00000000001100010010000000100011;
ROM[41445] <= 32'b00000000010000010000000100010011;
ROM[41446] <= 32'b00000000010000010010000000100011;
ROM[41447] <= 32'b00000000010000010000000100010011;
ROM[41448] <= 32'b00000000010100010010000000100011;
ROM[41449] <= 32'b00000000010000010000000100010011;
ROM[41450] <= 32'b00000000011000010010000000100011;
ROM[41451] <= 32'b00000000010000010000000100010011;
ROM[41452] <= 32'b00000001010000000000001110010011;
ROM[41453] <= 32'b00000000100000111000001110010011;
ROM[41454] <= 32'b01000000011100010000001110110011;
ROM[41455] <= 32'b00000000011100000000001000110011;
ROM[41456] <= 32'b00000000001000000000000110110011;
ROM[41457] <= 32'b11000011110011101101000011101111;
ROM[41458] <= 32'b11111111110000010000000100010011;
ROM[41459] <= 32'b00000000000000010010001110000011;
ROM[41460] <= 32'b00000000011101100010000000100011;
ROM[41461] <= 32'b00000000100100000000001110010011;
ROM[41462] <= 32'b00000000011100010010000000100011;
ROM[41463] <= 32'b00000000010000010000000100010011;
ROM[41464] <= 32'b00000000000000101001001110110111;
ROM[41465] <= 32'b10000010110000111000001110010011;
ROM[41466] <= 32'b00000000111000111000001110110011;
ROM[41467] <= 32'b00000000011100010010000000100011;
ROM[41468] <= 32'b00000000010000010000000100010011;
ROM[41469] <= 32'b00000000001100010010000000100011;
ROM[41470] <= 32'b00000000010000010000000100010011;
ROM[41471] <= 32'b00000000010000010010000000100011;
ROM[41472] <= 32'b00000000010000010000000100010011;
ROM[41473] <= 32'b00000000010100010010000000100011;
ROM[41474] <= 32'b00000000010000010000000100010011;
ROM[41475] <= 32'b00000000011000010010000000100011;
ROM[41476] <= 32'b00000000010000010000000100010011;
ROM[41477] <= 32'b00000001010000000000001110010011;
ROM[41478] <= 32'b00000000010000111000001110010011;
ROM[41479] <= 32'b01000000011100010000001110110011;
ROM[41480] <= 32'b00000000011100000000001000110011;
ROM[41481] <= 32'b00000000001000000000000110110011;
ROM[41482] <= 32'b01110001010100000000000011101111;
ROM[41483] <= 32'b00000010000000000000001110010011;
ROM[41484] <= 32'b00000000011100010010000000100011;
ROM[41485] <= 32'b00000000010000010000000100010011;
ROM[41486] <= 32'b00000000000000101001001110110111;
ROM[41487] <= 32'b10001000010000111000001110010011;
ROM[41488] <= 32'b00000000111000111000001110110011;
ROM[41489] <= 32'b00000000011100010010000000100011;
ROM[41490] <= 32'b00000000010000010000000100010011;
ROM[41491] <= 32'b00000000001100010010000000100011;
ROM[41492] <= 32'b00000000010000010000000100010011;
ROM[41493] <= 32'b00000000010000010010000000100011;
ROM[41494] <= 32'b00000000010000010000000100010011;
ROM[41495] <= 32'b00000000010100010010000000100011;
ROM[41496] <= 32'b00000000010000010000000100010011;
ROM[41497] <= 32'b00000000011000010010000000100011;
ROM[41498] <= 32'b00000000010000010000000100010011;
ROM[41499] <= 32'b00000001010000000000001110010011;
ROM[41500] <= 32'b00000000100000111000001110010011;
ROM[41501] <= 32'b01000000011100010000001110110011;
ROM[41502] <= 32'b00000000011100000000001000110011;
ROM[41503] <= 32'b00000000001000000000000110110011;
ROM[41504] <= 32'b00110010110000000001000011101111;
ROM[41505] <= 32'b00000010000000000000001110010011;
ROM[41506] <= 32'b00000000011100010010000000100011;
ROM[41507] <= 32'b00000000010000010000000100010011;
ROM[41508] <= 32'b00000000000000101001001110110111;
ROM[41509] <= 32'b10001101110000111000001110010011;
ROM[41510] <= 32'b00000000111000111000001110110011;
ROM[41511] <= 32'b00000000011100010010000000100011;
ROM[41512] <= 32'b00000000010000010000000100010011;
ROM[41513] <= 32'b00000000001100010010000000100011;
ROM[41514] <= 32'b00000000010000010000000100010011;
ROM[41515] <= 32'b00000000010000010010000000100011;
ROM[41516] <= 32'b00000000010000010000000100010011;
ROM[41517] <= 32'b00000000010100010010000000100011;
ROM[41518] <= 32'b00000000010000010000000100010011;
ROM[41519] <= 32'b00000000011000010010000000100011;
ROM[41520] <= 32'b00000000010000010000000100010011;
ROM[41521] <= 32'b00000001010000000000001110010011;
ROM[41522] <= 32'b00000000100000111000001110010011;
ROM[41523] <= 32'b01000000011100010000001110110011;
ROM[41524] <= 32'b00000000011100000000001000110011;
ROM[41525] <= 32'b00000000001000000000000110110011;
ROM[41526] <= 32'b00101101010000000001000011101111;
ROM[41527] <= 32'b00000010000000000000001110010011;
ROM[41528] <= 32'b00000000011100010010000000100011;
ROM[41529] <= 32'b00000000010000010000000100010011;
ROM[41530] <= 32'b00000000000000101001001110110111;
ROM[41531] <= 32'b10010011010000111000001110010011;
ROM[41532] <= 32'b00000000111000111000001110110011;
ROM[41533] <= 32'b00000000011100010010000000100011;
ROM[41534] <= 32'b00000000010000010000000100010011;
ROM[41535] <= 32'b00000000001100010010000000100011;
ROM[41536] <= 32'b00000000010000010000000100010011;
ROM[41537] <= 32'b00000000010000010010000000100011;
ROM[41538] <= 32'b00000000010000010000000100010011;
ROM[41539] <= 32'b00000000010100010010000000100011;
ROM[41540] <= 32'b00000000010000010000000100010011;
ROM[41541] <= 32'b00000000011000010010000000100011;
ROM[41542] <= 32'b00000000010000010000000100010011;
ROM[41543] <= 32'b00000001010000000000001110010011;
ROM[41544] <= 32'b00000000100000111000001110010011;
ROM[41545] <= 32'b01000000011100010000001110110011;
ROM[41546] <= 32'b00000000011100000000001000110011;
ROM[41547] <= 32'b00000000001000000000000110110011;
ROM[41548] <= 32'b00100111110000000001000011101111;
ROM[41549] <= 32'b00000010000000000000001110010011;
ROM[41550] <= 32'b00000000011100010010000000100011;
ROM[41551] <= 32'b00000000010000010000000100010011;
ROM[41552] <= 32'b00000000000000101001001110110111;
ROM[41553] <= 32'b10011000110000111000001110010011;
ROM[41554] <= 32'b00000000111000111000001110110011;
ROM[41555] <= 32'b00000000011100010010000000100011;
ROM[41556] <= 32'b00000000010000010000000100010011;
ROM[41557] <= 32'b00000000001100010010000000100011;
ROM[41558] <= 32'b00000000010000010000000100010011;
ROM[41559] <= 32'b00000000010000010010000000100011;
ROM[41560] <= 32'b00000000010000010000000100010011;
ROM[41561] <= 32'b00000000010100010010000000100011;
ROM[41562] <= 32'b00000000010000010000000100010011;
ROM[41563] <= 32'b00000000011000010010000000100011;
ROM[41564] <= 32'b00000000010000010000000100010011;
ROM[41565] <= 32'b00000001010000000000001110010011;
ROM[41566] <= 32'b00000000100000111000001110010011;
ROM[41567] <= 32'b01000000011100010000001110110011;
ROM[41568] <= 32'b00000000011100000000001000110011;
ROM[41569] <= 32'b00000000001000000000000110110011;
ROM[41570] <= 32'b00100010010000000001000011101111;
ROM[41571] <= 32'b00000010000000000000001110010011;
ROM[41572] <= 32'b00000000011100010010000000100011;
ROM[41573] <= 32'b00000000010000010000000100010011;
ROM[41574] <= 32'b00000000000000101001001110110111;
ROM[41575] <= 32'b10011110010000111000001110010011;
ROM[41576] <= 32'b00000000111000111000001110110011;
ROM[41577] <= 32'b00000000011100010010000000100011;
ROM[41578] <= 32'b00000000010000010000000100010011;
ROM[41579] <= 32'b00000000001100010010000000100011;
ROM[41580] <= 32'b00000000010000010000000100010011;
ROM[41581] <= 32'b00000000010000010010000000100011;
ROM[41582] <= 32'b00000000010000010000000100010011;
ROM[41583] <= 32'b00000000010100010010000000100011;
ROM[41584] <= 32'b00000000010000010000000100010011;
ROM[41585] <= 32'b00000000011000010010000000100011;
ROM[41586] <= 32'b00000000010000010000000100010011;
ROM[41587] <= 32'b00000001010000000000001110010011;
ROM[41588] <= 32'b00000000100000111000001110010011;
ROM[41589] <= 32'b01000000011100010000001110110011;
ROM[41590] <= 32'b00000000011100000000001000110011;
ROM[41591] <= 32'b00000000001000000000000110110011;
ROM[41592] <= 32'b00011100110000000001000011101111;
ROM[41593] <= 32'b00000010000000000000001110010011;
ROM[41594] <= 32'b00000000011100010010000000100011;
ROM[41595] <= 32'b00000000010000010000000100010011;
ROM[41596] <= 32'b00000000000000101001001110110111;
ROM[41597] <= 32'b10100011110000111000001110010011;
ROM[41598] <= 32'b00000000111000111000001110110011;
ROM[41599] <= 32'b00000000011100010010000000100011;
ROM[41600] <= 32'b00000000010000010000000100010011;
ROM[41601] <= 32'b00000000001100010010000000100011;
ROM[41602] <= 32'b00000000010000010000000100010011;
ROM[41603] <= 32'b00000000010000010010000000100011;
ROM[41604] <= 32'b00000000010000010000000100010011;
ROM[41605] <= 32'b00000000010100010010000000100011;
ROM[41606] <= 32'b00000000010000010000000100010011;
ROM[41607] <= 32'b00000000011000010010000000100011;
ROM[41608] <= 32'b00000000010000010000000100010011;
ROM[41609] <= 32'b00000001010000000000001110010011;
ROM[41610] <= 32'b00000000100000111000001110010011;
ROM[41611] <= 32'b01000000011100010000001110110011;
ROM[41612] <= 32'b00000000011100000000001000110011;
ROM[41613] <= 32'b00000000001000000000000110110011;
ROM[41614] <= 32'b00010111010000000001000011101111;
ROM[41615] <= 32'b00000010000000000000001110010011;
ROM[41616] <= 32'b00000000011100010010000000100011;
ROM[41617] <= 32'b00000000010000010000000100010011;
ROM[41618] <= 32'b00000000000000101001001110110111;
ROM[41619] <= 32'b10101001010000111000001110010011;
ROM[41620] <= 32'b00000000111000111000001110110011;
ROM[41621] <= 32'b00000000011100010010000000100011;
ROM[41622] <= 32'b00000000010000010000000100010011;
ROM[41623] <= 32'b00000000001100010010000000100011;
ROM[41624] <= 32'b00000000010000010000000100010011;
ROM[41625] <= 32'b00000000010000010010000000100011;
ROM[41626] <= 32'b00000000010000010000000100010011;
ROM[41627] <= 32'b00000000010100010010000000100011;
ROM[41628] <= 32'b00000000010000010000000100010011;
ROM[41629] <= 32'b00000000011000010010000000100011;
ROM[41630] <= 32'b00000000010000010000000100010011;
ROM[41631] <= 32'b00000001010000000000001110010011;
ROM[41632] <= 32'b00000000100000111000001110010011;
ROM[41633] <= 32'b01000000011100010000001110110011;
ROM[41634] <= 32'b00000000011100000000001000110011;
ROM[41635] <= 32'b00000000001000000000000110110011;
ROM[41636] <= 32'b00010001110000000001000011101111;
ROM[41637] <= 32'b00000010000000000000001110010011;
ROM[41638] <= 32'b00000000011100010010000000100011;
ROM[41639] <= 32'b00000000010000010000000100010011;
ROM[41640] <= 32'b00000000000000101001001110110111;
ROM[41641] <= 32'b10101110110000111000001110010011;
ROM[41642] <= 32'b00000000111000111000001110110011;
ROM[41643] <= 32'b00000000011100010010000000100011;
ROM[41644] <= 32'b00000000010000010000000100010011;
ROM[41645] <= 32'b00000000001100010010000000100011;
ROM[41646] <= 32'b00000000010000010000000100010011;
ROM[41647] <= 32'b00000000010000010010000000100011;
ROM[41648] <= 32'b00000000010000010000000100010011;
ROM[41649] <= 32'b00000000010100010010000000100011;
ROM[41650] <= 32'b00000000010000010000000100010011;
ROM[41651] <= 32'b00000000011000010010000000100011;
ROM[41652] <= 32'b00000000010000010000000100010011;
ROM[41653] <= 32'b00000001010000000000001110010011;
ROM[41654] <= 32'b00000000100000111000001110010011;
ROM[41655] <= 32'b01000000011100010000001110110011;
ROM[41656] <= 32'b00000000011100000000001000110011;
ROM[41657] <= 32'b00000000001000000000000110110011;
ROM[41658] <= 32'b00001100010000000001000011101111;
ROM[41659] <= 32'b00000010000000000000001110010011;
ROM[41660] <= 32'b00000000011100010010000000100011;
ROM[41661] <= 32'b00000000010000010000000100010011;
ROM[41662] <= 32'b00000000000000101001001110110111;
ROM[41663] <= 32'b10110100010000111000001110010011;
ROM[41664] <= 32'b00000000111000111000001110110011;
ROM[41665] <= 32'b00000000011100010010000000100011;
ROM[41666] <= 32'b00000000010000010000000100010011;
ROM[41667] <= 32'b00000000001100010010000000100011;
ROM[41668] <= 32'b00000000010000010000000100010011;
ROM[41669] <= 32'b00000000010000010010000000100011;
ROM[41670] <= 32'b00000000010000010000000100010011;
ROM[41671] <= 32'b00000000010100010010000000100011;
ROM[41672] <= 32'b00000000010000010000000100010011;
ROM[41673] <= 32'b00000000011000010010000000100011;
ROM[41674] <= 32'b00000000010000010000000100010011;
ROM[41675] <= 32'b00000001010000000000001110010011;
ROM[41676] <= 32'b00000000100000111000001110010011;
ROM[41677] <= 32'b01000000011100010000001110110011;
ROM[41678] <= 32'b00000000011100000000001000110011;
ROM[41679] <= 32'b00000000001000000000000110110011;
ROM[41680] <= 32'b00000110110000000001000011101111;
ROM[41681] <= 32'b11111111110000010000000100010011;
ROM[41682] <= 32'b00000000000000010010001110000011;
ROM[41683] <= 32'b00000000011100011010000000100011;
ROM[41684] <= 32'b00000000000000011010001110000011;
ROM[41685] <= 32'b00000000011100010010000000100011;
ROM[41686] <= 32'b00000000010000010000000100010011;
ROM[41687] <= 32'b00000000000000101001001110110111;
ROM[41688] <= 32'b10111010100000111000001110010011;
ROM[41689] <= 32'b00000000111000111000001110110011;
ROM[41690] <= 32'b00000000011100010010000000100011;
ROM[41691] <= 32'b00000000010000010000000100010011;
ROM[41692] <= 32'b00000000001100010010000000100011;
ROM[41693] <= 32'b00000000010000010000000100010011;
ROM[41694] <= 32'b00000000010000010010000000100011;
ROM[41695] <= 32'b00000000010000010000000100010011;
ROM[41696] <= 32'b00000000010100010010000000100011;
ROM[41697] <= 32'b00000000010000010000000100010011;
ROM[41698] <= 32'b00000000011000010010000000100011;
ROM[41699] <= 32'b00000000010000010000000100010011;
ROM[41700] <= 32'b00000001010000000000001110010011;
ROM[41701] <= 32'b00000000010000111000001110010011;
ROM[41702] <= 32'b01000000011100010000001110110011;
ROM[41703] <= 32'b00000000011100000000001000110011;
ROM[41704] <= 32'b00000000001000000000000110110011;
ROM[41705] <= 32'b10111100010011101110000011101111;
ROM[41706] <= 32'b11111111110000010000000100010011;
ROM[41707] <= 32'b00000000000000010010001110000011;
ROM[41708] <= 32'b00000000011101100010000000100011;
ROM[41709] <= 32'b00000000000000011010001110000011;
ROM[41710] <= 32'b00000000011100010010000000100011;
ROM[41711] <= 32'b00000000010000010000000100010011;
ROM[41712] <= 32'b00000000000000101001001110110111;
ROM[41713] <= 32'b11000000110000111000001110010011;
ROM[41714] <= 32'b00000000111000111000001110110011;
ROM[41715] <= 32'b00000000011100010010000000100011;
ROM[41716] <= 32'b00000000010000010000000100010011;
ROM[41717] <= 32'b00000000001100010010000000100011;
ROM[41718] <= 32'b00000000010000010000000100010011;
ROM[41719] <= 32'b00000000010000010010000000100011;
ROM[41720] <= 32'b00000000010000010000000100010011;
ROM[41721] <= 32'b00000000010100010010000000100011;
ROM[41722] <= 32'b00000000010000010000000100010011;
ROM[41723] <= 32'b00000000011000010010000000100011;
ROM[41724] <= 32'b00000000010000010000000100010011;
ROM[41725] <= 32'b00000001010000000000001110010011;
ROM[41726] <= 32'b00000000010000111000001110010011;
ROM[41727] <= 32'b01000000011100010000001110110011;
ROM[41728] <= 32'b00000000011100000000001000110011;
ROM[41729] <= 32'b00000000001000000000000110110011;
ROM[41730] <= 32'b00010000100000000010000011101111;
ROM[41731] <= 32'b11111111110000010000000100010011;
ROM[41732] <= 32'b00000000000000010010001110000011;
ROM[41733] <= 32'b00000000011101100010000000100011;
ROM[41734] <= 32'b00000000000000000000001110010011;
ROM[41735] <= 32'b00000000011100010010000000100011;
ROM[41736] <= 32'b00000000010000010000000100010011;
ROM[41737] <= 32'b00000001010000000000001110010011;
ROM[41738] <= 32'b01000000011100011000001110110011;
ROM[41739] <= 32'b00000000000000111010000010000011;
ROM[41740] <= 32'b11111111110000010000000100010011;
ROM[41741] <= 32'b00000000000000010010001110000011;
ROM[41742] <= 32'b00000000011100100010000000100011;
ROM[41743] <= 32'b00000000010000100000000100010011;
ROM[41744] <= 32'b00000001010000000000001110010011;
ROM[41745] <= 32'b01000000011100011000001110110011;
ROM[41746] <= 32'b00000000010000111010000110000011;
ROM[41747] <= 32'b00000000100000111010001000000011;
ROM[41748] <= 32'b00000000110000111010001010000011;
ROM[41749] <= 32'b00000001000000111010001100000011;
ROM[41750] <= 32'b00000000000000001000000011100111;
ROM[41751] <= 32'b00000000000000010010000000100011;
ROM[41752] <= 32'b00000000010000010000000100010011;
ROM[41753] <= 32'b00000000000000100010001110000011;
ROM[41754] <= 32'b00000000011100010010000000100011;
ROM[41755] <= 32'b00000000010000010000000100010011;
ROM[41756] <= 32'b11111111110000010000000100010011;
ROM[41757] <= 32'b00000000000000010010001110000011;
ROM[41758] <= 32'b00000000000000111000001010010011;
ROM[41759] <= 32'b00000001011000000000001110010011;
ROM[41760] <= 32'b00000000011100010010000000100011;
ROM[41761] <= 32'b00000000010000010000000100010011;
ROM[41762] <= 32'b00000000110000000000001110010011;
ROM[41763] <= 32'b00000000011100010010000000100011;
ROM[41764] <= 32'b00000000010000010000000100010011;
ROM[41765] <= 32'b00000000000000101001001110110111;
ROM[41766] <= 32'b11001110000000111000001110010011;
ROM[41767] <= 32'b00000000111000111000001110110011;
ROM[41768] <= 32'b00000000011100010010000000100011;
ROM[41769] <= 32'b00000000010000010000000100010011;
ROM[41770] <= 32'b00000000001100010010000000100011;
ROM[41771] <= 32'b00000000010000010000000100010011;
ROM[41772] <= 32'b00000000010000010010000000100011;
ROM[41773] <= 32'b00000000010000010000000100010011;
ROM[41774] <= 32'b00000000010100010010000000100011;
ROM[41775] <= 32'b00000000010000010000000100010011;
ROM[41776] <= 32'b00000000011000010010000000100011;
ROM[41777] <= 32'b00000000010000010000000100010011;
ROM[41778] <= 32'b00000001010000000000001110010011;
ROM[41779] <= 32'b00000000100000111000001110010011;
ROM[41780] <= 32'b01000000011100010000001110110011;
ROM[41781] <= 32'b00000000011100000000001000110011;
ROM[41782] <= 32'b00000000001000000000000110110011;
ROM[41783] <= 32'b11110010010111101100000011101111;
ROM[41784] <= 32'b11111111110000010000000100010011;
ROM[41785] <= 32'b00000000000000010010001110000011;
ROM[41786] <= 32'b00000000011101100010000000100011;
ROM[41787] <= 32'b00000000101100000000001110010011;
ROM[41788] <= 32'b00000000011100010010000000100011;
ROM[41789] <= 32'b00000000010000010000000100010011;
ROM[41790] <= 32'b00000000000000101001001110110111;
ROM[41791] <= 32'b11010100010000111000001110010011;
ROM[41792] <= 32'b00000000111000111000001110110011;
ROM[41793] <= 32'b00000000011100010010000000100011;
ROM[41794] <= 32'b00000000010000010000000100010011;
ROM[41795] <= 32'b00000000001100010010000000100011;
ROM[41796] <= 32'b00000000010000010000000100010011;
ROM[41797] <= 32'b00000000010000010010000000100011;
ROM[41798] <= 32'b00000000010000010000000100010011;
ROM[41799] <= 32'b00000000010100010010000000100011;
ROM[41800] <= 32'b00000000010000010000000100010011;
ROM[41801] <= 32'b00000000011000010010000000100011;
ROM[41802] <= 32'b00000000010000010000000100010011;
ROM[41803] <= 32'b00000001010000000000001110010011;
ROM[41804] <= 32'b00000000010000111000001110010011;
ROM[41805] <= 32'b01000000011100010000001110110011;
ROM[41806] <= 32'b00000000011100000000001000110011;
ROM[41807] <= 32'b00000000001000000000000110110011;
ROM[41808] <= 32'b00011111110100000000000011101111;
ROM[41809] <= 32'b00000010000000000000001110010011;
ROM[41810] <= 32'b00000000011100010010000000100011;
ROM[41811] <= 32'b00000000010000010000000100010011;
ROM[41812] <= 32'b00000000000000101001001110110111;
ROM[41813] <= 32'b11011001110000111000001110010011;
ROM[41814] <= 32'b00000000111000111000001110110011;
ROM[41815] <= 32'b00000000011100010010000000100011;
ROM[41816] <= 32'b00000000010000010000000100010011;
ROM[41817] <= 32'b00000000001100010010000000100011;
ROM[41818] <= 32'b00000000010000010000000100010011;
ROM[41819] <= 32'b00000000010000010010000000100011;
ROM[41820] <= 32'b00000000010000010000000100010011;
ROM[41821] <= 32'b00000000010100010010000000100011;
ROM[41822] <= 32'b00000000010000010000000100010011;
ROM[41823] <= 32'b00000000011000010010000000100011;
ROM[41824] <= 32'b00000000010000010000000100010011;
ROM[41825] <= 32'b00000001010000000000001110010011;
ROM[41826] <= 32'b00000000100000111000001110010011;
ROM[41827] <= 32'b01000000011100010000001110110011;
ROM[41828] <= 32'b00000000011100000000001000110011;
ROM[41829] <= 32'b00000000001000000000000110110011;
ROM[41830] <= 32'b01100001010100000000000011101111;
ROM[41831] <= 32'b00000101101100000000001110010011;
ROM[41832] <= 32'b00000000011100010010000000100011;
ROM[41833] <= 32'b00000000010000010000000100010011;
ROM[41834] <= 32'b00000000000000101001001110110111;
ROM[41835] <= 32'b11011111010000111000001110010011;
ROM[41836] <= 32'b00000000111000111000001110110011;
ROM[41837] <= 32'b00000000011100010010000000100011;
ROM[41838] <= 32'b00000000010000010000000100010011;
ROM[41839] <= 32'b00000000001100010010000000100011;
ROM[41840] <= 32'b00000000010000010000000100010011;
ROM[41841] <= 32'b00000000010000010010000000100011;
ROM[41842] <= 32'b00000000010000010000000100010011;
ROM[41843] <= 32'b00000000010100010010000000100011;
ROM[41844] <= 32'b00000000010000010000000100010011;
ROM[41845] <= 32'b00000000011000010010000000100011;
ROM[41846] <= 32'b00000000010000010000000100010011;
ROM[41847] <= 32'b00000001010000000000001110010011;
ROM[41848] <= 32'b00000000100000111000001110010011;
ROM[41849] <= 32'b01000000011100010000001110110011;
ROM[41850] <= 32'b00000000011100000000001000110011;
ROM[41851] <= 32'b00000000001000000000000110110011;
ROM[41852] <= 32'b01011011110100000000000011101111;
ROM[41853] <= 32'b00000100010000000000001110010011;
ROM[41854] <= 32'b00000000011100010010000000100011;
ROM[41855] <= 32'b00000000010000010000000100010011;
ROM[41856] <= 32'b00000000000000101001001110110111;
ROM[41857] <= 32'b11100100110000111000001110010011;
ROM[41858] <= 32'b00000000111000111000001110110011;
ROM[41859] <= 32'b00000000011100010010000000100011;
ROM[41860] <= 32'b00000000010000010000000100010011;
ROM[41861] <= 32'b00000000001100010010000000100011;
ROM[41862] <= 32'b00000000010000010000000100010011;
ROM[41863] <= 32'b00000000010000010010000000100011;
ROM[41864] <= 32'b00000000010000010000000100010011;
ROM[41865] <= 32'b00000000010100010010000000100011;
ROM[41866] <= 32'b00000000010000010000000100010011;
ROM[41867] <= 32'b00000000011000010010000000100011;
ROM[41868] <= 32'b00000000010000010000000100010011;
ROM[41869] <= 32'b00000001010000000000001110010011;
ROM[41870] <= 32'b00000000100000111000001110010011;
ROM[41871] <= 32'b01000000011100010000001110110011;
ROM[41872] <= 32'b00000000011100000000001000110011;
ROM[41873] <= 32'b00000000001000000000000110110011;
ROM[41874] <= 32'b01010110010100000000000011101111;
ROM[41875] <= 32'b00000100111100000000001110010011;
ROM[41876] <= 32'b00000000011100010010000000100011;
ROM[41877] <= 32'b00000000010000010000000100010011;
ROM[41878] <= 32'b00000000000000101001001110110111;
ROM[41879] <= 32'b11101010010000111000001110010011;
ROM[41880] <= 32'b00000000111000111000001110110011;
ROM[41881] <= 32'b00000000011100010010000000100011;
ROM[41882] <= 32'b00000000010000010000000100010011;
ROM[41883] <= 32'b00000000001100010010000000100011;
ROM[41884] <= 32'b00000000010000010000000100010011;
ROM[41885] <= 32'b00000000010000010010000000100011;
ROM[41886] <= 32'b00000000010000010000000100010011;
ROM[41887] <= 32'b00000000010100010010000000100011;
ROM[41888] <= 32'b00000000010000010000000100010011;
ROM[41889] <= 32'b00000000011000010010000000100011;
ROM[41890] <= 32'b00000000010000010000000100010011;
ROM[41891] <= 32'b00000001010000000000001110010011;
ROM[41892] <= 32'b00000000100000111000001110010011;
ROM[41893] <= 32'b01000000011100010000001110110011;
ROM[41894] <= 32'b00000000011100000000001000110011;
ROM[41895] <= 32'b00000000001000000000000110110011;
ROM[41896] <= 32'b01010000110100000000000011101111;
ROM[41897] <= 32'b00000100111000000000001110010011;
ROM[41898] <= 32'b00000000011100010010000000100011;
ROM[41899] <= 32'b00000000010000010000000100010011;
ROM[41900] <= 32'b00000000000000101001001110110111;
ROM[41901] <= 32'b11101111110000111000001110010011;
ROM[41902] <= 32'b00000000111000111000001110110011;
ROM[41903] <= 32'b00000000011100010010000000100011;
ROM[41904] <= 32'b00000000010000010000000100010011;
ROM[41905] <= 32'b00000000001100010010000000100011;
ROM[41906] <= 32'b00000000010000010000000100010011;
ROM[41907] <= 32'b00000000010000010010000000100011;
ROM[41908] <= 32'b00000000010000010000000100010011;
ROM[41909] <= 32'b00000000010100010010000000100011;
ROM[41910] <= 32'b00000000010000010000000100010011;
ROM[41911] <= 32'b00000000011000010010000000100011;
ROM[41912] <= 32'b00000000010000010000000100010011;
ROM[41913] <= 32'b00000001010000000000001110010011;
ROM[41914] <= 32'b00000000100000111000001110010011;
ROM[41915] <= 32'b01000000011100010000001110110011;
ROM[41916] <= 32'b00000000011100000000001000110011;
ROM[41917] <= 32'b00000000001000000000000110110011;
ROM[41918] <= 32'b01001011010100000000000011101111;
ROM[41919] <= 32'b00000100010100000000001110010011;
ROM[41920] <= 32'b00000000011100010010000000100011;
ROM[41921] <= 32'b00000000010000010000000100010011;
ROM[41922] <= 32'b00000000000000101001001110110111;
ROM[41923] <= 32'b11110101010000111000001110010011;
ROM[41924] <= 32'b00000000111000111000001110110011;
ROM[41925] <= 32'b00000000011100010010000000100011;
ROM[41926] <= 32'b00000000010000010000000100010011;
ROM[41927] <= 32'b00000000001100010010000000100011;
ROM[41928] <= 32'b00000000010000010000000100010011;
ROM[41929] <= 32'b00000000010000010010000000100011;
ROM[41930] <= 32'b00000000010000010000000100010011;
ROM[41931] <= 32'b00000000010100010010000000100011;
ROM[41932] <= 32'b00000000010000010000000100010011;
ROM[41933] <= 32'b00000000011000010010000000100011;
ROM[41934] <= 32'b00000000010000010000000100010011;
ROM[41935] <= 32'b00000001010000000000001110010011;
ROM[41936] <= 32'b00000000100000111000001110010011;
ROM[41937] <= 32'b01000000011100010000001110110011;
ROM[41938] <= 32'b00000000011100000000001000110011;
ROM[41939] <= 32'b00000000001000000000000110110011;
ROM[41940] <= 32'b01000101110100000000000011101111;
ROM[41941] <= 32'b00000010101000000000001110010011;
ROM[41942] <= 32'b00000000011100010010000000100011;
ROM[41943] <= 32'b00000000010000010000000100010011;
ROM[41944] <= 32'b00000000000000101001001110110111;
ROM[41945] <= 32'b11111010110000111000001110010011;
ROM[41946] <= 32'b00000000111000111000001110110011;
ROM[41947] <= 32'b00000000011100010010000000100011;
ROM[41948] <= 32'b00000000010000010000000100010011;
ROM[41949] <= 32'b00000000001100010010000000100011;
ROM[41950] <= 32'b00000000010000010000000100010011;
ROM[41951] <= 32'b00000000010000010010000000100011;
ROM[41952] <= 32'b00000000010000010000000100010011;
ROM[41953] <= 32'b00000000010100010010000000100011;
ROM[41954] <= 32'b00000000010000010000000100010011;
ROM[41955] <= 32'b00000000011000010010000000100011;
ROM[41956] <= 32'b00000000010000010000000100010011;
ROM[41957] <= 32'b00000001010000000000001110010011;
ROM[41958] <= 32'b00000000100000111000001110010011;
ROM[41959] <= 32'b01000000011100010000001110110011;
ROM[41960] <= 32'b00000000011100000000001000110011;
ROM[41961] <= 32'b00000000001000000000000110110011;
ROM[41962] <= 32'b01000000010100000000000011101111;
ROM[41963] <= 32'b00000011010000000000001110010011;
ROM[41964] <= 32'b00000000011100010010000000100011;
ROM[41965] <= 32'b00000000010000010000000100010011;
ROM[41966] <= 32'b00000000000000101001001110110111;
ROM[41967] <= 32'b00000000010000111000001110010011;
ROM[41968] <= 32'b00000000111000111000001110110011;
ROM[41969] <= 32'b00000000011100010010000000100011;
ROM[41970] <= 32'b00000000010000010000000100010011;
ROM[41971] <= 32'b00000000001100010010000000100011;
ROM[41972] <= 32'b00000000010000010000000100010011;
ROM[41973] <= 32'b00000000010000010010000000100011;
ROM[41974] <= 32'b00000000010000010000000100010011;
ROM[41975] <= 32'b00000000010100010010000000100011;
ROM[41976] <= 32'b00000000010000010000000100010011;
ROM[41977] <= 32'b00000000011000010010000000100011;
ROM[41978] <= 32'b00000000010000010000000100010011;
ROM[41979] <= 32'b00000001010000000000001110010011;
ROM[41980] <= 32'b00000000100000111000001110010011;
ROM[41981] <= 32'b01000000011100010000001110110011;
ROM[41982] <= 32'b00000000011100000000001000110011;
ROM[41983] <= 32'b00000000001000000000000110110011;
ROM[41984] <= 32'b00111010110100000000000011101111;
ROM[41985] <= 32'b00000101110100000000001110010011;
ROM[41986] <= 32'b00000000011100010010000000100011;
ROM[41987] <= 32'b00000000010000010000000100010011;
ROM[41988] <= 32'b00000000000000101001001110110111;
ROM[41989] <= 32'b00000101110000111000001110010011;
ROM[41990] <= 32'b00000000111000111000001110110011;
ROM[41991] <= 32'b00000000011100010010000000100011;
ROM[41992] <= 32'b00000000010000010000000100010011;
ROM[41993] <= 32'b00000000001100010010000000100011;
ROM[41994] <= 32'b00000000010000010000000100010011;
ROM[41995] <= 32'b00000000010000010010000000100011;
ROM[41996] <= 32'b00000000010000010000000100010011;
ROM[41997] <= 32'b00000000010100010010000000100011;
ROM[41998] <= 32'b00000000010000010000000100010011;
ROM[41999] <= 32'b00000000011000010010000000100011;
ROM[42000] <= 32'b00000000010000010000000100010011;
ROM[42001] <= 32'b00000001010000000000001110010011;
ROM[42002] <= 32'b00000000100000111000001110010011;
ROM[42003] <= 32'b01000000011100010000001110110011;
ROM[42004] <= 32'b00000000011100000000001000110011;
ROM[42005] <= 32'b00000000001000000000000110110011;
ROM[42006] <= 32'b00110101010100000000000011101111;
ROM[42007] <= 32'b00000010000000000000001110010011;
ROM[42008] <= 32'b00000000011100010010000000100011;
ROM[42009] <= 32'b00000000010000010000000100010011;
ROM[42010] <= 32'b00000000000000101001001110110111;
ROM[42011] <= 32'b00001011010000111000001110010011;
ROM[42012] <= 32'b00000000111000111000001110110011;
ROM[42013] <= 32'b00000000011100010010000000100011;
ROM[42014] <= 32'b00000000010000010000000100010011;
ROM[42015] <= 32'b00000000001100010010000000100011;
ROM[42016] <= 32'b00000000010000010000000100010011;
ROM[42017] <= 32'b00000000010000010010000000100011;
ROM[42018] <= 32'b00000000010000010000000100010011;
ROM[42019] <= 32'b00000000010100010010000000100011;
ROM[42020] <= 32'b00000000010000010000000100010011;
ROM[42021] <= 32'b00000000011000010010000000100011;
ROM[42022] <= 32'b00000000010000010000000100010011;
ROM[42023] <= 32'b00000001010000000000001110010011;
ROM[42024] <= 32'b00000000100000111000001110010011;
ROM[42025] <= 32'b01000000011100010000001110110011;
ROM[42026] <= 32'b00000000011100000000001000110011;
ROM[42027] <= 32'b00000000001000000000000110110011;
ROM[42028] <= 32'b00101111110100000000000011101111;
ROM[42029] <= 32'b00000010000000000000001110010011;
ROM[42030] <= 32'b00000000011100010010000000100011;
ROM[42031] <= 32'b00000000010000010000000100010011;
ROM[42032] <= 32'b00000000000000101001001110110111;
ROM[42033] <= 32'b00010000110000111000001110010011;
ROM[42034] <= 32'b00000000111000111000001110110011;
ROM[42035] <= 32'b00000000011100010010000000100011;
ROM[42036] <= 32'b00000000010000010000000100010011;
ROM[42037] <= 32'b00000000001100010010000000100011;
ROM[42038] <= 32'b00000000010000010000000100010011;
ROM[42039] <= 32'b00000000010000010010000000100011;
ROM[42040] <= 32'b00000000010000010000000100010011;
ROM[42041] <= 32'b00000000010100010010000000100011;
ROM[42042] <= 32'b00000000010000010000000100010011;
ROM[42043] <= 32'b00000000011000010010000000100011;
ROM[42044] <= 32'b00000000010000010000000100010011;
ROM[42045] <= 32'b00000001010000000000001110010011;
ROM[42046] <= 32'b00000000100000111000001110010011;
ROM[42047] <= 32'b01000000011100010000001110110011;
ROM[42048] <= 32'b00000000011100000000001000110011;
ROM[42049] <= 32'b00000000001000000000000110110011;
ROM[42050] <= 32'b00101010010100000000000011101111;
ROM[42051] <= 32'b11111111110000010000000100010011;
ROM[42052] <= 32'b00000000000000010010001110000011;
ROM[42053] <= 32'b00000000011100011010000000100011;
ROM[42054] <= 32'b00000000000000011010001110000011;
ROM[42055] <= 32'b00000000011100010010000000100011;
ROM[42056] <= 32'b00000000010000010000000100010011;
ROM[42057] <= 32'b00000000000000101001001110110111;
ROM[42058] <= 32'b00010111000000111000001110010011;
ROM[42059] <= 32'b00000000111000111000001110110011;
ROM[42060] <= 32'b00000000011100010010000000100011;
ROM[42061] <= 32'b00000000010000010000000100010011;
ROM[42062] <= 32'b00000000001100010010000000100011;
ROM[42063] <= 32'b00000000010000010000000100010011;
ROM[42064] <= 32'b00000000010000010010000000100011;
ROM[42065] <= 32'b00000000010000010000000100010011;
ROM[42066] <= 32'b00000000010100010010000000100011;
ROM[42067] <= 32'b00000000010000010000000100010011;
ROM[42068] <= 32'b00000000011000010010000000100011;
ROM[42069] <= 32'b00000000010000010000000100010011;
ROM[42070] <= 32'b00000001010000000000001110010011;
ROM[42071] <= 32'b00000000010000111000001110010011;
ROM[42072] <= 32'b01000000011100010000001110110011;
ROM[42073] <= 32'b00000000011100000000001000110011;
ROM[42074] <= 32'b00000000001000000000000110110011;
ROM[42075] <= 32'b11011111110111101101000011101111;
ROM[42076] <= 32'b11111111110000010000000100010011;
ROM[42077] <= 32'b00000000000000010010001110000011;
ROM[42078] <= 32'b00000000011101100010000000100011;
ROM[42079] <= 32'b00000000000000011010001110000011;
ROM[42080] <= 32'b00000000011100010010000000100011;
ROM[42081] <= 32'b00000000010000010000000100010011;
ROM[42082] <= 32'b00000000000000101001001110110111;
ROM[42083] <= 32'b00011101010000111000001110010011;
ROM[42084] <= 32'b00000000111000111000001110110011;
ROM[42085] <= 32'b00000000011100010010000000100011;
ROM[42086] <= 32'b00000000010000010000000100010011;
ROM[42087] <= 32'b00000000001100010010000000100011;
ROM[42088] <= 32'b00000000010000010000000100010011;
ROM[42089] <= 32'b00000000010000010010000000100011;
ROM[42090] <= 32'b00000000010000010000000100010011;
ROM[42091] <= 32'b00000000010100010010000000100011;
ROM[42092] <= 32'b00000000010000010000000100010011;
ROM[42093] <= 32'b00000000011000010010000000100011;
ROM[42094] <= 32'b00000000010000010000000100010011;
ROM[42095] <= 32'b00000001010000000000001110010011;
ROM[42096] <= 32'b00000000010000111000001110010011;
ROM[42097] <= 32'b01000000011100010000001110110011;
ROM[42098] <= 32'b00000000011100000000001000110011;
ROM[42099] <= 32'b00000000001000000000000110110011;
ROM[42100] <= 32'b00110100000100000001000011101111;
ROM[42101] <= 32'b11111111110000010000000100010011;
ROM[42102] <= 32'b00000000000000010010001110000011;
ROM[42103] <= 32'b00000000011101100010000000100011;
ROM[42104] <= 32'b00000000000000000000001110010011;
ROM[42105] <= 32'b00000000011100010010000000100011;
ROM[42106] <= 32'b00000000010000010000000100010011;
ROM[42107] <= 32'b00000001010000000000001110010011;
ROM[42108] <= 32'b01000000011100011000001110110011;
ROM[42109] <= 32'b00000000000000111010000010000011;
ROM[42110] <= 32'b11111111110000010000000100010011;
ROM[42111] <= 32'b00000000000000010010001110000011;
ROM[42112] <= 32'b00000000011100100010000000100011;
ROM[42113] <= 32'b00000000010000100000000100010011;
ROM[42114] <= 32'b00000001010000000000001110010011;
ROM[42115] <= 32'b01000000011100011000001110110011;
ROM[42116] <= 32'b00000000010000111010000110000011;
ROM[42117] <= 32'b00000000100000111010001000000011;
ROM[42118] <= 32'b00000000110000111010001010000011;
ROM[42119] <= 32'b00000001000000111010001100000011;
ROM[42120] <= 32'b00000000000000001000000011100111;
ROM[42121] <= 32'b00000000000000010010000000100011;
ROM[42122] <= 32'b00000000010000010000000100010011;
ROM[42123] <= 32'b00000000000000100010001110000011;
ROM[42124] <= 32'b00000000011100010010000000100011;
ROM[42125] <= 32'b00000000010000010000000100010011;
ROM[42126] <= 32'b11111111110000010000000100010011;
ROM[42127] <= 32'b00000000000000010010001110000011;
ROM[42128] <= 32'b00000000000000111000001010010011;
ROM[42129] <= 32'b00000001011000000000001110010011;
ROM[42130] <= 32'b00000000011100010010000000100011;
ROM[42131] <= 32'b00000000010000010000000100010011;
ROM[42132] <= 32'b00000000110000000000001110010011;
ROM[42133] <= 32'b00000000011100010010000000100011;
ROM[42134] <= 32'b00000000010000010000000100010011;
ROM[42135] <= 32'b00000000000000101001001110110111;
ROM[42136] <= 32'b00101010100000111000001110010011;
ROM[42137] <= 32'b00000000111000111000001110110011;
ROM[42138] <= 32'b00000000011100010010000000100011;
ROM[42139] <= 32'b00000000010000010000000100010011;
ROM[42140] <= 32'b00000000001100010010000000100011;
ROM[42141] <= 32'b00000000010000010000000100010011;
ROM[42142] <= 32'b00000000010000010010000000100011;
ROM[42143] <= 32'b00000000010000010000000100010011;
ROM[42144] <= 32'b00000000010100010010000000100011;
ROM[42145] <= 32'b00000000010000010000000100010011;
ROM[42146] <= 32'b00000000011000010010000000100011;
ROM[42147] <= 32'b00000000010000010000000100010011;
ROM[42148] <= 32'b00000001010000000000001110010011;
ROM[42149] <= 32'b00000000100000111000001110010011;
ROM[42150] <= 32'b01000000011100010000001110110011;
ROM[42151] <= 32'b00000000011100000000001000110011;
ROM[42152] <= 32'b00000000001000000000000110110011;
ROM[42153] <= 32'b10010101110111101100000011101111;
ROM[42154] <= 32'b11111111110000010000000100010011;
ROM[42155] <= 32'b00000000000000010010001110000011;
ROM[42156] <= 32'b00000000011101100010000000100011;
ROM[42157] <= 32'b00000000100100000000001110010011;
ROM[42158] <= 32'b00000000011100010010000000100011;
ROM[42159] <= 32'b00000000010000010000000100010011;
ROM[42160] <= 32'b00000000000000101001001110110111;
ROM[42161] <= 32'b00110000110000111000001110010011;
ROM[42162] <= 32'b00000000111000111000001110110011;
ROM[42163] <= 32'b00000000011100010010000000100011;
ROM[42164] <= 32'b00000000010000010000000100010011;
ROM[42165] <= 32'b00000000001100010010000000100011;
ROM[42166] <= 32'b00000000010000010000000100010011;
ROM[42167] <= 32'b00000000010000010010000000100011;
ROM[42168] <= 32'b00000000010000010000000100010011;
ROM[42169] <= 32'b00000000010100010010000000100011;
ROM[42170] <= 32'b00000000010000010000000100010011;
ROM[42171] <= 32'b00000000011000010010000000100011;
ROM[42172] <= 32'b00000000010000010000000100010011;
ROM[42173] <= 32'b00000001010000000000001110010011;
ROM[42174] <= 32'b00000000010000111000001110010011;
ROM[42175] <= 32'b01000000011100010000001110110011;
ROM[42176] <= 32'b00000000011100000000001000110011;
ROM[42177] <= 32'b00000000001000000000000110110011;
ROM[42178] <= 32'b01000011010000000000000011101111;
ROM[42179] <= 32'b00000010101000000000001110010011;
ROM[42180] <= 32'b00000000011100010010000000100011;
ROM[42181] <= 32'b00000000010000010000000100010011;
ROM[42182] <= 32'b00000000000000101001001110110111;
ROM[42183] <= 32'b00110110010000111000001110010011;
ROM[42184] <= 32'b00000000111000111000001110110011;
ROM[42185] <= 32'b00000000011100010010000000100011;
ROM[42186] <= 32'b00000000010000010000000100010011;
ROM[42187] <= 32'b00000000001100010010000000100011;
ROM[42188] <= 32'b00000000010000010000000100010011;
ROM[42189] <= 32'b00000000010000010010000000100011;
ROM[42190] <= 32'b00000000010000010000000100010011;
ROM[42191] <= 32'b00000000010100010010000000100011;
ROM[42192] <= 32'b00000000010000010000000100010011;
ROM[42193] <= 32'b00000000011000010010000000100011;
ROM[42194] <= 32'b00000000010000010000000100010011;
ROM[42195] <= 32'b00000001010000000000001110010011;
ROM[42196] <= 32'b00000000100000111000001110010011;
ROM[42197] <= 32'b01000000011100010000001110110011;
ROM[42198] <= 32'b00000000011100000000001000110011;
ROM[42199] <= 32'b00000000001000000000000110110011;
ROM[42200] <= 32'b00000100110100000000000011101111;
ROM[42201] <= 32'b00000100001100000000001110010011;
ROM[42202] <= 32'b00000000011100010010000000100011;
ROM[42203] <= 32'b00000000010000010000000100010011;
ROM[42204] <= 32'b00000000000000101001001110110111;
ROM[42205] <= 32'b00111011110000111000001110010011;
ROM[42206] <= 32'b00000000111000111000001110110011;
ROM[42207] <= 32'b00000000011100010010000000100011;
ROM[42208] <= 32'b00000000010000010000000100010011;
ROM[42209] <= 32'b00000000001100010010000000100011;
ROM[42210] <= 32'b00000000010000010000000100010011;
ROM[42211] <= 32'b00000000010000010010000000100011;
ROM[42212] <= 32'b00000000010000010000000100010011;
ROM[42213] <= 32'b00000000010100010010000000100011;
ROM[42214] <= 32'b00000000010000010000000100010011;
ROM[42215] <= 32'b00000000011000010010000000100011;
ROM[42216] <= 32'b00000000010000010000000100010011;
ROM[42217] <= 32'b00000001010000000000001110010011;
ROM[42218] <= 32'b00000000100000111000001110010011;
ROM[42219] <= 32'b01000000011100010000001110110011;
ROM[42220] <= 32'b00000000011100000000001000110011;
ROM[42221] <= 32'b00000000001000000000000110110011;
ROM[42222] <= 32'b01111111010000000000000011101111;
ROM[42223] <= 32'b00000101001000000000001110010011;
ROM[42224] <= 32'b00000000011100010010000000100011;
ROM[42225] <= 32'b00000000010000010000000100010011;
ROM[42226] <= 32'b00000000000000101001001110110111;
ROM[42227] <= 32'b01000001010000111000001110010011;
ROM[42228] <= 32'b00000000111000111000001110110011;
ROM[42229] <= 32'b00000000011100010010000000100011;
ROM[42230] <= 32'b00000000010000010000000100010011;
ROM[42231] <= 32'b00000000001100010010000000100011;
ROM[42232] <= 32'b00000000010000010000000100010011;
ROM[42233] <= 32'b00000000010000010010000000100011;
ROM[42234] <= 32'b00000000010000010000000100010011;
ROM[42235] <= 32'b00000000010100010010000000100011;
ROM[42236] <= 32'b00000000010000010000000100010011;
ROM[42237] <= 32'b00000000011000010010000000100011;
ROM[42238] <= 32'b00000000010000010000000100010011;
ROM[42239] <= 32'b00000001010000000000001110010011;
ROM[42240] <= 32'b00000000100000111000001110010011;
ROM[42241] <= 32'b01000000011100010000001110110011;
ROM[42242] <= 32'b00000000011100000000001000110011;
ROM[42243] <= 32'b00000000001000000000000110110011;
ROM[42244] <= 32'b01111001110000000000000011101111;
ROM[42245] <= 32'b00000100000100000000001110010011;
ROM[42246] <= 32'b00000000011100010010000000100011;
ROM[42247] <= 32'b00000000010000010000000100010011;
ROM[42248] <= 32'b00000000000000101001001110110111;
ROM[42249] <= 32'b01000110110000111000001110010011;
ROM[42250] <= 32'b00000000111000111000001110110011;
ROM[42251] <= 32'b00000000011100010010000000100011;
ROM[42252] <= 32'b00000000010000010000000100010011;
ROM[42253] <= 32'b00000000001100010010000000100011;
ROM[42254] <= 32'b00000000010000010000000100010011;
ROM[42255] <= 32'b00000000010000010010000000100011;
ROM[42256] <= 32'b00000000010000010000000100010011;
ROM[42257] <= 32'b00000000010100010010000000100011;
ROM[42258] <= 32'b00000000010000010000000100010011;
ROM[42259] <= 32'b00000000011000010010000000100011;
ROM[42260] <= 32'b00000000010000010000000100010011;
ROM[42261] <= 32'b00000001010000000000001110010011;
ROM[42262] <= 32'b00000000100000111000001110010011;
ROM[42263] <= 32'b01000000011100010000001110110011;
ROM[42264] <= 32'b00000000011100000000001000110011;
ROM[42265] <= 32'b00000000001000000000000110110011;
ROM[42266] <= 32'b01110100010000000000000011101111;
ROM[42267] <= 32'b00000101001100000000001110010011;
ROM[42268] <= 32'b00000000011100010010000000100011;
ROM[42269] <= 32'b00000000010000010000000100010011;
ROM[42270] <= 32'b00000000000000101001001110110111;
ROM[42271] <= 32'b01001100010000111000001110010011;
ROM[42272] <= 32'b00000000111000111000001110110011;
ROM[42273] <= 32'b00000000011100010010000000100011;
ROM[42274] <= 32'b00000000010000010000000100010011;
ROM[42275] <= 32'b00000000001100010010000000100011;
ROM[42276] <= 32'b00000000010000010000000100010011;
ROM[42277] <= 32'b00000000010000010010000000100011;
ROM[42278] <= 32'b00000000010000010000000100010011;
ROM[42279] <= 32'b00000000010100010010000000100011;
ROM[42280] <= 32'b00000000010000010000000100010011;
ROM[42281] <= 32'b00000000011000010010000000100011;
ROM[42282] <= 32'b00000000010000010000000100010011;
ROM[42283] <= 32'b00000001010000000000001110010011;
ROM[42284] <= 32'b00000000100000111000001110010011;
ROM[42285] <= 32'b01000000011100010000001110110011;
ROM[42286] <= 32'b00000000011100000000001000110011;
ROM[42287] <= 32'b00000000001000000000000110110011;
ROM[42288] <= 32'b01101110110000000000000011101111;
ROM[42289] <= 32'b00000100100000000000001110010011;
ROM[42290] <= 32'b00000000011100010010000000100011;
ROM[42291] <= 32'b00000000010000010000000100010011;
ROM[42292] <= 32'b00000000000000101001001110110111;
ROM[42293] <= 32'b01010001110000111000001110010011;
ROM[42294] <= 32'b00000000111000111000001110110011;
ROM[42295] <= 32'b00000000011100010010000000100011;
ROM[42296] <= 32'b00000000010000010000000100010011;
ROM[42297] <= 32'b00000000001100010010000000100011;
ROM[42298] <= 32'b00000000010000010000000100010011;
ROM[42299] <= 32'b00000000010000010010000000100011;
ROM[42300] <= 32'b00000000010000010000000100010011;
ROM[42301] <= 32'b00000000010100010010000000100011;
ROM[42302] <= 32'b00000000010000010000000100010011;
ROM[42303] <= 32'b00000000011000010010000000100011;
ROM[42304] <= 32'b00000000010000010000000100010011;
ROM[42305] <= 32'b00000001010000000000001110010011;
ROM[42306] <= 32'b00000000100000111000001110010011;
ROM[42307] <= 32'b01000000011100010000001110110011;
ROM[42308] <= 32'b00000000011100000000001000110011;
ROM[42309] <= 32'b00000000001000000000000110110011;
ROM[42310] <= 32'b01101001010000000000000011101111;
ROM[42311] <= 32'b00000100010100000000001110010011;
ROM[42312] <= 32'b00000000011100010010000000100011;
ROM[42313] <= 32'b00000000010000010000000100010011;
ROM[42314] <= 32'b00000000000000101001001110110111;
ROM[42315] <= 32'b01010111010000111000001110010011;
ROM[42316] <= 32'b00000000111000111000001110110011;
ROM[42317] <= 32'b00000000011100010010000000100011;
ROM[42318] <= 32'b00000000010000010000000100010011;
ROM[42319] <= 32'b00000000001100010010000000100011;
ROM[42320] <= 32'b00000000010000010000000100010011;
ROM[42321] <= 32'b00000000010000010010000000100011;
ROM[42322] <= 32'b00000000010000010000000100010011;
ROM[42323] <= 32'b00000000010100010010000000100011;
ROM[42324] <= 32'b00000000010000010000000100010011;
ROM[42325] <= 32'b00000000011000010010000000100011;
ROM[42326] <= 32'b00000000010000010000000100010011;
ROM[42327] <= 32'b00000001010000000000001110010011;
ROM[42328] <= 32'b00000000100000111000001110010011;
ROM[42329] <= 32'b01000000011100010000001110110011;
ROM[42330] <= 32'b00000000011100000000001000110011;
ROM[42331] <= 32'b00000000001000000000000110110011;
ROM[42332] <= 32'b01100011110000000000000011101111;
ROM[42333] <= 32'b00000100010000000000001110010011;
ROM[42334] <= 32'b00000000011100010010000000100011;
ROM[42335] <= 32'b00000000010000010000000100010011;
ROM[42336] <= 32'b00000000000000101001001110110111;
ROM[42337] <= 32'b01011100110000111000001110010011;
ROM[42338] <= 32'b00000000111000111000001110110011;
ROM[42339] <= 32'b00000000011100010010000000100011;
ROM[42340] <= 32'b00000000010000010000000100010011;
ROM[42341] <= 32'b00000000001100010010000000100011;
ROM[42342] <= 32'b00000000010000010000000100010011;
ROM[42343] <= 32'b00000000010000010010000000100011;
ROM[42344] <= 32'b00000000010000010000000100010011;
ROM[42345] <= 32'b00000000010100010010000000100011;
ROM[42346] <= 32'b00000000010000010000000100010011;
ROM[42347] <= 32'b00000000011000010010000000100011;
ROM[42348] <= 32'b00000000010000010000000100010011;
ROM[42349] <= 32'b00000001010000000000001110010011;
ROM[42350] <= 32'b00000000100000111000001110010011;
ROM[42351] <= 32'b01000000011100010000001110110011;
ROM[42352] <= 32'b00000000011100000000001000110011;
ROM[42353] <= 32'b00000000001000000000000110110011;
ROM[42354] <= 32'b01011110010000000000000011101111;
ROM[42355] <= 32'b00000010101000000000001110010011;
ROM[42356] <= 32'b00000000011100010010000000100011;
ROM[42357] <= 32'b00000000010000010000000100010011;
ROM[42358] <= 32'b00000000000000101001001110110111;
ROM[42359] <= 32'b01100010010000111000001110010011;
ROM[42360] <= 32'b00000000111000111000001110110011;
ROM[42361] <= 32'b00000000011100010010000000100011;
ROM[42362] <= 32'b00000000010000010000000100010011;
ROM[42363] <= 32'b00000000001100010010000000100011;
ROM[42364] <= 32'b00000000010000010000000100010011;
ROM[42365] <= 32'b00000000010000010010000000100011;
ROM[42366] <= 32'b00000000010000010000000100010011;
ROM[42367] <= 32'b00000000010100010010000000100011;
ROM[42368] <= 32'b00000000010000010000000100010011;
ROM[42369] <= 32'b00000000011000010010000000100011;
ROM[42370] <= 32'b00000000010000010000000100010011;
ROM[42371] <= 32'b00000001010000000000001110010011;
ROM[42372] <= 32'b00000000100000111000001110010011;
ROM[42373] <= 32'b01000000011100010000001110110011;
ROM[42374] <= 32'b00000000011100000000001000110011;
ROM[42375] <= 32'b00000000001000000000000110110011;
ROM[42376] <= 32'b01011000110000000000000011101111;
ROM[42377] <= 32'b11111111110000010000000100010011;
ROM[42378] <= 32'b00000000000000010010001110000011;
ROM[42379] <= 32'b00000000011100011010000000100011;
ROM[42380] <= 32'b00000000000000011010001110000011;
ROM[42381] <= 32'b00000000011100010010000000100011;
ROM[42382] <= 32'b00000000010000010000000100010011;
ROM[42383] <= 32'b00000000000000101001001110110111;
ROM[42384] <= 32'b01101000100000111000001110010011;
ROM[42385] <= 32'b00000000111000111000001110110011;
ROM[42386] <= 32'b00000000011100010010000000100011;
ROM[42387] <= 32'b00000000010000010000000100010011;
ROM[42388] <= 32'b00000000001100010010000000100011;
ROM[42389] <= 32'b00000000010000010000000100010011;
ROM[42390] <= 32'b00000000010000010010000000100011;
ROM[42391] <= 32'b00000000010000010000000100010011;
ROM[42392] <= 32'b00000000010100010010000000100011;
ROM[42393] <= 32'b00000000010000010000000100010011;
ROM[42394] <= 32'b00000000011000010010000000100011;
ROM[42395] <= 32'b00000000010000010000000100010011;
ROM[42396] <= 32'b00000001010000000000001110010011;
ROM[42397] <= 32'b00000000010000111000001110010011;
ROM[42398] <= 32'b01000000011100010000001110110011;
ROM[42399] <= 32'b00000000011100000000001000110011;
ROM[42400] <= 32'b00000000001000000000000110110011;
ROM[42401] <= 32'b10001110010111101101000011101111;
ROM[42402] <= 32'b11111111110000010000000100010011;
ROM[42403] <= 32'b00000000000000010010001110000011;
ROM[42404] <= 32'b00000000011101100010000000100011;
ROM[42405] <= 32'b00000000000000011010001110000011;
ROM[42406] <= 32'b00000000011100010010000000100011;
ROM[42407] <= 32'b00000000010000010000000100010011;
ROM[42408] <= 32'b00000000000000101001001110110111;
ROM[42409] <= 32'b01101110110000111000001110010011;
ROM[42410] <= 32'b00000000111000111000001110110011;
ROM[42411] <= 32'b00000000011100010010000000100011;
ROM[42412] <= 32'b00000000010000010000000100010011;
ROM[42413] <= 32'b00000000001100010010000000100011;
ROM[42414] <= 32'b00000000010000010000000100010011;
ROM[42415] <= 32'b00000000010000010010000000100011;
ROM[42416] <= 32'b00000000010000010000000100010011;
ROM[42417] <= 32'b00000000010100010010000000100011;
ROM[42418] <= 32'b00000000010000010000000100010011;
ROM[42419] <= 32'b00000000011000010010000000100011;
ROM[42420] <= 32'b00000000010000010000000100010011;
ROM[42421] <= 32'b00000001010000000000001110010011;
ROM[42422] <= 32'b00000000010000111000001110010011;
ROM[42423] <= 32'b01000000011100010000001110110011;
ROM[42424] <= 32'b00000000011100000000001000110011;
ROM[42425] <= 32'b00000000001000000000000110110011;
ROM[42426] <= 32'b01100010100000000001000011101111;
ROM[42427] <= 32'b11111111110000010000000100010011;
ROM[42428] <= 32'b00000000000000010010001110000011;
ROM[42429] <= 32'b00000000011101100010000000100011;
ROM[42430] <= 32'b00000000000000000000001110010011;
ROM[42431] <= 32'b00000000011100010010000000100011;
ROM[42432] <= 32'b00000000010000010000000100010011;
ROM[42433] <= 32'b00000001010000000000001110010011;
ROM[42434] <= 32'b01000000011100011000001110110011;
ROM[42435] <= 32'b00000000000000111010000010000011;
ROM[42436] <= 32'b11111111110000010000000100010011;
ROM[42437] <= 32'b00000000000000010010001110000011;
ROM[42438] <= 32'b00000000011100100010000000100011;
ROM[42439] <= 32'b00000000010000100000000100010011;
ROM[42440] <= 32'b00000001010000000000001110010011;
ROM[42441] <= 32'b01000000011100011000001110110011;
ROM[42442] <= 32'b00000000010000111010000110000011;
ROM[42443] <= 32'b00000000100000111010001000000011;
ROM[42444] <= 32'b00000000110000111010001010000011;
ROM[42445] <= 32'b00000001000000111010001100000011;
ROM[42446] <= 32'b00000000000000001000000011100111;
ROM[42447] <= 32'b00000000001100000000001110010011;
ROM[42448] <= 32'b00000000011100010010000000100011;
ROM[42449] <= 32'b00000000010000010000000100010011;
ROM[42450] <= 32'b00000000000000101001001110110111;
ROM[42451] <= 32'b01111001010000111000001110010011;
ROM[42452] <= 32'b00000000111000111000001110110011;
ROM[42453] <= 32'b00000000011100010010000000100011;
ROM[42454] <= 32'b00000000010000010000000100010011;
ROM[42455] <= 32'b00000000001100010010000000100011;
ROM[42456] <= 32'b00000000010000010000000100010011;
ROM[42457] <= 32'b00000000010000010010000000100011;
ROM[42458] <= 32'b00000000010000010000000100010011;
ROM[42459] <= 32'b00000000010100010010000000100011;
ROM[42460] <= 32'b00000000010000010000000100010011;
ROM[42461] <= 32'b00000000011000010010000000100011;
ROM[42462] <= 32'b00000000010000010000000100010011;
ROM[42463] <= 32'b00000001010000000000001110010011;
ROM[42464] <= 32'b00000000010000111000001110010011;
ROM[42465] <= 32'b01000000011100010000001110110011;
ROM[42466] <= 32'b00000000011100000000001000110011;
ROM[42467] <= 32'b00000000001000000000000110110011;
ROM[42468] <= 32'b11110100010111101010000011101111;
ROM[42469] <= 32'b11111111110000010000000100010011;
ROM[42470] <= 32'b00000000000000010010001110000011;
ROM[42471] <= 32'b00000000000000111000001010010011;
ROM[42472] <= 32'b00000000000000100010001110000011;
ROM[42473] <= 32'b00000000011100010010000000100011;
ROM[42474] <= 32'b00000000010000010000000100010011;
ROM[42475] <= 32'b00000000000000000000001110010011;
ROM[42476] <= 32'b00000000011100010010000000100011;
ROM[42477] <= 32'b00000000010000010000000100010011;
ROM[42478] <= 32'b11111111110000010000000100010011;
ROM[42479] <= 32'b00000000000000010010001110000011;
ROM[42480] <= 32'b11111111110000010000000100010011;
ROM[42481] <= 32'b00000000000000010010010000000011;
ROM[42482] <= 32'b00000000011101000010010010110011;
ROM[42483] <= 32'b00000000100000111010010100110011;
ROM[42484] <= 32'b00000000101001001000001110110011;
ROM[42485] <= 32'b00000000000100111000001110010011;
ROM[42486] <= 32'b00000000000100111111001110010011;
ROM[42487] <= 32'b00000000011100010010000000100011;
ROM[42488] <= 32'b00000000010000010000000100010011;
ROM[42489] <= 32'b11111111110000010000000100010011;
ROM[42490] <= 32'b00000000000000010010001110000011;
ROM[42491] <= 32'b00000000000000111000101001100011;
ROM[42492] <= 32'b00000000000000101010001110110111;
ROM[42493] <= 32'b10000000010000111000001110010011;
ROM[42494] <= 32'b00000000111000111000001110110011;
ROM[42495] <= 32'b00000000000000111000000011100111;
ROM[42496] <= 32'b00000001110000000000000011101111;
ROM[42497] <= 32'b00000000000100000000001110010011;
ROM[42498] <= 32'b00000000011100010010000000100011;
ROM[42499] <= 32'b00000000010000010000000100010011;
ROM[42500] <= 32'b11111111110000010000000100010011;
ROM[42501] <= 32'b00000000000000010010001110000011;
ROM[42502] <= 32'b00000000011100100010000000100011;
ROM[42503] <= 32'b00000000000000000000001110010011;
ROM[42504] <= 32'b00000000011100010010000000100011;
ROM[42505] <= 32'b00000000010000010000000100010011;
ROM[42506] <= 32'b11111111110000010000000100010011;
ROM[42507] <= 32'b00000000000000010010001110000011;
ROM[42508] <= 32'b00000000110100101000010000110011;
ROM[42509] <= 32'b00000000011101000010001000100011;
ROM[42510] <= 32'b00000000000000100010001110000011;
ROM[42511] <= 32'b00000000011100010010000000100011;
ROM[42512] <= 32'b00000000010000010000000100010011;
ROM[42513] <= 32'b11111111110000010000000100010011;
ROM[42514] <= 32'b00000000000000010010001110000011;
ROM[42515] <= 32'b00000000110100101000010000110011;
ROM[42516] <= 32'b00000000011101000010000000100011;
ROM[42517] <= 32'b00000000000000100010001110000011;
ROM[42518] <= 32'b00000000011100010010000000100011;
ROM[42519] <= 32'b00000000010000010000000100010011;
ROM[42520] <= 32'b00000000000000101010001110110111;
ROM[42521] <= 32'b10001010110000111000001110010011;
ROM[42522] <= 32'b00000000111000111000001110110011;
ROM[42523] <= 32'b00000000011100010010000000100011;
ROM[42524] <= 32'b00000000010000010000000100010011;
ROM[42525] <= 32'b00000000001100010010000000100011;
ROM[42526] <= 32'b00000000010000010000000100010011;
ROM[42527] <= 32'b00000000010000010010000000100011;
ROM[42528] <= 32'b00000000010000010000000100010011;
ROM[42529] <= 32'b00000000010100010010000000100011;
ROM[42530] <= 32'b00000000010000010000000100010011;
ROM[42531] <= 32'b00000000011000010010000000100011;
ROM[42532] <= 32'b00000000010000010000000100010011;
ROM[42533] <= 32'b00000001010000000000001110010011;
ROM[42534] <= 32'b00000000010000111000001110010011;
ROM[42535] <= 32'b01000000011100010000001110110011;
ROM[42536] <= 32'b00000000011100000000001000110011;
ROM[42537] <= 32'b00000000001000000000000110110011;
ROM[42538] <= 32'b11111101100011010110000011101111;
ROM[42539] <= 32'b11111111110000010000000100010011;
ROM[42540] <= 32'b00000000000000010010001110000011;
ROM[42541] <= 32'b00000000110100101000010000110011;
ROM[42542] <= 32'b00000000011101000010010000100011;
ROM[42543] <= 32'b00000000010100010010000000100011;
ROM[42544] <= 32'b00000000010000010000000100010011;
ROM[42545] <= 32'b00000001010000000000001110010011;
ROM[42546] <= 32'b01000000011100011000001110110011;
ROM[42547] <= 32'b00000000000000111010000010000011;
ROM[42548] <= 32'b11111111110000010000000100010011;
ROM[42549] <= 32'b00000000000000010010001110000011;
ROM[42550] <= 32'b00000000011100100010000000100011;
ROM[42551] <= 32'b00000000010000100000000100010011;
ROM[42552] <= 32'b00000001010000000000001110010011;
ROM[42553] <= 32'b01000000011100011000001110110011;
ROM[42554] <= 32'b00000000010000111010000110000011;
ROM[42555] <= 32'b00000000100000111010001000000011;
ROM[42556] <= 32'b00000000110000111010001010000011;
ROM[42557] <= 32'b00000001000000111010001100000011;
ROM[42558] <= 32'b00000000000000001000000011100111;
ROM[42559] <= 32'b00000000000000100010001110000011;
ROM[42560] <= 32'b00000000011100010010000000100011;
ROM[42561] <= 32'b00000000010000010000000100010011;
ROM[42562] <= 32'b11111111110000010000000100010011;
ROM[42563] <= 32'b00000000000000010010001110000011;
ROM[42564] <= 32'b00000000000000111000001010010011;
ROM[42565] <= 32'b00000000110100101000010000110011;
ROM[42566] <= 32'b00000000010001000010001110000011;
ROM[42567] <= 32'b00000000011100010010000000100011;
ROM[42568] <= 32'b00000000010000010000000100010011;
ROM[42569] <= 32'b00000001010000000000001110010011;
ROM[42570] <= 32'b01000000011100011000001110110011;
ROM[42571] <= 32'b00000000000000111010000010000011;
ROM[42572] <= 32'b11111111110000010000000100010011;
ROM[42573] <= 32'b00000000000000010010001110000011;
ROM[42574] <= 32'b00000000011100100010000000100011;
ROM[42575] <= 32'b00000000010000100000000100010011;
ROM[42576] <= 32'b00000001010000000000001110010011;
ROM[42577] <= 32'b01000000011100011000001110110011;
ROM[42578] <= 32'b00000000010000111010000110000011;
ROM[42579] <= 32'b00000000100000111010001000000011;
ROM[42580] <= 32'b00000000110000111010001010000011;
ROM[42581] <= 32'b00000001000000111010001100000011;
ROM[42582] <= 32'b00000000000000001000000011100111;
ROM[42583] <= 32'b00000000000000010010000000100011;
ROM[42584] <= 32'b00000000010000010000000100010011;
ROM[42585] <= 32'b00000000000000100010001110000011;
ROM[42586] <= 32'b00000000011100010010000000100011;
ROM[42587] <= 32'b00000000010000010000000100010011;
ROM[42588] <= 32'b11111111110000010000000100010011;
ROM[42589] <= 32'b00000000000000010010001110000011;
ROM[42590] <= 32'b00000000000000111000001010010011;
ROM[42591] <= 32'b00000000010000100010001110000011;
ROM[42592] <= 32'b00000000011100010010000000100011;
ROM[42593] <= 32'b00000000010000010000000100010011;
ROM[42594] <= 32'b00000000010000000000001110010011;
ROM[42595] <= 32'b00000000011100010010000000100011;
ROM[42596] <= 32'b00000000010000010000000100010011;
ROM[42597] <= 32'b00000000000000101010001110110111;
ROM[42598] <= 32'b10011110000000111000001110010011;
ROM[42599] <= 32'b00000000111000111000001110110011;
ROM[42600] <= 32'b00000000011100010010000000100011;
ROM[42601] <= 32'b00000000010000010000000100010011;
ROM[42602] <= 32'b00000000001100010010000000100011;
ROM[42603] <= 32'b00000000010000010000000100010011;
ROM[42604] <= 32'b00000000010000010010000000100011;
ROM[42605] <= 32'b00000000010000010000000100010011;
ROM[42606] <= 32'b00000000010100010010000000100011;
ROM[42607] <= 32'b00000000010000010000000100010011;
ROM[42608] <= 32'b00000000011000010010000000100011;
ROM[42609] <= 32'b00000000010000010000000100010011;
ROM[42610] <= 32'b00000001010000000000001110010011;
ROM[42611] <= 32'b00000000100000111000001110010011;
ROM[42612] <= 32'b01000000011100010000001110110011;
ROM[42613] <= 32'b00000000011100000000001000110011;
ROM[42614] <= 32'b00000000001000000000000110110011;
ROM[42615] <= 32'b11100101000111100111000011101111;
ROM[42616] <= 32'b11111111110000010000000100010011;
ROM[42617] <= 32'b00000000000000010010001110000011;
ROM[42618] <= 32'b00000000011100011010000000100011;
ROM[42619] <= 32'b00000000110100101000010000110011;
ROM[42620] <= 32'b00000000100001000010001110000011;
ROM[42621] <= 32'b00000000011100010010000000100011;
ROM[42622] <= 32'b00000000010000010000000100010011;
ROM[42623] <= 32'b00000000000000011010001110000011;
ROM[42624] <= 32'b00000000011100010010000000100011;
ROM[42625] <= 32'b00000000010000010000000100010011;
ROM[42626] <= 32'b11111111110000010000000100010011;
ROM[42627] <= 32'b00000000000000010010001110000011;
ROM[42628] <= 32'b11111111110000010000000100010011;
ROM[42629] <= 32'b00000000000000010010010000000011;
ROM[42630] <= 32'b00000000011101000000001110110011;
ROM[42631] <= 32'b00000000011100010010000000100011;
ROM[42632] <= 32'b00000000010000010000000100010011;
ROM[42633] <= 32'b11111111110000010000000100010011;
ROM[42634] <= 32'b00000000000000010010001110000011;
ROM[42635] <= 32'b00000000000000111000001100010011;
ROM[42636] <= 32'b00000000110100110000010000110011;
ROM[42637] <= 32'b00000000000001000010001110000011;
ROM[42638] <= 32'b00000000011100010010000000100011;
ROM[42639] <= 32'b00000000010000010000000100010011;
ROM[42640] <= 32'b00000001010000000000001110010011;
ROM[42641] <= 32'b01000000011100011000001110110011;
ROM[42642] <= 32'b00000000000000111010000010000011;
ROM[42643] <= 32'b11111111110000010000000100010011;
ROM[42644] <= 32'b00000000000000010010001110000011;
ROM[42645] <= 32'b00000000011100100010000000100011;
ROM[42646] <= 32'b00000000010000100000000100010011;
ROM[42647] <= 32'b00000001010000000000001110010011;
ROM[42648] <= 32'b01000000011100011000001110110011;
ROM[42649] <= 32'b00000000010000111010000110000011;
ROM[42650] <= 32'b00000000100000111010001000000011;
ROM[42651] <= 32'b00000000110000111010001010000011;
ROM[42652] <= 32'b00000001000000111010001100000011;
ROM[42653] <= 32'b00000000000000001000000011100111;
ROM[42654] <= 32'b00000000000000010010000000100011;
ROM[42655] <= 32'b00000000010000010000000100010011;
ROM[42656] <= 32'b00000000000000100010001110000011;
ROM[42657] <= 32'b00000000011100010010000000100011;
ROM[42658] <= 32'b00000000010000010000000100010011;
ROM[42659] <= 32'b11111111110000010000000100010011;
ROM[42660] <= 32'b00000000000000010010001110000011;
ROM[42661] <= 32'b00000000000000111000001010010011;
ROM[42662] <= 32'b00000000010000100010001110000011;
ROM[42663] <= 32'b00000000011100010010000000100011;
ROM[42664] <= 32'b00000000010000010000000100010011;
ROM[42665] <= 32'b00000000010000000000001110010011;
ROM[42666] <= 32'b00000000011100010010000000100011;
ROM[42667] <= 32'b00000000010000010000000100010011;
ROM[42668] <= 32'b00000000000000101010001110110111;
ROM[42669] <= 32'b10101111110000111000001110010011;
ROM[42670] <= 32'b00000000111000111000001110110011;
ROM[42671] <= 32'b00000000011100010010000000100011;
ROM[42672] <= 32'b00000000010000010000000100010011;
ROM[42673] <= 32'b00000000001100010010000000100011;
ROM[42674] <= 32'b00000000010000010000000100010011;
ROM[42675] <= 32'b00000000010000010010000000100011;
ROM[42676] <= 32'b00000000010000010000000100010011;
ROM[42677] <= 32'b00000000010100010010000000100011;
ROM[42678] <= 32'b00000000010000010000000100010011;
ROM[42679] <= 32'b00000000011000010010000000100011;
ROM[42680] <= 32'b00000000010000010000000100010011;
ROM[42681] <= 32'b00000001010000000000001110010011;
ROM[42682] <= 32'b00000000100000111000001110010011;
ROM[42683] <= 32'b01000000011100010000001110110011;
ROM[42684] <= 32'b00000000011100000000001000110011;
ROM[42685] <= 32'b00000000001000000000000110110011;
ROM[42686] <= 32'b11010011010111100111000011101111;
ROM[42687] <= 32'b11111111110000010000000100010011;
ROM[42688] <= 32'b00000000000000010010001110000011;
ROM[42689] <= 32'b00000000011100011010000000100011;
ROM[42690] <= 32'b00000000100000100010001110000011;
ROM[42691] <= 32'b00000000011100010010000000100011;
ROM[42692] <= 32'b00000000010000010000000100010011;
ROM[42693] <= 32'b00000000110100101000010000110011;
ROM[42694] <= 32'b00000000100001000010001110000011;
ROM[42695] <= 32'b00000000011100010010000000100011;
ROM[42696] <= 32'b00000000010000010000000100010011;
ROM[42697] <= 32'b00000000000000011010001110000011;
ROM[42698] <= 32'b00000000011100010010000000100011;
ROM[42699] <= 32'b00000000010000010000000100010011;
ROM[42700] <= 32'b11111111110000010000000100010011;
ROM[42701] <= 32'b00000000000000010010001110000011;
ROM[42702] <= 32'b11111111110000010000000100010011;
ROM[42703] <= 32'b00000000000000010010010000000011;
ROM[42704] <= 32'b00000000011101000000001110110011;
ROM[42705] <= 32'b00000000011100010010000000100011;
ROM[42706] <= 32'b00000000010000010000000100010011;
ROM[42707] <= 32'b11111111110000010000000100010011;
ROM[42708] <= 32'b00000000000000010010001110000011;
ROM[42709] <= 32'b00000000000000111000001100010011;
ROM[42710] <= 32'b11111111110000010000000100010011;
ROM[42711] <= 32'b00000000000000010010001110000011;
ROM[42712] <= 32'b00000000110100110000010000110011;
ROM[42713] <= 32'b00000000011101000010000000100011;
ROM[42714] <= 32'b00000000000000000000001110010011;
ROM[42715] <= 32'b00000000011100010010000000100011;
ROM[42716] <= 32'b00000000010000010000000100010011;
ROM[42717] <= 32'b00000001010000000000001110010011;
ROM[42718] <= 32'b01000000011100011000001110110011;
ROM[42719] <= 32'b00000000000000111010000010000011;
ROM[42720] <= 32'b11111111110000010000000100010011;
ROM[42721] <= 32'b00000000000000010010001110000011;
ROM[42722] <= 32'b00000000011100100010000000100011;
ROM[42723] <= 32'b00000000010000100000000100010011;
ROM[42724] <= 32'b00000001010000000000001110010011;
ROM[42725] <= 32'b01000000011100011000001110110011;
ROM[42726] <= 32'b00000000010000111010000110000011;
ROM[42727] <= 32'b00000000100000111010001000000011;
ROM[42728] <= 32'b00000000110000111010001010000011;
ROM[42729] <= 32'b00000001000000111010001100000011;
ROM[42730] <= 32'b00000000000000001000000011100111;
ROM[42731] <= 32'b00000000000000010010000000100011;
ROM[42732] <= 32'b00000000010000010000000100010011;
ROM[42733] <= 32'b00000000000000100010001110000011;
ROM[42734] <= 32'b00000000011100010010000000100011;
ROM[42735] <= 32'b00000000010000010000000100010011;
ROM[42736] <= 32'b11111111110000010000000100010011;
ROM[42737] <= 32'b00000000000000010010001110000011;
ROM[42738] <= 32'b00000000000000111000001010010011;
ROM[42739] <= 32'b00000000110100101000010000110011;
ROM[42740] <= 32'b00000000010001000010001110000011;
ROM[42741] <= 32'b00000000011100010010000000100011;
ROM[42742] <= 32'b00000000010000010000000100010011;
ROM[42743] <= 32'b00000000010000000000001110010011;
ROM[42744] <= 32'b00000000011100010010000000100011;
ROM[42745] <= 32'b00000000010000010000000100010011;
ROM[42746] <= 32'b00000000000000101010001110110111;
ROM[42747] <= 32'b11000011010000111000001110010011;
ROM[42748] <= 32'b00000000111000111000001110110011;
ROM[42749] <= 32'b00000000011100010010000000100011;
ROM[42750] <= 32'b00000000010000010000000100010011;
ROM[42751] <= 32'b00000000001100010010000000100011;
ROM[42752] <= 32'b00000000010000010000000100010011;
ROM[42753] <= 32'b00000000010000010010000000100011;
ROM[42754] <= 32'b00000000010000010000000100010011;
ROM[42755] <= 32'b00000000010100010010000000100011;
ROM[42756] <= 32'b00000000010000010000000100010011;
ROM[42757] <= 32'b00000000011000010010000000100011;
ROM[42758] <= 32'b00000000010000010000000100010011;
ROM[42759] <= 32'b00000001010000000000001110010011;
ROM[42760] <= 32'b00000000100000111000001110010011;
ROM[42761] <= 32'b01000000011100010000001110110011;
ROM[42762] <= 32'b00000000011100000000001000110011;
ROM[42763] <= 32'b00000000001000000000000110110011;
ROM[42764] <= 32'b10111111110111100111000011101111;
ROM[42765] <= 32'b11111111110000010000000100010011;
ROM[42766] <= 32'b00000000000000010010001110000011;
ROM[42767] <= 32'b00000000011100011010000000100011;
ROM[42768] <= 32'b00000000110100101000010000110011;
ROM[42769] <= 32'b00000000010001000010001110000011;
ROM[42770] <= 32'b00000000011100010010000000100011;
ROM[42771] <= 32'b00000000010000010000000100010011;
ROM[42772] <= 32'b00000000110100101000010000110011;
ROM[42773] <= 32'b00000000000001000010001110000011;
ROM[42774] <= 32'b00000000011100010010000000100011;
ROM[42775] <= 32'b00000000010000010000000100010011;
ROM[42776] <= 32'b11111111110000010000000100010011;
ROM[42777] <= 32'b00000000000000010010001110000011;
ROM[42778] <= 32'b11111111110000010000000100010011;
ROM[42779] <= 32'b00000000000000010010010000000011;
ROM[42780] <= 32'b00000000011101000010001110110011;
ROM[42781] <= 32'b00000000011100010010000000100011;
ROM[42782] <= 32'b00000000010000010000000100010011;
ROM[42783] <= 32'b11111111110000010000000100010011;
ROM[42784] <= 32'b00000000000000010010001110000011;
ROM[42785] <= 32'b00000000000000111000101001100011;
ROM[42786] <= 32'b00000000000000101010001110110111;
ROM[42787] <= 32'b11001001110000111000001110010011;
ROM[42788] <= 32'b00000000111000111000001110110011;
ROM[42789] <= 32'b00000000000000111000000011100111;
ROM[42790] <= 32'b00001010110000000000000011101111;
ROM[42791] <= 32'b00000000010000100010001110000011;
ROM[42792] <= 32'b00000000011100010010000000100011;
ROM[42793] <= 32'b00000000010000010000000100010011;
ROM[42794] <= 32'b00000000110100101000010000110011;
ROM[42795] <= 32'b00000000100001000010001110000011;
ROM[42796] <= 32'b00000000011100010010000000100011;
ROM[42797] <= 32'b00000000010000010000000100010011;
ROM[42798] <= 32'b00000000000000011010001110000011;
ROM[42799] <= 32'b00000000011100010010000000100011;
ROM[42800] <= 32'b00000000010000010000000100010011;
ROM[42801] <= 32'b11111111110000010000000100010011;
ROM[42802] <= 32'b00000000000000010010001110000011;
ROM[42803] <= 32'b11111111110000010000000100010011;
ROM[42804] <= 32'b00000000000000010010010000000011;
ROM[42805] <= 32'b00000000011101000000001110110011;
ROM[42806] <= 32'b00000000011100010010000000100011;
ROM[42807] <= 32'b00000000010000010000000100010011;
ROM[42808] <= 32'b11111111110000010000000100010011;
ROM[42809] <= 32'b00000000000000010010001110000011;
ROM[42810] <= 32'b00000000000000111000001100010011;
ROM[42811] <= 32'b11111111110000010000000100010011;
ROM[42812] <= 32'b00000000000000010010001110000011;
ROM[42813] <= 32'b00000000110100110000010000110011;
ROM[42814] <= 32'b00000000011101000010000000100011;
ROM[42815] <= 32'b00000000110100101000010000110011;
ROM[42816] <= 32'b00000000010001000010001110000011;
ROM[42817] <= 32'b00000000011100010010000000100011;
ROM[42818] <= 32'b00000000010000010000000100010011;
ROM[42819] <= 32'b00000000000100000000001110010011;
ROM[42820] <= 32'b00000000011100010010000000100011;
ROM[42821] <= 32'b00000000010000010000000100010011;
ROM[42822] <= 32'b11111111110000010000000100010011;
ROM[42823] <= 32'b00000000000000010010001110000011;
ROM[42824] <= 32'b11111111110000010000000100010011;
ROM[42825] <= 32'b00000000000000010010010000000011;
ROM[42826] <= 32'b00000000011101000000001110110011;
ROM[42827] <= 32'b00000000011100010010000000100011;
ROM[42828] <= 32'b00000000010000010000000100010011;
ROM[42829] <= 32'b11111111110000010000000100010011;
ROM[42830] <= 32'b00000000000000010010001110000011;
ROM[42831] <= 32'b00000000110100101000010000110011;
ROM[42832] <= 32'b00000000011101000010001000100011;
ROM[42833] <= 32'b00000000110100101000010000110011;
ROM[42834] <= 32'b00000000100001000010001110000011;
ROM[42835] <= 32'b00000000011100010010000000100011;
ROM[42836] <= 32'b00000000010000010000000100010011;
ROM[42837] <= 32'b00000001010000000000001110010011;
ROM[42838] <= 32'b01000000011100011000001110110011;
ROM[42839] <= 32'b00000000000000111010000010000011;
ROM[42840] <= 32'b11111111110000010000000100010011;
ROM[42841] <= 32'b00000000000000010010001110000011;
ROM[42842] <= 32'b00000000011100100010000000100011;
ROM[42843] <= 32'b00000000010000100000000100010011;
ROM[42844] <= 32'b00000001010000000000001110010011;
ROM[42845] <= 32'b01000000011100011000001110110011;
ROM[42846] <= 32'b00000000010000111010000110000011;
ROM[42847] <= 32'b00000000100000111010001000000011;
ROM[42848] <= 32'b00000000110000111010001010000011;
ROM[42849] <= 32'b00000001000000111010001100000011;
ROM[42850] <= 32'b00000000000000001000000011100111;
ROM[42851] <= 32'b00000000000000100010001110000011;
ROM[42852] <= 32'b00000000011100010010000000100011;
ROM[42853] <= 32'b00000000010000010000000100010011;
ROM[42854] <= 32'b11111111110000010000000100010011;
ROM[42855] <= 32'b00000000000000010010001110000011;
ROM[42856] <= 32'b00000000000000111000001010010011;
ROM[42857] <= 32'b00000000110100101000010000110011;
ROM[42858] <= 32'b00000000010001000010001110000011;
ROM[42859] <= 32'b00000000011100010010000000100011;
ROM[42860] <= 32'b00000000010000010000000100010011;
ROM[42861] <= 32'b00000000000000000000001110010011;
ROM[42862] <= 32'b00000000011100010010000000100011;
ROM[42863] <= 32'b00000000010000010000000100010011;
ROM[42864] <= 32'b11111111110000010000000100010011;
ROM[42865] <= 32'b00000000000000010010001110000011;
ROM[42866] <= 32'b11111111110000010000000100010011;
ROM[42867] <= 32'b00000000000000010010010000000011;
ROM[42868] <= 32'b00000000100000111010001110110011;
ROM[42869] <= 32'b00000000011100010010000000100011;
ROM[42870] <= 32'b00000000010000010000000100010011;
ROM[42871] <= 32'b11111111110000010000000100010011;
ROM[42872] <= 32'b00000000000000010010001110000011;
ROM[42873] <= 32'b00000000000000111000101001100011;
ROM[42874] <= 32'b00000000000000101010001110110111;
ROM[42875] <= 32'b11011111110000111000001110010011;
ROM[42876] <= 32'b00000000111000111000001110110011;
ROM[42877] <= 32'b00000000000000111000000011100111;
ROM[42878] <= 32'b00000100110000000000000011101111;
ROM[42879] <= 32'b00000000110100101000010000110011;
ROM[42880] <= 32'b00000000010001000010001110000011;
ROM[42881] <= 32'b00000000011100010010000000100011;
ROM[42882] <= 32'b00000000010000010000000100010011;
ROM[42883] <= 32'b00000000000100000000001110010011;
ROM[42884] <= 32'b00000000011100010010000000100011;
ROM[42885] <= 32'b00000000010000010000000100010011;
ROM[42886] <= 32'b11111111110000010000000100010011;
ROM[42887] <= 32'b00000000000000010010001110000011;
ROM[42888] <= 32'b11111111110000010000000100010011;
ROM[42889] <= 32'b00000000000000010010010000000011;
ROM[42890] <= 32'b01000000011101000000001110110011;
ROM[42891] <= 32'b00000000011100010010000000100011;
ROM[42892] <= 32'b00000000010000010000000100010011;
ROM[42893] <= 32'b11111111110000010000000100010011;
ROM[42894] <= 32'b00000000000000010010001110000011;
ROM[42895] <= 32'b00000000110100101000010000110011;
ROM[42896] <= 32'b00000000011101000010001000100011;
ROM[42897] <= 32'b00000000000000000000001110010011;
ROM[42898] <= 32'b00000000011100010010000000100011;
ROM[42899] <= 32'b00000000010000010000000100010011;
ROM[42900] <= 32'b00000001010000000000001110010011;
ROM[42901] <= 32'b01000000011100011000001110110011;
ROM[42902] <= 32'b00000000000000111010000010000011;
ROM[42903] <= 32'b11111111110000010000000100010011;
ROM[42904] <= 32'b00000000000000010010001110000011;
ROM[42905] <= 32'b00000000011100100010000000100011;
ROM[42906] <= 32'b00000000010000100000000100010011;
ROM[42907] <= 32'b00000001010000000000001110010011;
ROM[42908] <= 32'b01000000011100011000001110110011;
ROM[42909] <= 32'b00000000010000111010000110000011;
ROM[42910] <= 32'b00000000100000111010001000000011;
ROM[42911] <= 32'b00000000110000111010001010000011;
ROM[42912] <= 32'b00000001000000111010001100000011;
ROM[42913] <= 32'b00000000000000001000000011100111;
ROM[42914] <= 32'b00000000000000010010000000100011;
ROM[42915] <= 32'b00000000010000010000000100010011;
ROM[42916] <= 32'b00000000000000010010000000100011;
ROM[42917] <= 32'b00000000010000010000000100010011;
ROM[42918] <= 32'b00000000000000010010000000100011;
ROM[42919] <= 32'b00000000010000010000000100010011;
ROM[42920] <= 32'b00000000000000100010001110000011;
ROM[42921] <= 32'b00000000011100010010000000100011;
ROM[42922] <= 32'b00000000010000010000000100010011;
ROM[42923] <= 32'b11111111110000010000000100010011;
ROM[42924] <= 32'b00000000000000010010001110000011;
ROM[42925] <= 32'b00000000000000111000001010010011;
ROM[42926] <= 32'b00000000000000000000001110010011;
ROM[42927] <= 32'b00000000011100010010000000100011;
ROM[42928] <= 32'b00000000010000010000000100010011;
ROM[42929] <= 32'b11111111110000010000000100010011;
ROM[42930] <= 32'b00000000000000010010001110000011;
ROM[42931] <= 32'b00000000011100011010000000100011;
ROM[42932] <= 32'b00000000110100101000010000110011;
ROM[42933] <= 32'b00000000010001000010001110000011;
ROM[42934] <= 32'b00000000011100010010000000100011;
ROM[42935] <= 32'b00000000010000010000000100010011;
ROM[42936] <= 32'b00000000000000000000001110010011;
ROM[42937] <= 32'b00000000011100010010000000100011;
ROM[42938] <= 32'b00000000010000010000000100010011;
ROM[42939] <= 32'b11111111110000010000000100010011;
ROM[42940] <= 32'b00000000000000010010001110000011;
ROM[42941] <= 32'b11111111110000010000000100010011;
ROM[42942] <= 32'b00000000000000010010010000000011;
ROM[42943] <= 32'b00000000100000111010001110110011;
ROM[42944] <= 32'b00000000011100010010000000100011;
ROM[42945] <= 32'b00000000010000010000000100010011;
ROM[42946] <= 32'b00000000110100101000010000110011;
ROM[42947] <= 32'b00000000100001000010001110000011;
ROM[42948] <= 32'b00000000011100010010000000100011;
ROM[42949] <= 32'b00000000010000010000000100010011;
ROM[42950] <= 32'b00000000000000000000001110010011;
ROM[42951] <= 32'b00000000011100010010000000100011;
ROM[42952] <= 32'b00000000010000010000000100010011;
ROM[42953] <= 32'b11111111110000010000000100010011;
ROM[42954] <= 32'b00000000000000010010001110000011;
ROM[42955] <= 32'b11111111110000010000000100010011;
ROM[42956] <= 32'b00000000000000010010010000000011;
ROM[42957] <= 32'b00000000011101000000001110110011;
ROM[42958] <= 32'b00000000011100010010000000100011;
ROM[42959] <= 32'b00000000010000010000000100010011;
ROM[42960] <= 32'b11111111110000010000000100010011;
ROM[42961] <= 32'b00000000000000010010001110000011;
ROM[42962] <= 32'b00000000000000111000001100010011;
ROM[42963] <= 32'b00000000110100110000010000110011;
ROM[42964] <= 32'b00000000000001000010001110000011;
ROM[42965] <= 32'b00000000011100010010000000100011;
ROM[42966] <= 32'b00000000010000010000000100010011;
ROM[42967] <= 32'b00000010110100000000001110010011;
ROM[42968] <= 32'b00000000011100010010000000100011;
ROM[42969] <= 32'b00000000010000010000000100010011;
ROM[42970] <= 32'b11111111110000010000000100010011;
ROM[42971] <= 32'b00000000000000010010001110000011;
ROM[42972] <= 32'b11111111110000010000000100010011;
ROM[42973] <= 32'b00000000000000010010010000000011;
ROM[42974] <= 32'b00000000011101000010010010110011;
ROM[42975] <= 32'b00000000100000111010010100110011;
ROM[42976] <= 32'b00000000101001001000001110110011;
ROM[42977] <= 32'b00000000000100111000001110010011;
ROM[42978] <= 32'b00000000000100111111001110010011;
ROM[42979] <= 32'b00000000011100010010000000100011;
ROM[42980] <= 32'b00000000010000010000000100010011;
ROM[42981] <= 32'b11111111110000010000000100010011;
ROM[42982] <= 32'b00000000000000010010001110000011;
ROM[42983] <= 32'b11111111110000010000000100010011;
ROM[42984] <= 32'b00000000000000010010010000000011;
ROM[42985] <= 32'b00000000011101000111001110110011;
ROM[42986] <= 32'b00000000011100010010000000100011;
ROM[42987] <= 32'b00000000010000010000000100010011;
ROM[42988] <= 32'b11111111110000010000000100010011;
ROM[42989] <= 32'b00000000000000010010001110000011;
ROM[42990] <= 32'b00000000000000111000101001100011;
ROM[42991] <= 32'b00000000000000101010001110110111;
ROM[42992] <= 32'b00000000000000111000001110010011;
ROM[42993] <= 32'b00000000111000111000001110110011;
ROM[42994] <= 32'b00000000000000111000000011100111;
ROM[42995] <= 32'b00000000000000000000001110010011;
ROM[42996] <= 32'b00000000011100010010000000100011;
ROM[42997] <= 32'b00000000010000010000000100010011;
ROM[42998] <= 32'b11111111110000010000000100010011;
ROM[42999] <= 32'b00000000000000010010001110000011;
ROM[43000] <= 32'b00000000011100011010010000100011;
ROM[43001] <= 32'b00000000000000000000001110010011;
ROM[43002] <= 32'b00000000011100010010000000100011;
ROM[43003] <= 32'b00000000010000010000000100010011;
ROM[43004] <= 32'b11111111110000010000000100010011;
ROM[43005] <= 32'b00000000000000010010001110000011;
ROM[43006] <= 32'b00000000011100011010001000100011;
ROM[43007] <= 32'b00000100100000000000000011101111;
ROM[43008] <= 32'b00000000000100000000001110010011;
ROM[43009] <= 32'b00000000011100010010000000100011;
ROM[43010] <= 32'b00000000010000010000000100010011;
ROM[43011] <= 32'b11111111110000010000000100010011;
ROM[43012] <= 32'b00000000000000010010001110000011;
ROM[43013] <= 32'b01000000011100000000001110110011;
ROM[43014] <= 32'b00000000011100010010000000100011;
ROM[43015] <= 32'b00000000010000010000000100010011;
ROM[43016] <= 32'b11111111110000010000000100010011;
ROM[43017] <= 32'b00000000000000010010001110000011;
ROM[43018] <= 32'b00000000011100011010010000100011;
ROM[43019] <= 32'b00000000000100000000001110010011;
ROM[43020] <= 32'b00000000011100010010000000100011;
ROM[43021] <= 32'b00000000010000010000000100010011;
ROM[43022] <= 32'b11111111110000010000000100010011;
ROM[43023] <= 32'b00000000000000010010001110000011;
ROM[43024] <= 32'b00000000011100011010001000100011;
ROM[43025] <= 32'b00000000010000011010001110000011;
ROM[43026] <= 32'b00000000011100010010000000100011;
ROM[43027] <= 32'b00000000010000010000000100010011;
ROM[43028] <= 32'b00000000110100101000010000110011;
ROM[43029] <= 32'b00000000010001000010001110000011;
ROM[43030] <= 32'b00000000011100010010000000100011;
ROM[43031] <= 32'b00000000010000010000000100010011;
ROM[43032] <= 32'b11111111110000010000000100010011;
ROM[43033] <= 32'b00000000000000010010001110000011;
ROM[43034] <= 32'b11111111110000010000000100010011;
ROM[43035] <= 32'b00000000000000010010010000000011;
ROM[43036] <= 32'b00000000011101000010001110110011;
ROM[43037] <= 32'b00000000011100010010000000100011;
ROM[43038] <= 32'b00000000010000010000000100010011;
ROM[43039] <= 32'b00000000110100101000010000110011;
ROM[43040] <= 32'b00000000100001000010001110000011;
ROM[43041] <= 32'b00000000011100010010000000100011;
ROM[43042] <= 32'b00000000010000010000000100010011;
ROM[43043] <= 32'b00000000010000000000001110010011;
ROM[43044] <= 32'b00000000011100010010000000100011;
ROM[43045] <= 32'b00000000010000010000000100010011;
ROM[43046] <= 32'b00000000010000011010001110000011;
ROM[43047] <= 32'b00000000011100010010000000100011;
ROM[43048] <= 32'b00000000010000010000000100010011;
ROM[43049] <= 32'b00000000000000101010001110110111;
ROM[43050] <= 32'b00001111000000111000001110010011;
ROM[43051] <= 32'b00000000111000111000001110110011;
ROM[43052] <= 32'b00000000011100010010000000100011;
ROM[43053] <= 32'b00000000010000010000000100010011;
ROM[43054] <= 32'b00000000001100010010000000100011;
ROM[43055] <= 32'b00000000010000010000000100010011;
ROM[43056] <= 32'b00000000010000010010000000100011;
ROM[43057] <= 32'b00000000010000010000000100010011;
ROM[43058] <= 32'b00000000010100010010000000100011;
ROM[43059] <= 32'b00000000010000010000000100010011;
ROM[43060] <= 32'b00000000011000010010000000100011;
ROM[43061] <= 32'b00000000010000010000000100010011;
ROM[43062] <= 32'b00000001010000000000001110010011;
ROM[43063] <= 32'b00000000100000111000001110010011;
ROM[43064] <= 32'b01000000011100010000001110110011;
ROM[43065] <= 32'b00000000011100000000001000110011;
ROM[43066] <= 32'b00000000001000000000000110110011;
ROM[43067] <= 32'b11110100000011100111000011101111;
ROM[43068] <= 32'b11111111110000010000000100010011;
ROM[43069] <= 32'b00000000000000010010001110000011;
ROM[43070] <= 32'b11111111110000010000000100010011;
ROM[43071] <= 32'b00000000000000010010010000000011;
ROM[43072] <= 32'b00000000011101000000001110110011;
ROM[43073] <= 32'b00000000011100010010000000100011;
ROM[43074] <= 32'b00000000010000010000000100010011;
ROM[43075] <= 32'b11111111110000010000000100010011;
ROM[43076] <= 32'b00000000000000010010001110000011;
ROM[43077] <= 32'b00000000000000111000001100010011;
ROM[43078] <= 32'b00000000110100110000010000110011;
ROM[43079] <= 32'b00000000000001000010001110000011;
ROM[43080] <= 32'b00000000011100010010000000100011;
ROM[43081] <= 32'b00000000010000010000000100010011;
ROM[43082] <= 32'b00000000000000101010001110110111;
ROM[43083] <= 32'b00010111010000111000001110010011;
ROM[43084] <= 32'b00000000111000111000001110110011;
ROM[43085] <= 32'b00000000011100010010000000100011;
ROM[43086] <= 32'b00000000010000010000000100010011;
ROM[43087] <= 32'b00000000001100010010000000100011;
ROM[43088] <= 32'b00000000010000010000000100010011;
ROM[43089] <= 32'b00000000010000010010000000100011;
ROM[43090] <= 32'b00000000010000010000000100010011;
ROM[43091] <= 32'b00000000010100010010000000100011;
ROM[43092] <= 32'b00000000010000010000000100010011;
ROM[43093] <= 32'b00000000011000010010000000100011;
ROM[43094] <= 32'b00000000010000010000000100010011;
ROM[43095] <= 32'b00000001010000000000001110010011;
ROM[43096] <= 32'b00000000010000111000001110010011;
ROM[43097] <= 32'b01000000011100010000001110110011;
ROM[43098] <= 32'b00000000011100000000001000110011;
ROM[43099] <= 32'b00000000001000000000000110110011;
ROM[43100] <= 32'b00101110010000000000000011101111;
ROM[43101] <= 32'b11111111110000010000000100010011;
ROM[43102] <= 32'b00000000000000010010001110000011;
ROM[43103] <= 32'b11111111110000010000000100010011;
ROM[43104] <= 32'b00000000000000010010010000000011;
ROM[43105] <= 32'b00000000011101000111001110110011;
ROM[43106] <= 32'b00000000011100010010000000100011;
ROM[43107] <= 32'b00000000010000010000000100010011;
ROM[43108] <= 32'b11111111110000010000000100010011;
ROM[43109] <= 32'b00000000000000010010001110000011;
ROM[43110] <= 32'b01000000011100000000001110110011;
ROM[43111] <= 32'b00000000000100111000001110010011;
ROM[43112] <= 32'b00000000011100010010000000100011;
ROM[43113] <= 32'b00000000010000010000000100010011;
ROM[43114] <= 32'b11111111110000010000000100010011;
ROM[43115] <= 32'b00000000000000010010001110000011;
ROM[43116] <= 32'b00000000000000111000101001100011;
ROM[43117] <= 32'b00000000000000101010001110110111;
ROM[43118] <= 32'b00111000110000111000001110010011;
ROM[43119] <= 32'b00000000111000111000001110110011;
ROM[43120] <= 32'b00000000000000111000000011100111;
ROM[43121] <= 32'b00000000000000011010001110000011;
ROM[43122] <= 32'b00000000011100010010000000100011;
ROM[43123] <= 32'b00000000010000010000000100010011;
ROM[43124] <= 32'b00000000101000000000001110010011;
ROM[43125] <= 32'b00000000011100010010000000100011;
ROM[43126] <= 32'b00000000010000010000000100010011;
ROM[43127] <= 32'b00000000000000101010001110110111;
ROM[43128] <= 32'b00100010100000111000001110010011;
ROM[43129] <= 32'b00000000111000111000001110110011;
ROM[43130] <= 32'b00000000011100010010000000100011;
ROM[43131] <= 32'b00000000010000010000000100010011;
ROM[43132] <= 32'b00000000001100010010000000100011;
ROM[43133] <= 32'b00000000010000010000000100010011;
ROM[43134] <= 32'b00000000010000010010000000100011;
ROM[43135] <= 32'b00000000010000010000000100010011;
ROM[43136] <= 32'b00000000010100010010000000100011;
ROM[43137] <= 32'b00000000010000010000000100010011;
ROM[43138] <= 32'b00000000011000010010000000100011;
ROM[43139] <= 32'b00000000010000010000000100010011;
ROM[43140] <= 32'b00000001010000000000001110010011;
ROM[43141] <= 32'b00000000100000111000001110010011;
ROM[43142] <= 32'b01000000011100010000001110110011;
ROM[43143] <= 32'b00000000011100000000001000110011;
ROM[43144] <= 32'b00000000001000000000000110110011;
ROM[43145] <= 32'b11100000100011100111000011101111;
ROM[43146] <= 32'b00000000110100101000010000110011;
ROM[43147] <= 32'b00000000100001000010001110000011;
ROM[43148] <= 32'b00000000011100010010000000100011;
ROM[43149] <= 32'b00000000010000010000000100010011;
ROM[43150] <= 32'b00000000010000000000001110010011;
ROM[43151] <= 32'b00000000011100010010000000100011;
ROM[43152] <= 32'b00000000010000010000000100010011;
ROM[43153] <= 32'b00000000010000011010001110000011;
ROM[43154] <= 32'b00000000011100010010000000100011;
ROM[43155] <= 32'b00000000010000010000000100010011;
ROM[43156] <= 32'b00000000000000101010001110110111;
ROM[43157] <= 32'b00101001110000111000001110010011;
ROM[43158] <= 32'b00000000111000111000001110110011;
ROM[43159] <= 32'b00000000011100010010000000100011;
ROM[43160] <= 32'b00000000010000010000000100010011;
ROM[43161] <= 32'b00000000001100010010000000100011;
ROM[43162] <= 32'b00000000010000010000000100010011;
ROM[43163] <= 32'b00000000010000010010000000100011;
ROM[43164] <= 32'b00000000010000010000000100010011;
ROM[43165] <= 32'b00000000010100010010000000100011;
ROM[43166] <= 32'b00000000010000010000000100010011;
ROM[43167] <= 32'b00000000011000010010000000100011;
ROM[43168] <= 32'b00000000010000010000000100010011;
ROM[43169] <= 32'b00000001010000000000001110010011;
ROM[43170] <= 32'b00000000100000111000001110010011;
ROM[43171] <= 32'b01000000011100010000001110110011;
ROM[43172] <= 32'b00000000011100000000001000110011;
ROM[43173] <= 32'b00000000001000000000000110110011;
ROM[43174] <= 32'b11011001010011100111000011101111;
ROM[43175] <= 32'b11111111110000010000000100010011;
ROM[43176] <= 32'b00000000000000010010001110000011;
ROM[43177] <= 32'b11111111110000010000000100010011;
ROM[43178] <= 32'b00000000000000010010010000000011;
ROM[43179] <= 32'b00000000011101000000001110110011;
ROM[43180] <= 32'b00000000011100010010000000100011;
ROM[43181] <= 32'b00000000010000010000000100010011;
ROM[43182] <= 32'b11111111110000010000000100010011;
ROM[43183] <= 32'b00000000000000010010001110000011;
ROM[43184] <= 32'b00000000000000111000001100010011;
ROM[43185] <= 32'b00000000110100110000010000110011;
ROM[43186] <= 32'b00000000000001000010001110000011;
ROM[43187] <= 32'b00000000011100010010000000100011;
ROM[43188] <= 32'b00000000010000010000000100010011;
ROM[43189] <= 32'b00000000000000101010001110110111;
ROM[43190] <= 32'b00110010000000111000001110010011;
ROM[43191] <= 32'b00000000111000111000001110110011;
ROM[43192] <= 32'b00000000011100010010000000100011;
ROM[43193] <= 32'b00000000010000010000000100010011;
ROM[43194] <= 32'b00000000001100010010000000100011;
ROM[43195] <= 32'b00000000010000010000000100010011;
ROM[43196] <= 32'b00000000010000010010000000100011;
ROM[43197] <= 32'b00000000010000010000000100010011;
ROM[43198] <= 32'b00000000010100010010000000100011;
ROM[43199] <= 32'b00000000010000010000000100010011;
ROM[43200] <= 32'b00000000011000010010000000100011;
ROM[43201] <= 32'b00000000010000010000000100010011;
ROM[43202] <= 32'b00000001010000000000001110010011;
ROM[43203] <= 32'b00000000010000111000001110010011;
ROM[43204] <= 32'b01000000011100010000001110110011;
ROM[43205] <= 32'b00000000011100000000001000110011;
ROM[43206] <= 32'b00000000001000000000000110110011;
ROM[43207] <= 32'b00100010010000000000000011101111;
ROM[43208] <= 32'b11111111110000010000000100010011;
ROM[43209] <= 32'b00000000000000010010001110000011;
ROM[43210] <= 32'b11111111110000010000000100010011;
ROM[43211] <= 32'b00000000000000010010010000000011;
ROM[43212] <= 32'b00000000011101000000001110110011;
ROM[43213] <= 32'b00000000011100010010000000100011;
ROM[43214] <= 32'b00000000010000010000000100010011;
ROM[43215] <= 32'b11111111110000010000000100010011;
ROM[43216] <= 32'b00000000000000010010001110000011;
ROM[43217] <= 32'b00000000011100011010000000100011;
ROM[43218] <= 32'b00000000010000011010001110000011;
ROM[43219] <= 32'b00000000011100010010000000100011;
ROM[43220] <= 32'b00000000010000010000000100010011;
ROM[43221] <= 32'b00000000000100000000001110010011;
ROM[43222] <= 32'b00000000011100010010000000100011;
ROM[43223] <= 32'b00000000010000010000000100010011;
ROM[43224] <= 32'b11111111110000010000000100010011;
ROM[43225] <= 32'b00000000000000010010001110000011;
ROM[43226] <= 32'b11111111110000010000000100010011;
ROM[43227] <= 32'b00000000000000010010010000000011;
ROM[43228] <= 32'b00000000011101000000001110110011;
ROM[43229] <= 32'b00000000011100010010000000100011;
ROM[43230] <= 32'b00000000010000010000000100010011;
ROM[43231] <= 32'b11111111110000010000000100010011;
ROM[43232] <= 32'b00000000000000010010001110000011;
ROM[43233] <= 32'b00000000011100011010001000100011;
ROM[43234] <= 32'b11001011110111111111000011101111;
ROM[43235] <= 32'b00000000100000011010001110000011;
ROM[43236] <= 32'b00000000011100010010000000100011;
ROM[43237] <= 32'b00000000010000010000000100010011;
ROM[43238] <= 32'b11111111110000010000000100010011;
ROM[43239] <= 32'b00000000000000010010001110000011;
ROM[43240] <= 32'b00000000000000111000101001100011;
ROM[43241] <= 32'b00000000000000101010001110110111;
ROM[43242] <= 32'b00111111110000111000001110010011;
ROM[43243] <= 32'b00000000111000111000001110110011;
ROM[43244] <= 32'b00000000000000111000000011100111;
ROM[43245] <= 32'b00000000000000011010001110000011;
ROM[43246] <= 32'b00000000011100010010000000100011;
ROM[43247] <= 32'b00000000010000010000000100010011;
ROM[43248] <= 32'b00000001010000000000001110010011;
ROM[43249] <= 32'b01000000011100011000001110110011;
ROM[43250] <= 32'b00000000000000111010000010000011;
ROM[43251] <= 32'b11111111110000010000000100010011;
ROM[43252] <= 32'b00000000000000010010001110000011;
ROM[43253] <= 32'b00000000011100100010000000100011;
ROM[43254] <= 32'b00000000010000100000000100010011;
ROM[43255] <= 32'b00000001010000000000001110010011;
ROM[43256] <= 32'b01000000011100011000001110110011;
ROM[43257] <= 32'b00000000010000111010000110000011;
ROM[43258] <= 32'b00000000100000111010001000000011;
ROM[43259] <= 32'b00000000110000111010001010000011;
ROM[43260] <= 32'b00000001000000111010001100000011;
ROM[43261] <= 32'b00000000000000001000000011100111;
ROM[43262] <= 32'b00000101110000000000000011101111;
ROM[43263] <= 32'b00000000000000011010001110000011;
ROM[43264] <= 32'b00000000011100010010000000100011;
ROM[43265] <= 32'b00000000010000010000000100010011;
ROM[43266] <= 32'b11111111110000010000000100010011;
ROM[43267] <= 32'b00000000000000010010001110000011;
ROM[43268] <= 32'b01000000011100000000001110110011;
ROM[43269] <= 32'b00000000011100010010000000100011;
ROM[43270] <= 32'b00000000010000010000000100010011;
ROM[43271] <= 32'b00000001010000000000001110010011;
ROM[43272] <= 32'b01000000011100011000001110110011;
ROM[43273] <= 32'b00000000000000111010000010000011;
ROM[43274] <= 32'b11111111110000010000000100010011;
ROM[43275] <= 32'b00000000000000010010001110000011;
ROM[43276] <= 32'b00000000011100100010000000100011;
ROM[43277] <= 32'b00000000010000100000000100010011;
ROM[43278] <= 32'b00000001010000000000001110010011;
ROM[43279] <= 32'b01000000011100011000001110110011;
ROM[43280] <= 32'b00000000010000111010000110000011;
ROM[43281] <= 32'b00000000100000111010001000000011;
ROM[43282] <= 32'b00000000110000111010001010000011;
ROM[43283] <= 32'b00000001000000111010001100000011;
ROM[43284] <= 32'b00000000000000001000000011100111;
ROM[43285] <= 32'b00000000000000100010001110000011;
ROM[43286] <= 32'b00000000011100010010000000100011;
ROM[43287] <= 32'b00000000010000010000000100010011;
ROM[43288] <= 32'b00000011000000000000001110010011;
ROM[43289] <= 32'b00000000011100010010000000100011;
ROM[43290] <= 32'b00000000010000010000000100010011;
ROM[43291] <= 32'b11111111110000010000000100010011;
ROM[43292] <= 32'b00000000000000010010001110000011;
ROM[43293] <= 32'b11111111110000010000000100010011;
ROM[43294] <= 32'b00000000000000010010010000000011;
ROM[43295] <= 32'b00000000011101000010001110110011;
ROM[43296] <= 32'b00000000011100010010000000100011;
ROM[43297] <= 32'b00000000010000010000000100010011;
ROM[43298] <= 32'b11111111110000010000000100010011;
ROM[43299] <= 32'b00000000000000010010001110000011;
ROM[43300] <= 32'b01000000011100000000001110110011;
ROM[43301] <= 32'b00000000000100111000001110010011;
ROM[43302] <= 32'b00000000011100010010000000100011;
ROM[43303] <= 32'b00000000010000010000000100010011;
ROM[43304] <= 32'b00000000000000100010001110000011;
ROM[43305] <= 32'b00000000011100010010000000100011;
ROM[43306] <= 32'b00000000010000010000000100010011;
ROM[43307] <= 32'b00000011100100000000001110010011;
ROM[43308] <= 32'b00000000011100010010000000100011;
ROM[43309] <= 32'b00000000010000010000000100010011;
ROM[43310] <= 32'b11111111110000010000000100010011;
ROM[43311] <= 32'b00000000000000010010001110000011;
ROM[43312] <= 32'b11111111110000010000000100010011;
ROM[43313] <= 32'b00000000000000010010010000000011;
ROM[43314] <= 32'b00000000100000111010001110110011;
ROM[43315] <= 32'b00000000011100010010000000100011;
ROM[43316] <= 32'b00000000010000010000000100010011;
ROM[43317] <= 32'b11111111110000010000000100010011;
ROM[43318] <= 32'b00000000000000010010001110000011;
ROM[43319] <= 32'b01000000011100000000001110110011;
ROM[43320] <= 32'b00000000000100111000001110010011;
ROM[43321] <= 32'b00000000011100010010000000100011;
ROM[43322] <= 32'b00000000010000010000000100010011;
ROM[43323] <= 32'b11111111110000010000000100010011;
ROM[43324] <= 32'b00000000000000010010001110000011;
ROM[43325] <= 32'b11111111110000010000000100010011;
ROM[43326] <= 32'b00000000000000010010010000000011;
ROM[43327] <= 32'b00000000011101000111001110110011;
ROM[43328] <= 32'b00000000011100010010000000100011;
ROM[43329] <= 32'b00000000010000010000000100010011;
ROM[43330] <= 32'b00000001010000000000001110010011;
ROM[43331] <= 32'b01000000011100011000001110110011;
ROM[43332] <= 32'b00000000000000111010000010000011;
ROM[43333] <= 32'b11111111110000010000000100010011;
ROM[43334] <= 32'b00000000000000010010001110000011;
ROM[43335] <= 32'b00000000011100100010000000100011;
ROM[43336] <= 32'b00000000010000100000000100010011;
ROM[43337] <= 32'b00000001010000000000001110010011;
ROM[43338] <= 32'b01000000011100011000001110110011;
ROM[43339] <= 32'b00000000010000111010000110000011;
ROM[43340] <= 32'b00000000100000111010001000000011;
ROM[43341] <= 32'b00000000110000111010001010000011;
ROM[43342] <= 32'b00000001000000111010001100000011;
ROM[43343] <= 32'b00000000000000001000000011100111;
ROM[43344] <= 32'b00000000000000100010001110000011;
ROM[43345] <= 32'b00000000011100010010000000100011;
ROM[43346] <= 32'b00000000010000010000000100010011;
ROM[43347] <= 32'b00000011000000000000001110010011;
ROM[43348] <= 32'b00000000011100010010000000100011;
ROM[43349] <= 32'b00000000010000010000000100010011;
ROM[43350] <= 32'b11111111110000010000000100010011;
ROM[43351] <= 32'b00000000000000010010001110000011;
ROM[43352] <= 32'b11111111110000010000000100010011;
ROM[43353] <= 32'b00000000000000010010010000000011;
ROM[43354] <= 32'b01000000011101000000001110110011;
ROM[43355] <= 32'b00000000011100010010000000100011;
ROM[43356] <= 32'b00000000010000010000000100010011;
ROM[43357] <= 32'b00000001010000000000001110010011;
ROM[43358] <= 32'b01000000011100011000001110110011;
ROM[43359] <= 32'b00000000000000111010000010000011;
ROM[43360] <= 32'b11111111110000010000000100010011;
ROM[43361] <= 32'b00000000000000010010001110000011;
ROM[43362] <= 32'b00000000011100100010000000100011;
ROM[43363] <= 32'b00000000010000100000000100010011;
ROM[43364] <= 32'b00000001010000000000001110010011;
ROM[43365] <= 32'b01000000011100011000001110110011;
ROM[43366] <= 32'b00000000010000111010000110000011;
ROM[43367] <= 32'b00000000100000111010001000000011;
ROM[43368] <= 32'b00000000110000111010001010000011;
ROM[43369] <= 32'b00000001000000111010001100000011;
ROM[43370] <= 32'b00000000000000001000000011100111;
ROM[43371] <= 32'b00000000000000100010001110000011;
ROM[43372] <= 32'b00000000011100010010000000100011;
ROM[43373] <= 32'b00000000010000010000000100010011;
ROM[43374] <= 32'b00000011000000000000001110010011;
ROM[43375] <= 32'b00000000011100010010000000100011;
ROM[43376] <= 32'b00000000010000010000000100010011;
ROM[43377] <= 32'b11111111110000010000000100010011;
ROM[43378] <= 32'b00000000000000010010001110000011;
ROM[43379] <= 32'b11111111110000010000000100010011;
ROM[43380] <= 32'b00000000000000010010010000000011;
ROM[43381] <= 32'b00000000011101000000001110110011;
ROM[43382] <= 32'b00000000011100010010000000100011;
ROM[43383] <= 32'b00000000010000010000000100010011;
ROM[43384] <= 32'b00000001010000000000001110010011;
ROM[43385] <= 32'b01000000011100011000001110110011;
ROM[43386] <= 32'b00000000000000111010000010000011;
ROM[43387] <= 32'b11111111110000010000000100010011;
ROM[43388] <= 32'b00000000000000010010001110000011;
ROM[43389] <= 32'b00000000011100100010000000100011;
ROM[43390] <= 32'b00000000010000100000000100010011;
ROM[43391] <= 32'b00000001010000000000001110010011;
ROM[43392] <= 32'b01000000011100011000001110110011;
ROM[43393] <= 32'b00000000010000111010000110000011;
ROM[43394] <= 32'b00000000100000111010001000000011;
ROM[43395] <= 32'b00000000110000111010001010000011;
ROM[43396] <= 32'b00000001000000111010001100000011;
ROM[43397] <= 32'b00000000000000001000000011100111;
ROM[43398] <= 32'b00000000000000100010001110000011;
ROM[43399] <= 32'b00000000011100010010000000100011;
ROM[43400] <= 32'b00000000010000010000000100010011;
ROM[43401] <= 32'b11111111110000010000000100010011;
ROM[43402] <= 32'b00000000000000010010001110000011;
ROM[43403] <= 32'b00000000000000111000001010010011;
ROM[43404] <= 32'b00000000000000000000001110010011;
ROM[43405] <= 32'b00000000011100010010000000100011;
ROM[43406] <= 32'b00000000010000010000000100010011;
ROM[43407] <= 32'b11111111110000010000000100010011;
ROM[43408] <= 32'b00000000000000010010001110000011;
ROM[43409] <= 32'b00000000110100101000010000110011;
ROM[43410] <= 32'b00000000011101000010001000100011;
ROM[43411] <= 32'b00000000000000000000001110010011;
ROM[43412] <= 32'b00000000011100010010000000100011;
ROM[43413] <= 32'b00000000010000010000000100010011;
ROM[43414] <= 32'b00000001010000000000001110010011;
ROM[43415] <= 32'b01000000011100011000001110110011;
ROM[43416] <= 32'b00000000000000111010000010000011;
ROM[43417] <= 32'b11111111110000010000000100010011;
ROM[43418] <= 32'b00000000000000010010001110000011;
ROM[43419] <= 32'b00000000011100100010000000100011;
ROM[43420] <= 32'b00000000010000100000000100010011;
ROM[43421] <= 32'b00000001010000000000001110010011;
ROM[43422] <= 32'b01000000011100011000001110110011;
ROM[43423] <= 32'b00000000010000111010000110000011;
ROM[43424] <= 32'b00000000100000111010001000000011;
ROM[43425] <= 32'b00000000110000111010001010000011;
ROM[43426] <= 32'b00000001000000111010001100000011;
ROM[43427] <= 32'b00000000000000001000000011100111;
ROM[43428] <= 32'b00000000000000100010001110000011;
ROM[43429] <= 32'b00000000011100010010000000100011;
ROM[43430] <= 32'b00000000010000010000000100010011;
ROM[43431] <= 32'b11111111110000010000000100010011;
ROM[43432] <= 32'b00000000000000010010001110000011;
ROM[43433] <= 32'b00000000000000111000001010010011;
ROM[43434] <= 32'b00000000010100010010000000100011;
ROM[43435] <= 32'b00000000010000010000000100010011;
ROM[43436] <= 32'b00000000000000101010001110110111;
ROM[43437] <= 32'b01101111110000111000001110010011;
ROM[43438] <= 32'b00000000111000111000001110110011;
ROM[43439] <= 32'b00000000011100010010000000100011;
ROM[43440] <= 32'b00000000010000010000000100010011;
ROM[43441] <= 32'b00000000001100010010000000100011;
ROM[43442] <= 32'b00000000010000010000000100010011;
ROM[43443] <= 32'b00000000010000010010000000100011;
ROM[43444] <= 32'b00000000010000010000000100010011;
ROM[43445] <= 32'b00000000010100010010000000100011;
ROM[43446] <= 32'b00000000010000010000000100010011;
ROM[43447] <= 32'b00000000011000010010000000100011;
ROM[43448] <= 32'b00000000010000010000000100010011;
ROM[43449] <= 32'b00000001010000000000001110010011;
ROM[43450] <= 32'b00000000010000111000001110010011;
ROM[43451] <= 32'b01000000011100010000001110110011;
ROM[43452] <= 32'b00000000011100000000001000110011;
ROM[43453] <= 32'b00000000001000000000000110110011;
ROM[43454] <= 32'b11110010000111111111000011101111;
ROM[43455] <= 32'b11111111110000010000000100010011;
ROM[43456] <= 32'b00000000000000010010001110000011;
ROM[43457] <= 32'b00000000011101100010000000100011;
ROM[43458] <= 32'b00000000000000000000001110010011;
ROM[43459] <= 32'b00000000011100010010000000100011;
ROM[43460] <= 32'b00000000010000010000000100010011;
ROM[43461] <= 32'b11111111110000010000000100010011;
ROM[43462] <= 32'b00000000000000010010001110000011;
ROM[43463] <= 32'b00000000110100101000010000110011;
ROM[43464] <= 32'b00000000011101000010001000100011;
ROM[43465] <= 32'b00000000010000100010001110000011;
ROM[43466] <= 32'b00000000011100010010000000100011;
ROM[43467] <= 32'b00000000010000010000000100010011;
ROM[43468] <= 32'b00000000000000000000001110010011;
ROM[43469] <= 32'b00000000011100010010000000100011;
ROM[43470] <= 32'b00000000010000010000000100010011;
ROM[43471] <= 32'b11111111110000010000000100010011;
ROM[43472] <= 32'b00000000000000010010001110000011;
ROM[43473] <= 32'b11111111110000010000000100010011;
ROM[43474] <= 32'b00000000000000010010010000000011;
ROM[43475] <= 32'b00000000011101000010001110110011;
ROM[43476] <= 32'b00000000011100010010000000100011;
ROM[43477] <= 32'b00000000010000010000000100010011;
ROM[43478] <= 32'b11111111110000010000000100010011;
ROM[43479] <= 32'b00000000000000010010001110000011;
ROM[43480] <= 32'b00000000000000111000101001100011;
ROM[43481] <= 32'b00000000000000101010001110110111;
ROM[43482] <= 32'b01110111100000111000001110010011;
ROM[43483] <= 32'b00000000111000111000001110110011;
ROM[43484] <= 32'b00000000000000111000000011100111;
ROM[43485] <= 32'b00001001110000000000000011101111;
ROM[43486] <= 32'b00000000010000100010001110000011;
ROM[43487] <= 32'b00000000011100010010000000100011;
ROM[43488] <= 32'b00000000010000010000000100010011;
ROM[43489] <= 32'b11111111110000010000000100010011;
ROM[43490] <= 32'b00000000000000010010001110000011;
ROM[43491] <= 32'b01000000011100000000001110110011;
ROM[43492] <= 32'b00000000011100010010000000100011;
ROM[43493] <= 32'b00000000010000010000000100010011;
ROM[43494] <= 32'b11111111110000010000000100010011;
ROM[43495] <= 32'b00000000000000010010001110000011;
ROM[43496] <= 32'b00000000011100100010001000100011;
ROM[43497] <= 32'b00000000010100010010000000100011;
ROM[43498] <= 32'b00000000010000010000000100010011;
ROM[43499] <= 32'b00000010110100000000001110010011;
ROM[43500] <= 32'b00000000011100010010000000100011;
ROM[43501] <= 32'b00000000010000010000000100010011;
ROM[43502] <= 32'b00000000000000101011001110110111;
ROM[43503] <= 32'b10000000010000111000001110010011;
ROM[43504] <= 32'b00000000111000111000001110110011;
ROM[43505] <= 32'b00000000011100010010000000100011;
ROM[43506] <= 32'b00000000010000010000000100010011;
ROM[43507] <= 32'b00000000001100010010000000100011;
ROM[43508] <= 32'b00000000010000010000000100010011;
ROM[43509] <= 32'b00000000010000010010000000100011;
ROM[43510] <= 32'b00000000010000010000000100010011;
ROM[43511] <= 32'b00000000010100010010000000100011;
ROM[43512] <= 32'b00000000010000010000000100010011;
ROM[43513] <= 32'b00000000011000010010000000100011;
ROM[43514] <= 32'b00000000010000010000000100010011;
ROM[43515] <= 32'b00000001010000000000001110010011;
ROM[43516] <= 32'b00000000100000111000001110010011;
ROM[43517] <= 32'b01000000011100010000001110110011;
ROM[43518] <= 32'b00000000011100000000001000110011;
ROM[43519] <= 32'b00000000001000000000000110110011;
ROM[43520] <= 32'b10111010110011111111000011101111;
ROM[43521] <= 32'b11111111110000010000000100010011;
ROM[43522] <= 32'b00000000000000010010001110000011;
ROM[43523] <= 32'b00000000011101100010000000100011;
ROM[43524] <= 32'b00000000010100010010000000100011;
ROM[43525] <= 32'b00000000010000010000000100010011;
ROM[43526] <= 32'b00000000010000100010001110000011;
ROM[43527] <= 32'b00000000011100010010000000100011;
ROM[43528] <= 32'b00000000010000010000000100010011;
ROM[43529] <= 32'b00000000000000101011001110110111;
ROM[43530] <= 32'b10000111000000111000001110010011;
ROM[43531] <= 32'b00000000111000111000001110110011;
ROM[43532] <= 32'b00000000011100010010000000100011;
ROM[43533] <= 32'b00000000010000010000000100010011;
ROM[43534] <= 32'b00000000001100010010000000100011;
ROM[43535] <= 32'b00000000010000010000000100010011;
ROM[43536] <= 32'b00000000010000010010000000100011;
ROM[43537] <= 32'b00000000010000010000000100010011;
ROM[43538] <= 32'b00000000010100010010000000100011;
ROM[43539] <= 32'b00000000010000010000000100010011;
ROM[43540] <= 32'b00000000011000010010000000100011;
ROM[43541] <= 32'b00000000010000010000000100010011;
ROM[43542] <= 32'b00000001010000000000001110010011;
ROM[43543] <= 32'b00000000100000111000001110010011;
ROM[43544] <= 32'b01000000011100010000001110110011;
ROM[43545] <= 32'b00000000011100000000001000110011;
ROM[43546] <= 32'b00000000001000000000000110110011;
ROM[43547] <= 32'b00000101010000000000000011101111;
ROM[43548] <= 32'b11111111110000010000000100010011;
ROM[43549] <= 32'b00000000000000010010001110000011;
ROM[43550] <= 32'b00000000011101100010000000100011;
ROM[43551] <= 32'b00000000000000000000001110010011;
ROM[43552] <= 32'b00000000011100010010000000100011;
ROM[43553] <= 32'b00000000010000010000000100010011;
ROM[43554] <= 32'b00000001010000000000001110010011;
ROM[43555] <= 32'b01000000011100011000001110110011;
ROM[43556] <= 32'b00000000000000111010000010000011;
ROM[43557] <= 32'b11111111110000010000000100010011;
ROM[43558] <= 32'b00000000000000010010001110000011;
ROM[43559] <= 32'b00000000011100100010000000100011;
ROM[43560] <= 32'b00000000010000100000000100010011;
ROM[43561] <= 32'b00000001010000000000001110010011;
ROM[43562] <= 32'b01000000011100011000001110110011;
ROM[43563] <= 32'b00000000010000111010000110000011;
ROM[43564] <= 32'b00000000100000111010001000000011;
ROM[43565] <= 32'b00000000110000111010001010000011;
ROM[43566] <= 32'b00000001000000111010001100000011;
ROM[43567] <= 32'b00000000000000001000000011100111;
ROM[43568] <= 32'b00000000000000010010000000100011;
ROM[43569] <= 32'b00000000010000010000000100010011;
ROM[43570] <= 32'b00000000000000100010001110000011;
ROM[43571] <= 32'b00000000011100010010000000100011;
ROM[43572] <= 32'b00000000010000010000000100010011;
ROM[43573] <= 32'b11111111110000010000000100010011;
ROM[43574] <= 32'b00000000000000010010001110000011;
ROM[43575] <= 32'b00000000000000111000001010010011;
ROM[43576] <= 32'b00000000010000100010001110000011;
ROM[43577] <= 32'b00000000011100010010000000100011;
ROM[43578] <= 32'b00000000010000010000000100010011;
ROM[43579] <= 32'b00000000101000000000001110010011;
ROM[43580] <= 32'b00000000011100010010000000100011;
ROM[43581] <= 32'b00000000010000010000000100010011;
ROM[43582] <= 32'b11111111110000010000000100010011;
ROM[43583] <= 32'b00000000000000010010001110000011;
ROM[43584] <= 32'b11111111110000010000000100010011;
ROM[43585] <= 32'b00000000000000010010010000000011;
ROM[43586] <= 32'b00000000011101000010001110110011;
ROM[43587] <= 32'b00000000011100010010000000100011;
ROM[43588] <= 32'b00000000010000010000000100010011;
ROM[43589] <= 32'b11111111110000010000000100010011;
ROM[43590] <= 32'b00000000000000010010001110000011;
ROM[43591] <= 32'b00000000000000111000101001100011;
ROM[43592] <= 32'b00000000000000101011001110110111;
ROM[43593] <= 32'b10110100100000111000001110010011;
ROM[43594] <= 32'b00000000111000111000001110110011;
ROM[43595] <= 32'b00000000000000111000000011100111;
ROM[43596] <= 32'b00000000010000100010001110000011;
ROM[43597] <= 32'b00000000011100010010000000100011;
ROM[43598] <= 32'b00000000010000010000000100010011;
ROM[43599] <= 32'b00000000101000000000001110010011;
ROM[43600] <= 32'b00000000011100010010000000100011;
ROM[43601] <= 32'b00000000010000010000000100010011;
ROM[43602] <= 32'b00000000000000101011001110110111;
ROM[43603] <= 32'b10011001010000111000001110010011;
ROM[43604] <= 32'b00000000111000111000001110110011;
ROM[43605] <= 32'b00000000011100010010000000100011;
ROM[43606] <= 32'b00000000010000010000000100010011;
ROM[43607] <= 32'b00000000001100010010000000100011;
ROM[43608] <= 32'b00000000010000010000000100010011;
ROM[43609] <= 32'b00000000010000010010000000100011;
ROM[43610] <= 32'b00000000010000010000000100010011;
ROM[43611] <= 32'b00000000010100010010000000100011;
ROM[43612] <= 32'b00000000010000010000000100010011;
ROM[43613] <= 32'b00000000011000010010000000100011;
ROM[43614] <= 32'b00000000010000010000000100010011;
ROM[43615] <= 32'b00000001010000000000001110010011;
ROM[43616] <= 32'b00000000100000111000001110010011;
ROM[43617] <= 32'b01000000011100010000001110110011;
ROM[43618] <= 32'b00000000011100000000001000110011;
ROM[43619] <= 32'b00000000001000000000000110110011;
ROM[43620] <= 32'b10100001100011100111000011101111;
ROM[43621] <= 32'b11111111110000010000000100010011;
ROM[43622] <= 32'b00000000000000010010001110000011;
ROM[43623] <= 32'b00000000011100011010000000100011;
ROM[43624] <= 32'b00000000010100010010000000100011;
ROM[43625] <= 32'b00000000010000010000000100010011;
ROM[43626] <= 32'b00000000000000011010001110000011;
ROM[43627] <= 32'b00000000011100010010000000100011;
ROM[43628] <= 32'b00000000010000010000000100010011;
ROM[43629] <= 32'b00000000000000101011001110110111;
ROM[43630] <= 32'b10100000000000111000001110010011;
ROM[43631] <= 32'b00000000111000111000001110110011;
ROM[43632] <= 32'b00000000011100010010000000100011;
ROM[43633] <= 32'b00000000010000010000000100010011;
ROM[43634] <= 32'b00000000001100010010000000100011;
ROM[43635] <= 32'b00000000010000010000000100010011;
ROM[43636] <= 32'b00000000010000010010000000100011;
ROM[43637] <= 32'b00000000010000010000000100010011;
ROM[43638] <= 32'b00000000010100010010000000100011;
ROM[43639] <= 32'b00000000010000010000000100010011;
ROM[43640] <= 32'b00000000011000010010000000100011;
ROM[43641] <= 32'b00000000010000010000000100010011;
ROM[43642] <= 32'b00000001010000000000001110010011;
ROM[43643] <= 32'b00000000100000111000001110010011;
ROM[43644] <= 32'b01000000011100010000001110110011;
ROM[43645] <= 32'b00000000011100000000001000110011;
ROM[43646] <= 32'b00000000001000000000000110110011;
ROM[43647] <= 32'b11101100010111111111000011101111;
ROM[43648] <= 32'b11111111110000010000000100010011;
ROM[43649] <= 32'b00000000000000010010001110000011;
ROM[43650] <= 32'b00000000011101100010000000100011;
ROM[43651] <= 32'b00000000010100010010000000100011;
ROM[43652] <= 32'b00000000010000010000000100010011;
ROM[43653] <= 32'b00000000010000100010001110000011;
ROM[43654] <= 32'b00000000011100010010000000100011;
ROM[43655] <= 32'b00000000010000010000000100010011;
ROM[43656] <= 32'b00000000000000011010001110000011;
ROM[43657] <= 32'b00000000011100010010000000100011;
ROM[43658] <= 32'b00000000010000010000000100010011;
ROM[43659] <= 32'b00000000101000000000001110010011;
ROM[43660] <= 32'b00000000011100010010000000100011;
ROM[43661] <= 32'b00000000010000010000000100010011;
ROM[43662] <= 32'b00000000000000101011001110110111;
ROM[43663] <= 32'b10101000010000111000001110010011;
ROM[43664] <= 32'b00000000111000111000001110110011;
ROM[43665] <= 32'b00000000011100010010000000100011;
ROM[43666] <= 32'b00000000010000010000000100010011;
ROM[43667] <= 32'b00000000001100010010000000100011;
ROM[43668] <= 32'b00000000010000010000000100010011;
ROM[43669] <= 32'b00000000010000010010000000100011;
ROM[43670] <= 32'b00000000010000010000000100010011;
ROM[43671] <= 32'b00000000010100010010000000100011;
ROM[43672] <= 32'b00000000010000010000000100010011;
ROM[43673] <= 32'b00000000011000010010000000100011;
ROM[43674] <= 32'b00000000010000010000000100010011;
ROM[43675] <= 32'b00000001010000000000001110010011;
ROM[43676] <= 32'b00000000100000111000001110010011;
ROM[43677] <= 32'b01000000011100010000001110110011;
ROM[43678] <= 32'b00000000011100000000001000110011;
ROM[43679] <= 32'b00000000001000000000000110110011;
ROM[43680] <= 32'b11011010110111100110000011101111;
ROM[43681] <= 32'b11111111110000010000000100010011;
ROM[43682] <= 32'b00000000000000010010001110000011;
ROM[43683] <= 32'b11111111110000010000000100010011;
ROM[43684] <= 32'b00000000000000010010010000000011;
ROM[43685] <= 32'b01000000011101000000001110110011;
ROM[43686] <= 32'b00000000011100010010000000100011;
ROM[43687] <= 32'b00000000010000010000000100010011;
ROM[43688] <= 32'b00000000000000101011001110110111;
ROM[43689] <= 32'b10101110110000111000001110010011;
ROM[43690] <= 32'b00000000111000111000001110110011;
ROM[43691] <= 32'b00000000011100010010000000100011;
ROM[43692] <= 32'b00000000010000010000000100010011;
ROM[43693] <= 32'b00000000001100010010000000100011;
ROM[43694] <= 32'b00000000010000010000000100010011;
ROM[43695] <= 32'b00000000010000010010000000100011;
ROM[43696] <= 32'b00000000010000010000000100010011;
ROM[43697] <= 32'b00000000010100010010000000100011;
ROM[43698] <= 32'b00000000010000010000000100010011;
ROM[43699] <= 32'b00000000011000010010000000100011;
ROM[43700] <= 32'b00000000010000010000000100010011;
ROM[43701] <= 32'b00000001010000000000001110010011;
ROM[43702] <= 32'b00000000010000111000001110010011;
ROM[43703] <= 32'b01000000011100010000001110110011;
ROM[43704] <= 32'b00000000011100000000001000110011;
ROM[43705] <= 32'b00000000001000000000000110110011;
ROM[43706] <= 32'b10101100010111111111000011101111;
ROM[43707] <= 32'b00000000000000101011001110110111;
ROM[43708] <= 32'b10110011100000111000001110010011;
ROM[43709] <= 32'b00000000111000111000001110110011;
ROM[43710] <= 32'b00000000011100010010000000100011;
ROM[43711] <= 32'b00000000010000010000000100010011;
ROM[43712] <= 32'b00000000001100010010000000100011;
ROM[43713] <= 32'b00000000010000010000000100010011;
ROM[43714] <= 32'b00000000010000010010000000100011;
ROM[43715] <= 32'b00000000010000010000000100010011;
ROM[43716] <= 32'b00000000010100010010000000100011;
ROM[43717] <= 32'b00000000010000010000000100010011;
ROM[43718] <= 32'b00000000011000010010000000100011;
ROM[43719] <= 32'b00000000010000010000000100010011;
ROM[43720] <= 32'b00000001010000000000001110010011;
ROM[43721] <= 32'b00000000100000111000001110010011;
ROM[43722] <= 32'b01000000011100010000001110110011;
ROM[43723] <= 32'b00000000011100000000001000110011;
ROM[43724] <= 32'b00000000001000000000000110110011;
ROM[43725] <= 32'b10000111100011111111000011101111;
ROM[43726] <= 32'b11111111110000010000000100010011;
ROM[43727] <= 32'b00000000000000010010001110000011;
ROM[43728] <= 32'b00000000011101100010000000100011;
ROM[43729] <= 32'b00001011110000000000000011101111;
ROM[43730] <= 32'b00000000010100010010000000100011;
ROM[43731] <= 32'b00000000010000010000000100010011;
ROM[43732] <= 32'b00000000010000100010001110000011;
ROM[43733] <= 32'b00000000011100010010000000100011;
ROM[43734] <= 32'b00000000010000010000000100010011;
ROM[43735] <= 32'b00000000000000101011001110110111;
ROM[43736] <= 32'b10111010100000111000001110010011;
ROM[43737] <= 32'b00000000111000111000001110110011;
ROM[43738] <= 32'b00000000011100010010000000100011;
ROM[43739] <= 32'b00000000010000010000000100010011;
ROM[43740] <= 32'b00000000001100010010000000100011;
ROM[43741] <= 32'b00000000010000010000000100010011;
ROM[43742] <= 32'b00000000010000010010000000100011;
ROM[43743] <= 32'b00000000010000010000000100010011;
ROM[43744] <= 32'b00000000010100010010000000100011;
ROM[43745] <= 32'b00000000010000010000000100010011;
ROM[43746] <= 32'b00000000011000010010000000100011;
ROM[43747] <= 32'b00000000010000010000000100010011;
ROM[43748] <= 32'b00000001010000000000001110010011;
ROM[43749] <= 32'b00000000010000111000001110010011;
ROM[43750] <= 32'b01000000011100010000001110110011;
ROM[43751] <= 32'b00000000011100000000001000110011;
ROM[43752] <= 32'b00000000001000000000000110110011;
ROM[43753] <= 32'b10100000100111111111000011101111;
ROM[43754] <= 32'b00000000000000101011001110110111;
ROM[43755] <= 32'b10111111010000111000001110010011;
ROM[43756] <= 32'b00000000111000111000001110110011;
ROM[43757] <= 32'b00000000011100010010000000100011;
ROM[43758] <= 32'b00000000010000010000000100010011;
ROM[43759] <= 32'b00000000001100010010000000100011;
ROM[43760] <= 32'b00000000010000010000000100010011;
ROM[43761] <= 32'b00000000010000010010000000100011;
ROM[43762] <= 32'b00000000010000010000000100010011;
ROM[43763] <= 32'b00000000010100010010000000100011;
ROM[43764] <= 32'b00000000010000010000000100010011;
ROM[43765] <= 32'b00000000011000010010000000100011;
ROM[43766] <= 32'b00000000010000010000000100010011;
ROM[43767] <= 32'b00000001010000000000001110010011;
ROM[43768] <= 32'b00000000100000111000001110010011;
ROM[43769] <= 32'b01000000011100010000001110110011;
ROM[43770] <= 32'b00000000011100000000001000110011;
ROM[43771] <= 32'b00000000001000000000000110110011;
ROM[43772] <= 32'b11111011110111111110000011101111;
ROM[43773] <= 32'b11111111110000010000000100010011;
ROM[43774] <= 32'b00000000000000010010001110000011;
ROM[43775] <= 32'b00000000011101100010000000100011;
ROM[43776] <= 32'b00000000000000000000001110010011;
ROM[43777] <= 32'b00000000011100010010000000100011;
ROM[43778] <= 32'b00000000010000010000000100010011;
ROM[43779] <= 32'b00000001010000000000001110010011;
ROM[43780] <= 32'b01000000011100011000001110110011;
ROM[43781] <= 32'b00000000000000111010000010000011;
ROM[43782] <= 32'b11111111110000010000000100010011;
ROM[43783] <= 32'b00000000000000010010001110000011;
ROM[43784] <= 32'b00000000011100100010000000100011;
ROM[43785] <= 32'b00000000010000100000000100010011;
ROM[43786] <= 32'b00000001010000000000001110010011;
ROM[43787] <= 32'b01000000011100011000001110110011;
ROM[43788] <= 32'b00000000010000111010000110000011;
ROM[43789] <= 32'b00000000100000111010001000000011;
ROM[43790] <= 32'b00000000110000111010001010000011;
ROM[43791] <= 32'b00000001000000111010001100000011;
ROM[43792] <= 32'b00000000000000001000000011100111;
ROM[43793] <= 32'b00000000110100000000001110010011;
ROM[43794] <= 32'b00000000011100010010000000100011;
ROM[43795] <= 32'b00000000010000010000000100010011;
ROM[43796] <= 32'b00000001010000000000001110010011;
ROM[43797] <= 32'b01000000011100011000001110110011;
ROM[43798] <= 32'b00000000000000111010000010000011;
ROM[43799] <= 32'b11111111110000010000000100010011;
ROM[43800] <= 32'b00000000000000010010001110000011;
ROM[43801] <= 32'b00000000011100100010000000100011;
ROM[43802] <= 32'b00000000010000100000000100010011;
ROM[43803] <= 32'b00000001010000000000001110010011;
ROM[43804] <= 32'b01000000011100011000001110110011;
ROM[43805] <= 32'b00000000010000111010000110000011;
ROM[43806] <= 32'b00000000100000111010001000000011;
ROM[43807] <= 32'b00000000110000111010001010000011;
ROM[43808] <= 32'b00000001000000111010001100000011;
ROM[43809] <= 32'b00000000000000001000000011100111;
ROM[43810] <= 32'b00000000100000000000001110010011;
ROM[43811] <= 32'b00000000011100010010000000100011;
ROM[43812] <= 32'b00000000010000010000000100010011;
ROM[43813] <= 32'b00000001010000000000001110010011;
ROM[43814] <= 32'b01000000011100011000001110110011;
ROM[43815] <= 32'b00000000000000111010000010000011;
ROM[43816] <= 32'b11111111110000010000000100010011;
ROM[43817] <= 32'b00000000000000010010001110000011;
ROM[43818] <= 32'b00000000011100100010000000100011;
ROM[43819] <= 32'b00000000010000100000000100010011;
ROM[43820] <= 32'b00000001010000000000001110010011;
ROM[43821] <= 32'b01000000011100011000001110110011;
ROM[43822] <= 32'b00000000010000111010000110000011;
ROM[43823] <= 32'b00000000100000111010001000000011;
ROM[43824] <= 32'b00000000110000111010001010000011;
ROM[43825] <= 32'b00000001000000111010001100000011;
ROM[43826] <= 32'b00000000000000001000000011100111;
ROM[43827] <= 32'b00000010001000000000001110010011;
ROM[43828] <= 32'b00000000011100010010000000100011;
ROM[43829] <= 32'b00000000010000010000000100010011;
ROM[43830] <= 32'b00000001010000000000001110010011;
ROM[43831] <= 32'b01000000011100011000001110110011;
ROM[43832] <= 32'b00000000000000111010000010000011;
ROM[43833] <= 32'b11111111110000010000000100010011;
ROM[43834] <= 32'b00000000000000010010001110000011;
ROM[43835] <= 32'b00000000011100100010000000100011;
ROM[43836] <= 32'b00000000010000100000000100010011;
ROM[43837] <= 32'b00000001010000000000001110010011;
ROM[43838] <= 32'b01000000011100011000001110110011;
ROM[43839] <= 32'b00000000010000111010000110000011;
ROM[43840] <= 32'b00000000100000111010001000000011;
ROM[43841] <= 32'b00000000110000111010001010000011;
ROM[43842] <= 32'b00000001000000111010001100000011;
ROM[43843] <= 32'b00000000000000001000000011100111;
ROM[43844] <= 32'b00000000000000100010001110000011;
ROM[43845] <= 32'b00000000011100010010000000100011;
ROM[43846] <= 32'b00000000010000010000000100010011;
ROM[43847] <= 32'b11111111110000010000000100010011;
ROM[43848] <= 32'b00000000000000010010001110000011;
ROM[43849] <= 32'b00000000000000111000001010010011;
ROM[43850] <= 32'b00000000110100101000010000110011;
ROM[43851] <= 32'b00000000100001000010001110000011;
ROM[43852] <= 32'b00000000011100010010000000100011;
ROM[43853] <= 32'b00000000010000010000000100010011;
ROM[43854] <= 32'b00000000000000101011001110110111;
ROM[43855] <= 32'b11011000010000111000001110010011;
ROM[43856] <= 32'b00000000111000111000001110110011;
ROM[43857] <= 32'b00000000011100010010000000100011;
ROM[43858] <= 32'b00000000010000010000000100010011;
ROM[43859] <= 32'b00000000001100010010000000100011;
ROM[43860] <= 32'b00000000010000010000000100010011;
ROM[43861] <= 32'b00000000010000010010000000100011;
ROM[43862] <= 32'b00000000010000010000000100010011;
ROM[43863] <= 32'b00000000010100010010000000100011;
ROM[43864] <= 32'b00000000010000010000000100010011;
ROM[43865] <= 32'b00000000011000010010000000100011;
ROM[43866] <= 32'b00000000010000010000000100010011;
ROM[43867] <= 32'b00000001010000000000001110010011;
ROM[43868] <= 32'b00000000010000111000001110010011;
ROM[43869] <= 32'b01000000011100010000001110110011;
ROM[43870] <= 32'b00000000011100000000001000110011;
ROM[43871] <= 32'b00000000001000000000000110110011;
ROM[43872] <= 32'b10111001000011010101000011101111;
ROM[43873] <= 32'b11111111110000010000000100010011;
ROM[43874] <= 32'b00000000000000010010001110000011;
ROM[43875] <= 32'b00000000011101100010000000100011;
ROM[43876] <= 32'b00000000000000000000001110010011;
ROM[43877] <= 32'b00000000011100010010000000100011;
ROM[43878] <= 32'b00000000010000010000000100010011;
ROM[43879] <= 32'b00000001010000000000001110010011;
ROM[43880] <= 32'b01000000011100011000001110110011;
ROM[43881] <= 32'b00000000000000111010000010000011;
ROM[43882] <= 32'b11111111110000010000000100010011;
ROM[43883] <= 32'b00000000000000010010001110000011;
ROM[43884] <= 32'b00000000011100100010000000100011;
ROM[43885] <= 32'b00000000010000100000000100010011;
ROM[43886] <= 32'b00000001010000000000001110010011;
ROM[43887] <= 32'b01000000011100011000001110110011;
ROM[43888] <= 32'b00000000010000111010000110000011;
ROM[43889] <= 32'b00000000100000111010001000000011;
ROM[43890] <= 32'b00000000110000111010001010000011;
ROM[43891] <= 32'b00000001000000111010001100000011;
ROM[43892] <= 32'b00000000000000001000000011100111;
ROM[43893] <= 32'b00000000000000101011001110110111;
ROM[43894] <= 32'b11100010000000111000001110010011;
ROM[43895] <= 32'b00000000111000111000001110110011;
ROM[43896] <= 32'b00000000011100010010000000100011;
ROM[43897] <= 32'b00000000010000010000000100010011;
ROM[43898] <= 32'b00000000001100010010000000100011;
ROM[43899] <= 32'b00000000010000010000000100010011;
ROM[43900] <= 32'b00000000010000010010000000100011;
ROM[43901] <= 32'b00000000010000010000000100010011;
ROM[43902] <= 32'b00000000010100010010000000100011;
ROM[43903] <= 32'b00000000010000010000000100010011;
ROM[43904] <= 32'b00000000011000010010000000100011;
ROM[43905] <= 32'b00000000010000010000000100010011;
ROM[43906] <= 32'b00000001010000000000001110010011;
ROM[43907] <= 32'b00000000000000111000001110010011;
ROM[43908] <= 32'b01000000011100010000001110110011;
ROM[43909] <= 32'b00000000011100000000001000110011;
ROM[43910] <= 32'b00000000001000000000000110110011;
ROM[43911] <= 32'b11000100100011101000000011101111;
ROM[43912] <= 32'b11111111110000010000000100010011;
ROM[43913] <= 32'b00000000000000010010001110000011;
ROM[43914] <= 32'b00000000011101100010000000100011;
ROM[43915] <= 32'b00000000000000101011001110110111;
ROM[43916] <= 32'b11100111100000111000001110010011;
ROM[43917] <= 32'b00000000111000111000001110110011;
ROM[43918] <= 32'b00000000011100010010000000100011;
ROM[43919] <= 32'b00000000010000010000000100010011;
ROM[43920] <= 32'b00000000001100010010000000100011;
ROM[43921] <= 32'b00000000010000010000000100010011;
ROM[43922] <= 32'b00000000010000010010000000100011;
ROM[43923] <= 32'b00000000010000010000000100010011;
ROM[43924] <= 32'b00000000010100010010000000100011;
ROM[43925] <= 32'b00000000010000010000000100010011;
ROM[43926] <= 32'b00000000011000010010000000100011;
ROM[43927] <= 32'b00000000010000010000000100010011;
ROM[43928] <= 32'b00000001010000000000001110010011;
ROM[43929] <= 32'b00000000000000111000001110010011;
ROM[43930] <= 32'b01000000011100010000001110110011;
ROM[43931] <= 32'b00000000011100000000001000110011;
ROM[43932] <= 32'b00000000001000000000000110110011;
ROM[43933] <= 32'b10100101000011100101000011101111;
ROM[43934] <= 32'b11111111110000010000000100010011;
ROM[43935] <= 32'b00000000000000010010001110000011;
ROM[43936] <= 32'b00000000011101100010000000100011;
ROM[43937] <= 32'b00000000000000101011001110110111;
ROM[43938] <= 32'b11101101000000111000001110010011;
ROM[43939] <= 32'b00000000111000111000001110110011;
ROM[43940] <= 32'b00000000011100010010000000100011;
ROM[43941] <= 32'b00000000010000010000000100010011;
ROM[43942] <= 32'b00000000001100010010000000100011;
ROM[43943] <= 32'b00000000010000010000000100010011;
ROM[43944] <= 32'b00000000010000010010000000100011;
ROM[43945] <= 32'b00000000010000010000000100010011;
ROM[43946] <= 32'b00000000010100010010000000100011;
ROM[43947] <= 32'b00000000010000010000000100010011;
ROM[43948] <= 32'b00000000011000010010000000100011;
ROM[43949] <= 32'b00000000010000010000000100010011;
ROM[43950] <= 32'b00000001010000000000001110010011;
ROM[43951] <= 32'b00000000000000111000001110010011;
ROM[43952] <= 32'b01000000011100010000001110110011;
ROM[43953] <= 32'b00000000011100000000001000110011;
ROM[43954] <= 32'b00000000001000000000000110110011;
ROM[43955] <= 32'b11101010110111101001000011101111;
ROM[43956] <= 32'b11111111110000010000000100010011;
ROM[43957] <= 32'b00000000000000010010001110000011;
ROM[43958] <= 32'b00000000011101100010000000100011;
ROM[43959] <= 32'b00000000000000101011001110110111;
ROM[43960] <= 32'b11110010100000111000001110010011;
ROM[43961] <= 32'b00000000111000111000001110110011;
ROM[43962] <= 32'b00000000011100010010000000100011;
ROM[43963] <= 32'b00000000010000010000000100010011;
ROM[43964] <= 32'b00000000001100010010000000100011;
ROM[43965] <= 32'b00000000010000010000000100010011;
ROM[43966] <= 32'b00000000010000010010000000100011;
ROM[43967] <= 32'b00000000010000010000000100010011;
ROM[43968] <= 32'b00000000010100010010000000100011;
ROM[43969] <= 32'b00000000010000010000000100010011;
ROM[43970] <= 32'b00000000011000010010000000100011;
ROM[43971] <= 32'b00000000010000010000000100010011;
ROM[43972] <= 32'b00000001010000000000001110010011;
ROM[43973] <= 32'b00000000000000111000001110010011;
ROM[43974] <= 32'b01000000011100010000001110110011;
ROM[43975] <= 32'b00000000011100000000001000110011;
ROM[43976] <= 32'b00000000001000000000000110110011;
ROM[43977] <= 32'b10000100010111100010000011101111;
ROM[43978] <= 32'b11111111110000010000000100010011;
ROM[43979] <= 32'b00000000000000010010001110000011;
ROM[43980] <= 32'b00000000011101100010000000100011;
ROM[43981] <= 32'b00000000000000101011001110110111;
ROM[43982] <= 32'b11111000000000111000001110010011;
ROM[43983] <= 32'b00000000111000111000001110110011;
ROM[43984] <= 32'b00000000011100010010000000100011;
ROM[43985] <= 32'b00000000010000010000000100010011;
ROM[43986] <= 32'b00000000001100010010000000100011;
ROM[43987] <= 32'b00000000010000010000000100010011;
ROM[43988] <= 32'b00000000010000010010000000100011;
ROM[43989] <= 32'b00000000010000010000000100010011;
ROM[43990] <= 32'b00000000010100010010000000100011;
ROM[43991] <= 32'b00000000010000010000000100010011;
ROM[43992] <= 32'b00000000011000010010000000100011;
ROM[43993] <= 32'b00000000010000010000000100010011;
ROM[43994] <= 32'b00000001010000000000001110010011;
ROM[43995] <= 32'b00000000000000111000001110010011;
ROM[43996] <= 32'b01000000011100010000001110110011;
ROM[43997] <= 32'b00000000011100000000001000110011;
ROM[43998] <= 32'b00000000001000000000000110110011;
ROM[43999] <= 32'b11010000000111110010000011101111;
ROM[44000] <= 32'b11111111110000010000000100010011;
ROM[44001] <= 32'b00000000000000010010001110000011;
ROM[44002] <= 32'b00000000011101100010000000100011;
ROM[44003] <= 32'b00000000000000101011001110110111;
ROM[44004] <= 32'b11111101100000111000001110010011;
ROM[44005] <= 32'b00000000111000111000001110110011;
ROM[44006] <= 32'b00000000011100010010000000100011;
ROM[44007] <= 32'b00000000010000010000000100010011;
ROM[44008] <= 32'b00000000001100010010000000100011;
ROM[44009] <= 32'b00000000010000010000000100010011;
ROM[44010] <= 32'b00000000010000010010000000100011;
ROM[44011] <= 32'b00000000010000010000000100010011;
ROM[44012] <= 32'b00000000010100010010000000100011;
ROM[44013] <= 32'b00000000010000010000000100010011;
ROM[44014] <= 32'b00000000011000010010000000100011;
ROM[44015] <= 32'b00000000010000010000000100010011;
ROM[44016] <= 32'b00000001010000000000001110010011;
ROM[44017] <= 32'b00000000000000111000001110010011;
ROM[44018] <= 32'b01000000011100010000001110110011;
ROM[44019] <= 32'b00000000011100000000001000110011;
ROM[44020] <= 32'b00000000001000000000000110110011;
ROM[44021] <= 32'b01010100100000000000000011101111;
ROM[44022] <= 32'b11111111110000010000000100010011;
ROM[44023] <= 32'b00000000000000010010001110000011;
ROM[44024] <= 32'b00000000011101100010000000100011;
ROM[44025] <= 32'b00000000000000000000001110010011;
ROM[44026] <= 32'b00000000011100010010000000100011;
ROM[44027] <= 32'b00000000010000010000000100010011;
ROM[44028] <= 32'b00000001010000000000001110010011;
ROM[44029] <= 32'b01000000011100011000001110110011;
ROM[44030] <= 32'b00000000000000111010000010000011;
ROM[44031] <= 32'b11111111110000010000000100010011;
ROM[44032] <= 32'b00000000000000010010001110000011;
ROM[44033] <= 32'b00000000011100100010000000100011;
ROM[44034] <= 32'b00000000010000100000000100010011;
ROM[44035] <= 32'b00000001010000000000001110010011;
ROM[44036] <= 32'b01000000011100011000001110110011;
ROM[44037] <= 32'b00000000010000111010000110000011;
ROM[44038] <= 32'b00000000100000111010001000000011;
ROM[44039] <= 32'b00000000110000111010001010000011;
ROM[44040] <= 32'b00000001000000111010001100000011;
ROM[44041] <= 32'b00000000000000001000000011100111;
ROM[44042] <= 32'b00000000000100000000001110010011;
ROM[44043] <= 32'b00000000011100010010000000100011;
ROM[44044] <= 32'b00000000010000010000000100010011;
ROM[44045] <= 32'b11111111110000010000000100010011;
ROM[44046] <= 32'b00000000000000010010001110000011;
ROM[44047] <= 32'b01000000011100000000001110110011;
ROM[44048] <= 32'b00000000011100010010000000100011;
ROM[44049] <= 32'b00000000010000010000000100010011;
ROM[44050] <= 32'b11111111110000010000000100010011;
ROM[44051] <= 32'b00000000000000010010001110000011;
ROM[44052] <= 32'b01000000011100000000001110110011;
ROM[44053] <= 32'b00000000000100111000001110010011;
ROM[44054] <= 32'b00000000011100010010000000100011;
ROM[44055] <= 32'b00000000010000010000000100010011;
ROM[44056] <= 32'b11111111110000010000000100010011;
ROM[44057] <= 32'b00000000000000010010001110000011;
ROM[44058] <= 32'b00000000000000111000101001100011;
ROM[44059] <= 32'b00000000000000101011001110110111;
ROM[44060] <= 32'b00001000000000111000001110010011;
ROM[44061] <= 32'b00000000111000111000001110110011;
ROM[44062] <= 32'b00000000000000111000000011100111;
ROM[44063] <= 32'b11111010110111111111000011101111;
ROM[44064] <= 32'b00000000000000000000001110010011;
ROM[44065] <= 32'b00000000011100010010000000100011;
ROM[44066] <= 32'b00000000010000010000000100010011;
ROM[44067] <= 32'b00000001010000000000001110010011;
ROM[44068] <= 32'b01000000011100011000001110110011;
ROM[44069] <= 32'b00000000000000111010000010000011;
ROM[44070] <= 32'b11111111110000010000000100010011;
ROM[44071] <= 32'b00000000000000010010001110000011;
ROM[44072] <= 32'b00000000011100100010000000100011;
ROM[44073] <= 32'b00000000010000100000000100010011;
ROM[44074] <= 32'b00000001010000000000001110010011;
ROM[44075] <= 32'b01000000011100011000001110110011;
ROM[44076] <= 32'b00000000010000111010000110000011;
ROM[44077] <= 32'b00000000100000111010001000000011;
ROM[44078] <= 32'b00000000110000111010001010000011;
ROM[44079] <= 32'b00000001000000111010001100000011;
ROM[44080] <= 32'b00000000000000001000000011100111;
ROM[44081] <= 32'b00000000000000010010000000100011;
ROM[44082] <= 32'b00000000010000010000000100010011;
ROM[44083] <= 32'b00000000000000010010000000100011;
ROM[44084] <= 32'b00000000010000010000000100010011;
ROM[44085] <= 32'b00000000000000000000001110010011;
ROM[44086] <= 32'b00000000011100010010000000100011;
ROM[44087] <= 32'b00000000010000010000000100010011;
ROM[44088] <= 32'b11111111110000010000000100010011;
ROM[44089] <= 32'b00000000000000010010001110000011;
ROM[44090] <= 32'b00000000011100011010000000100011;
ROM[44091] <= 32'b00000000000000011010001110000011;
ROM[44092] <= 32'b00000000011100010010000000100011;
ROM[44093] <= 32'b00000000010000010000000100010011;
ROM[44094] <= 32'b00000000000000100010001110000011;
ROM[44095] <= 32'b00000000011100010010000000100011;
ROM[44096] <= 32'b00000000010000010000000100010011;
ROM[44097] <= 32'b11111111110000010000000100010011;
ROM[44098] <= 32'b00000000000000010010001110000011;
ROM[44099] <= 32'b11111111110000010000000100010011;
ROM[44100] <= 32'b00000000000000010010010000000011;
ROM[44101] <= 32'b00000000011101000010001110110011;
ROM[44102] <= 32'b00000000011100010010000000100011;
ROM[44103] <= 32'b00000000010000010000000100010011;
ROM[44104] <= 32'b11111111110000010000000100010011;
ROM[44105] <= 32'b00000000000000010010001110000011;
ROM[44106] <= 32'b01000000011100000000001110110011;
ROM[44107] <= 32'b00000000000100111000001110010011;
ROM[44108] <= 32'b00000000011100010010000000100011;
ROM[44109] <= 32'b00000000010000010000000100010011;
ROM[44110] <= 32'b11111111110000010000000100010011;
ROM[44111] <= 32'b00000000000000010010001110000011;
ROM[44112] <= 32'b00000000000000111000101001100011;
ROM[44113] <= 32'b00000000000000101011001110110111;
ROM[44114] <= 32'b00100101110000111000001110010011;
ROM[44115] <= 32'b00000000111000111000001110110011;
ROM[44116] <= 32'b00000000000000111000000011100111;
ROM[44117] <= 32'b00000000000000000000001110010011;
ROM[44118] <= 32'b00000000011100010010000000100011;
ROM[44119] <= 32'b00000000010000010000000100010011;
ROM[44120] <= 32'b11111111110000010000000100010011;
ROM[44121] <= 32'b00000000000000010010001110000011;
ROM[44122] <= 32'b00000000011100011010001000100011;
ROM[44123] <= 32'b00000000010000011010001110000011;
ROM[44124] <= 32'b00000000011100010010000000100011;
ROM[44125] <= 32'b00000000010000010000000100010011;
ROM[44126] <= 32'b00000110010000000000001110010011;
ROM[44127] <= 32'b00000000011100010010000000100011;
ROM[44128] <= 32'b00000000010000010000000100010011;
ROM[44129] <= 32'b11111111110000010000000100010011;
ROM[44130] <= 32'b00000000000000010010001110000011;
ROM[44131] <= 32'b11111111110000010000000100010011;
ROM[44132] <= 32'b00000000000000010010010000000011;
ROM[44133] <= 32'b00000000011101000010001110110011;
ROM[44134] <= 32'b00000000011100010010000000100011;
ROM[44135] <= 32'b00000000010000010000000100010011;
ROM[44136] <= 32'b11111111110000010000000100010011;
ROM[44137] <= 32'b00000000000000010010001110000011;
ROM[44138] <= 32'b01000000011100000000001110110011;
ROM[44139] <= 32'b00000000000100111000001110010011;
ROM[44140] <= 32'b00000000011100010010000000100011;
ROM[44141] <= 32'b00000000010000010000000100010011;
ROM[44142] <= 32'b11111111110000010000000100010011;
ROM[44143] <= 32'b00000000000000010010001110000011;
ROM[44144] <= 32'b00000000000000111000101001100011;
ROM[44145] <= 32'b00000000000000101011001110110111;
ROM[44146] <= 32'b00100001100000111000001110010011;
ROM[44147] <= 32'b00000000111000111000001110110011;
ROM[44148] <= 32'b00000000000000111000000011100111;
ROM[44149] <= 32'b00000000010000011010001110000011;
ROM[44150] <= 32'b00000000011100010010000000100011;
ROM[44151] <= 32'b00000000010000010000000100010011;
ROM[44152] <= 32'b00000000000100000000001110010011;
ROM[44153] <= 32'b00000000011100010010000000100011;
ROM[44154] <= 32'b00000000010000010000000100010011;
ROM[44155] <= 32'b11111111110000010000000100010011;
ROM[44156] <= 32'b00000000000000010010001110000011;
ROM[44157] <= 32'b11111111110000010000000100010011;
ROM[44158] <= 32'b00000000000000010010010000000011;
ROM[44159] <= 32'b00000000011101000000001110110011;
ROM[44160] <= 32'b00000000011100010010000000100011;
ROM[44161] <= 32'b00000000010000010000000100010011;
ROM[44162] <= 32'b11111111110000010000000100010011;
ROM[44163] <= 32'b00000000000000010010001110000011;
ROM[44164] <= 32'b00000000011100011010001000100011;
ROM[44165] <= 32'b11110101100111111111000011101111;
ROM[44166] <= 32'b00000000000000011010001110000011;
ROM[44167] <= 32'b00000000011100010010000000100011;
ROM[44168] <= 32'b00000000010000010000000100010011;
ROM[44169] <= 32'b00000000000100000000001110010011;
ROM[44170] <= 32'b00000000011100010010000000100011;
ROM[44171] <= 32'b00000000010000010000000100010011;
ROM[44172] <= 32'b11111111110000010000000100010011;
ROM[44173] <= 32'b00000000000000010010001110000011;
ROM[44174] <= 32'b11111111110000010000000100010011;
ROM[44175] <= 32'b00000000000000010010010000000011;
ROM[44176] <= 32'b00000000011101000000001110110011;
ROM[44177] <= 32'b00000000011100010010000000100011;
ROM[44178] <= 32'b00000000010000010000000100010011;
ROM[44179] <= 32'b11111111110000010000000100010011;
ROM[44180] <= 32'b00000000000000010010001110000011;
ROM[44181] <= 32'b00000000011100011010000000100011;
ROM[44182] <= 32'b11101001010111111111000011101111;
ROM[44183] <= 32'b00000000000000000000001110010011;
ROM[44184] <= 32'b00000000011100010010000000100011;
ROM[44185] <= 32'b00000000010000010000000100010011;
ROM[44186] <= 32'b00000001010000000000001110010011;
ROM[44187] <= 32'b01000000011100011000001110110011;
ROM[44188] <= 32'b00000000000000111010000010000011;
ROM[44189] <= 32'b11111111110000010000000100010011;
ROM[44190] <= 32'b00000000000000010010001110000011;
ROM[44191] <= 32'b00000000011100100010000000100011;
ROM[44192] <= 32'b00000000010000100000000100010011;
ROM[44193] <= 32'b00000001010000000000001110010011;
ROM[44194] <= 32'b01000000011100011000001110110011;
ROM[44195] <= 32'b00000000010000111010000110000011;
ROM[44196] <= 32'b00000000100000111010001000000011;
ROM[44197] <= 32'b00000000110000111010001010000011;
ROM[44198] <= 32'b00000001000000111010001100000011;
ROM[44199] <= 32'b00000000000000001000000011100111;
ROM[44200] <= 32'b00000000000000010010000000100011;
ROM[44201] <= 32'b00000000010000010000000100010011;
ROM[44202] <= 32'b00000000000000010010000000100011;
ROM[44203] <= 32'b00000000010000010000000100010011;
ROM[44204] <= 32'b00000000010000000000001110010011;
ROM[44205] <= 32'b00000000011100010010000000100011;
ROM[44206] <= 32'b00000000010000010000000100010011;
ROM[44207] <= 32'b00000000000000101011001110110111;
ROM[44208] <= 32'b00110000100000111000001110010011;
ROM[44209] <= 32'b00000000111000111000001110110011;
ROM[44210] <= 32'b00000000011100010010000000100011;
ROM[44211] <= 32'b00000000010000010000000100010011;
ROM[44212] <= 32'b00000000001100010010000000100011;
ROM[44213] <= 32'b00000000010000010000000100010011;
ROM[44214] <= 32'b00000000010000010010000000100011;
ROM[44215] <= 32'b00000000010000010000000100010011;
ROM[44216] <= 32'b00000000010100010010000000100011;
ROM[44217] <= 32'b00000000010000010000000100010011;
ROM[44218] <= 32'b00000000011000010010000000100011;
ROM[44219] <= 32'b00000000010000010000000100010011;
ROM[44220] <= 32'b00000001010000000000001110010011;
ROM[44221] <= 32'b00000000010000111000001110010011;
ROM[44222] <= 32'b01000000011100010000001110110011;
ROM[44223] <= 32'b00000000011100000000001000110011;
ROM[44224] <= 32'b00000000001000000000000110110011;
ROM[44225] <= 32'b11000011100011111110000011101111;
ROM[44226] <= 32'b00000100000100000000001110010011;
ROM[44227] <= 32'b00000000011100010010000000100011;
ROM[44228] <= 32'b00000000010000010000000100010011;
ROM[44229] <= 32'b00000000000000101011001110110111;
ROM[44230] <= 32'b00110110000000111000001110010011;
ROM[44231] <= 32'b00000000111000111000001110110011;
ROM[44232] <= 32'b00000000011100010010000000100011;
ROM[44233] <= 32'b00000000010000010000000100010011;
ROM[44234] <= 32'b00000000001100010010000000100011;
ROM[44235] <= 32'b00000000010000010000000100010011;
ROM[44236] <= 32'b00000000010000010010000000100011;
ROM[44237] <= 32'b00000000010000010000000100010011;
ROM[44238] <= 32'b00000000010100010010000000100011;
ROM[44239] <= 32'b00000000010000010000000100010011;
ROM[44240] <= 32'b00000000011000010010000000100011;
ROM[44241] <= 32'b00000000010000010000000100010011;
ROM[44242] <= 32'b00000001010000000000001110010011;
ROM[44243] <= 32'b00000000100000111000001110010011;
ROM[44244] <= 32'b01000000011100010000001110110011;
ROM[44245] <= 32'b00000000011100000000001000110011;
ROM[44246] <= 32'b00000000001000000000000110110011;
ROM[44247] <= 32'b10000101000111111110000011101111;
ROM[44248] <= 32'b00000100001000000000001110010011;
ROM[44249] <= 32'b00000000011100010010000000100011;
ROM[44250] <= 32'b00000000010000010000000100010011;
ROM[44251] <= 32'b00000000000000101011001110110111;
ROM[44252] <= 32'b00111011100000111000001110010011;
ROM[44253] <= 32'b00000000111000111000001110110011;
ROM[44254] <= 32'b00000000011100010010000000100011;
ROM[44255] <= 32'b00000000010000010000000100010011;
ROM[44256] <= 32'b00000000001100010010000000100011;
ROM[44257] <= 32'b00000000010000010000000100010011;
ROM[44258] <= 32'b00000000010000010010000000100011;
ROM[44259] <= 32'b00000000010000010000000100010011;
ROM[44260] <= 32'b00000000010100010010000000100011;
ROM[44261] <= 32'b00000000010000010000000100010011;
ROM[44262] <= 32'b00000000011000010010000000100011;
ROM[44263] <= 32'b00000000010000010000000100010011;
ROM[44264] <= 32'b00000001010000000000001110010011;
ROM[44265] <= 32'b00000000100000111000001110010011;
ROM[44266] <= 32'b01000000011100010000001110110011;
ROM[44267] <= 32'b00000000011100000000001000110011;
ROM[44268] <= 32'b00000000001000000000000110110011;
ROM[44269] <= 32'b11111111100011111110000011101111;
ROM[44270] <= 32'b00000100001100000000001110010011;
ROM[44271] <= 32'b00000000011100010010000000100011;
ROM[44272] <= 32'b00000000010000010000000100010011;
ROM[44273] <= 32'b00000000000000101011001110110111;
ROM[44274] <= 32'b01000001000000111000001110010011;
ROM[44275] <= 32'b00000000111000111000001110110011;
ROM[44276] <= 32'b00000000011100010010000000100011;
ROM[44277] <= 32'b00000000010000010000000100010011;
ROM[44278] <= 32'b00000000001100010010000000100011;
ROM[44279] <= 32'b00000000010000010000000100010011;
ROM[44280] <= 32'b00000000010000010010000000100011;
ROM[44281] <= 32'b00000000010000010000000100010011;
ROM[44282] <= 32'b00000000010100010010000000100011;
ROM[44283] <= 32'b00000000010000010000000100010011;
ROM[44284] <= 32'b00000000011000010010000000100011;
ROM[44285] <= 32'b00000000010000010000000100010011;
ROM[44286] <= 32'b00000001010000000000001110010011;
ROM[44287] <= 32'b00000000100000111000001110010011;
ROM[44288] <= 32'b01000000011100010000001110110011;
ROM[44289] <= 32'b00000000011100000000001000110011;
ROM[44290] <= 32'b00000000001000000000000110110011;
ROM[44291] <= 32'b11111010000011111110000011101111;
ROM[44292] <= 32'b00000100010000000000001110010011;
ROM[44293] <= 32'b00000000011100010010000000100011;
ROM[44294] <= 32'b00000000010000010000000100010011;
ROM[44295] <= 32'b00000000000000101011001110110111;
ROM[44296] <= 32'b01000110100000111000001110010011;
ROM[44297] <= 32'b00000000111000111000001110110011;
ROM[44298] <= 32'b00000000011100010010000000100011;
ROM[44299] <= 32'b00000000010000010000000100010011;
ROM[44300] <= 32'b00000000001100010010000000100011;
ROM[44301] <= 32'b00000000010000010000000100010011;
ROM[44302] <= 32'b00000000010000010010000000100011;
ROM[44303] <= 32'b00000000010000010000000100010011;
ROM[44304] <= 32'b00000000010100010010000000100011;
ROM[44305] <= 32'b00000000010000010000000100010011;
ROM[44306] <= 32'b00000000011000010010000000100011;
ROM[44307] <= 32'b00000000010000010000000100010011;
ROM[44308] <= 32'b00000001010000000000001110010011;
ROM[44309] <= 32'b00000000100000111000001110010011;
ROM[44310] <= 32'b01000000011100010000001110110011;
ROM[44311] <= 32'b00000000011100000000001000110011;
ROM[44312] <= 32'b00000000001000000000000110110011;
ROM[44313] <= 32'b11110100100011111110000011101111;
ROM[44314] <= 32'b11111111110000010000000100010011;
ROM[44315] <= 32'b00000000000000010010001110000011;
ROM[44316] <= 32'b00000000011100011010001000100011;
ROM[44317] <= 32'b00000000010000011010001110000011;
ROM[44318] <= 32'b00000000011100010010000000100011;
ROM[44319] <= 32'b00000000010000010000000100010011;
ROM[44320] <= 32'b00000000000000101011001110110111;
ROM[44321] <= 32'b01001100110000111000001110010011;
ROM[44322] <= 32'b00000000111000111000001110110011;
ROM[44323] <= 32'b00000000011100010010000000100011;
ROM[44324] <= 32'b00000000010000010000000100010011;
ROM[44325] <= 32'b00000000001100010010000000100011;
ROM[44326] <= 32'b00000000010000010000000100010011;
ROM[44327] <= 32'b00000000010000010010000000100011;
ROM[44328] <= 32'b00000000010000010000000100010011;
ROM[44329] <= 32'b00000000010100010010000000100011;
ROM[44330] <= 32'b00000000010000010000000100010011;
ROM[44331] <= 32'b00000000011000010010000000100011;
ROM[44332] <= 32'b00000000010000010000000100010011;
ROM[44333] <= 32'b00000001010000000000001110010011;
ROM[44334] <= 32'b00000000010000111000001110010011;
ROM[44335] <= 32'b01000000011100010000001110110011;
ROM[44336] <= 32'b00000000011100000000001000110011;
ROM[44337] <= 32'b00000000001000000000000110110011;
ROM[44338] <= 32'b11110010000011100010000011101111;
ROM[44339] <= 32'b11111111110000010000000100010011;
ROM[44340] <= 32'b00000000000000010010001110000011;
ROM[44341] <= 32'b00000000011100011010000000100011;
ROM[44342] <= 32'b00000000000000000000001110010011;
ROM[44343] <= 32'b00000000011100010010000000100011;
ROM[44344] <= 32'b00000000010000010000000100010011;
ROM[44345] <= 32'b00000001010000000000001110010011;
ROM[44346] <= 32'b01000000011100011000001110110011;
ROM[44347] <= 32'b00000000000000111010000010000011;
ROM[44348] <= 32'b11111111110000010000000100010011;
ROM[44349] <= 32'b00000000000000010010001110000011;
ROM[44350] <= 32'b00000000011100100010000000100011;
ROM[44351] <= 32'b00000000010000100000000100010011;
ROM[44352] <= 32'b00000001010000000000001110010011;
ROM[44353] <= 32'b01000000011100011000001110110011;
ROM[44354] <= 32'b00000000010000111010000110000011;
ROM[44355] <= 32'b00000000100000111010001000000011;
ROM[44356] <= 32'b00000000110000111010001010000011;
ROM[44357] <= 32'b00000001000000111010001100000011;
ROM[44358] <= 32'b00000000000000001000000011100111;
ROM[44359] <= 32'b00000000000000000000001110010011;
ROM[44360] <= 32'b00000000011100010010000000100011;
ROM[44361] <= 32'b00000000010000010000000100010011;
ROM[44362] <= 32'b00010011111100000000001110010011;
ROM[44363] <= 32'b00000000011100010010000000100011;
ROM[44364] <= 32'b00000000010000010000000100010011;
ROM[44365] <= 32'b00000000000000000000001110010011;
ROM[44366] <= 32'b00000000011100010010000000100011;
ROM[44367] <= 32'b00000000010000010000000100010011;
ROM[44368] <= 32'b00000000000000101011001110110111;
ROM[44369] <= 32'b01011000110000111000001110010011;
ROM[44370] <= 32'b00000000111000111000001110110011;
ROM[44371] <= 32'b00000000011100010010000000100011;
ROM[44372] <= 32'b00000000010000010000000100010011;
ROM[44373] <= 32'b00000000001100010010000000100011;
ROM[44374] <= 32'b00000000010000010000000100010011;
ROM[44375] <= 32'b00000000010000010010000000100011;
ROM[44376] <= 32'b00000000010000010000000100010011;
ROM[44377] <= 32'b00000000010100010010000000100011;
ROM[44378] <= 32'b00000000010000010000000100010011;
ROM[44379] <= 32'b00000000011000010010000000100011;
ROM[44380] <= 32'b00000000010000010000000100010011;
ROM[44381] <= 32'b00000001010000000000001110010011;
ROM[44382] <= 32'b00000000110000111000001110010011;
ROM[44383] <= 32'b01000000011100010000001110110011;
ROM[44384] <= 32'b00000000011100000000001000110011;
ROM[44385] <= 32'b00000000001000000000000110110011;
ROM[44386] <= 32'b10100010010111110011000011101111;
ROM[44387] <= 32'b11111111110000010000000100010011;
ROM[44388] <= 32'b00000000000000010010001110000011;
ROM[44389] <= 32'b00000000011101100010000000100011;
ROM[44390] <= 32'b00000000000000000000001110010011;
ROM[44391] <= 32'b00000000011100010010000000100011;
ROM[44392] <= 32'b00000000010000010000000100010011;
ROM[44393] <= 32'b00010011111100000000001110010011;
ROM[44394] <= 32'b00000000011100010010000000100011;
ROM[44395] <= 32'b00000000010000010000000100010011;
ROM[44396] <= 32'b00001110111100000000001110010011;
ROM[44397] <= 32'b00000000011100010010000000100011;
ROM[44398] <= 32'b00000000010000010000000100010011;
ROM[44399] <= 32'b00000000000000101011001110110111;
ROM[44400] <= 32'b01100000100000111000001110010011;
ROM[44401] <= 32'b00000000111000111000001110110011;
ROM[44402] <= 32'b00000000011100010010000000100011;
ROM[44403] <= 32'b00000000010000010000000100010011;
ROM[44404] <= 32'b00000000001100010010000000100011;
ROM[44405] <= 32'b00000000010000010000000100010011;
ROM[44406] <= 32'b00000000010000010010000000100011;
ROM[44407] <= 32'b00000000010000010000000100010011;
ROM[44408] <= 32'b00000000010100010010000000100011;
ROM[44409] <= 32'b00000000010000010000000100010011;
ROM[44410] <= 32'b00000000011000010010000000100011;
ROM[44411] <= 32'b00000000010000010000000100010011;
ROM[44412] <= 32'b00000001010000000000001110010011;
ROM[44413] <= 32'b00000000110000111000001110010011;
ROM[44414] <= 32'b01000000011100010000001110110011;
ROM[44415] <= 32'b00000000011100000000001000110011;
ROM[44416] <= 32'b00000000001000000000000110110011;
ROM[44417] <= 32'b10011010100111110011000011101111;
ROM[44418] <= 32'b11111111110000010000000100010011;
ROM[44419] <= 32'b00000000000000010010001110000011;
ROM[44420] <= 32'b00000000011101100010000000100011;
ROM[44421] <= 32'b00000000000000000000001110010011;
ROM[44422] <= 32'b00000000011100010010000000100011;
ROM[44423] <= 32'b00000000010000010000000100010011;
ROM[44424] <= 32'b00000000000000000000001110010011;
ROM[44425] <= 32'b00000000011100010010000000100011;
ROM[44426] <= 32'b00000000010000010000000100010011;
ROM[44427] <= 32'b00001110111100000000001110010011;
ROM[44428] <= 32'b00000000011100010010000000100011;
ROM[44429] <= 32'b00000000010000010000000100010011;
ROM[44430] <= 32'b00000000000000101011001110110111;
ROM[44431] <= 32'b01101000010000111000001110010011;
ROM[44432] <= 32'b00000000111000111000001110110011;
ROM[44433] <= 32'b00000000011100010010000000100011;
ROM[44434] <= 32'b00000000010000010000000100010011;
ROM[44435] <= 32'b00000000001100010010000000100011;
ROM[44436] <= 32'b00000000010000010000000100010011;
ROM[44437] <= 32'b00000000010000010010000000100011;
ROM[44438] <= 32'b00000000010000010000000100010011;
ROM[44439] <= 32'b00000000010100010010000000100011;
ROM[44440] <= 32'b00000000010000010000000100010011;
ROM[44441] <= 32'b00000000011000010010000000100011;
ROM[44442] <= 32'b00000000010000010000000100010011;
ROM[44443] <= 32'b00000001010000000000001110010011;
ROM[44444] <= 32'b00000000110000111000001110010011;
ROM[44445] <= 32'b01000000011100010000001110110011;
ROM[44446] <= 32'b00000000011100000000001000110011;
ROM[44447] <= 32'b00000000001000000000000110110011;
ROM[44448] <= 32'b10110100100111110011000011101111;
ROM[44449] <= 32'b11111111110000010000000100010011;
ROM[44450] <= 32'b00000000000000010010001110000011;
ROM[44451] <= 32'b00000000011101100010000000100011;
ROM[44452] <= 32'b00010011111100000000001110010011;
ROM[44453] <= 32'b00000000011100010010000000100011;
ROM[44454] <= 32'b00000000010000010000000100010011;
ROM[44455] <= 32'b00000000000000000000001110010011;
ROM[44456] <= 32'b00000000011100010010000000100011;
ROM[44457] <= 32'b00000000010000010000000100010011;
ROM[44458] <= 32'b00001110111100000000001110010011;
ROM[44459] <= 32'b00000000011100010010000000100011;
ROM[44460] <= 32'b00000000010000010000000100010011;
ROM[44461] <= 32'b00000000000000101011001110110111;
ROM[44462] <= 32'b01110000000000111000001110010011;
ROM[44463] <= 32'b00000000111000111000001110110011;
ROM[44464] <= 32'b00000000011100010010000000100011;
ROM[44465] <= 32'b00000000010000010000000100010011;
ROM[44466] <= 32'b00000000001100010010000000100011;
ROM[44467] <= 32'b00000000010000010000000100010011;
ROM[44468] <= 32'b00000000010000010010000000100011;
ROM[44469] <= 32'b00000000010000010000000100010011;
ROM[44470] <= 32'b00000000010100010010000000100011;
ROM[44471] <= 32'b00000000010000010000000100010011;
ROM[44472] <= 32'b00000000011000010010000000100011;
ROM[44473] <= 32'b00000000010000010000000100010011;
ROM[44474] <= 32'b00000001010000000000001110010011;
ROM[44475] <= 32'b00000000110000111000001110010011;
ROM[44476] <= 32'b01000000011100010000001110110011;
ROM[44477] <= 32'b00000000011100000000001000110011;
ROM[44478] <= 32'b00000000001000000000000110110011;
ROM[44479] <= 32'b10101100110111110011000011101111;
ROM[44480] <= 32'b11111111110000010000000100010011;
ROM[44481] <= 32'b00000000000000010010001110000011;
ROM[44482] <= 32'b00000000011101100010000000100011;
ROM[44483] <= 32'b00000011001000000000001110010011;
ROM[44484] <= 32'b00000000011100010010000000100011;
ROM[44485] <= 32'b00000000010000010000000100010011;
ROM[44486] <= 32'b00000110010000000000001110010011;
ROM[44487] <= 32'b00000000011100010010000000100011;
ROM[44488] <= 32'b00000000010000010000000100010011;
ROM[44489] <= 32'b00000011001000000000001110010011;
ROM[44490] <= 32'b00000000011100010010000000100011;
ROM[44491] <= 32'b00000000010000010000000100010011;
ROM[44492] <= 32'b00000000000000101011001110110111;
ROM[44493] <= 32'b01110111110000111000001110010011;
ROM[44494] <= 32'b00000000111000111000001110110011;
ROM[44495] <= 32'b00000000011100010010000000100011;
ROM[44496] <= 32'b00000000010000010000000100010011;
ROM[44497] <= 32'b00000000001100010010000000100011;
ROM[44498] <= 32'b00000000010000010000000100010011;
ROM[44499] <= 32'b00000000010000010010000000100011;
ROM[44500] <= 32'b00000000010000010000000100010011;
ROM[44501] <= 32'b00000000010100010010000000100011;
ROM[44502] <= 32'b00000000010000010000000100010011;
ROM[44503] <= 32'b00000000011000010010000000100011;
ROM[44504] <= 32'b00000000010000010000000100010011;
ROM[44505] <= 32'b00000001010000000000001110010011;
ROM[44506] <= 32'b00000000110000111000001110010011;
ROM[44507] <= 32'b01000000011100010000001110110011;
ROM[44508] <= 32'b00000000011100000000001000110011;
ROM[44509] <= 32'b00000000001000000000000110110011;
ROM[44510] <= 32'b10000011010111110011000011101111;
ROM[44511] <= 32'b11111111110000010000000100010011;
ROM[44512] <= 32'b00000000000000010010001110000011;
ROM[44513] <= 32'b00000000011101100010000000100011;
ROM[44514] <= 32'b00000011001000000000001110010011;
ROM[44515] <= 32'b00000000011100010010000000100011;
ROM[44516] <= 32'b00000000010000010000000100010011;
ROM[44517] <= 32'b00000110010000000000001110010011;
ROM[44518] <= 32'b00000000011100010010000000100011;
ROM[44519] <= 32'b00000000010000010000000100010011;
ROM[44520] <= 32'b00000110010000000000001110010011;
ROM[44521] <= 32'b00000000011100010010000000100011;
ROM[44522] <= 32'b00000000010000010000000100010011;
ROM[44523] <= 32'b00000000000000101011001110110111;
ROM[44524] <= 32'b01111111100000111000001110010011;
ROM[44525] <= 32'b00000000111000111000001110110011;
ROM[44526] <= 32'b00000000011100010010000000100011;
ROM[44527] <= 32'b00000000010000010000000100010011;
ROM[44528] <= 32'b00000000001100010010000000100011;
ROM[44529] <= 32'b00000000010000010000000100010011;
ROM[44530] <= 32'b00000000010000010010000000100011;
ROM[44531] <= 32'b00000000010000010000000100010011;
ROM[44532] <= 32'b00000000010100010010000000100011;
ROM[44533] <= 32'b00000000010000010000000100010011;
ROM[44534] <= 32'b00000000011000010010000000100011;
ROM[44535] <= 32'b00000000010000010000000100010011;
ROM[44536] <= 32'b00000001010000000000001110010011;
ROM[44537] <= 32'b00000000110000111000001110010011;
ROM[44538] <= 32'b01000000011100010000001110110011;
ROM[44539] <= 32'b00000000011100000000001000110011;
ROM[44540] <= 32'b00000000001000000000000110110011;
ROM[44541] <= 32'b11111011100011110011000011101111;
ROM[44542] <= 32'b11111111110000010000000100010011;
ROM[44543] <= 32'b00000000000000010010001110000011;
ROM[44544] <= 32'b00000000011101100010000000100011;
ROM[44545] <= 32'b00000011001000000000001110010011;
ROM[44546] <= 32'b00000000011100010010000000100011;
ROM[44547] <= 32'b00000000010000010000000100010011;
ROM[44548] <= 32'b00000110010000000000001110010011;
ROM[44549] <= 32'b00000000011100010010000000100011;
ROM[44550] <= 32'b00000000010000010000000100010011;
ROM[44551] <= 32'b00000011001000000000001110010011;
ROM[44552] <= 32'b00000000011100010010000000100011;
ROM[44553] <= 32'b00000000010000010000000100010011;
ROM[44554] <= 32'b00000000000000101100001110110111;
ROM[44555] <= 32'b10000111010000111000001110010011;
ROM[44556] <= 32'b00000000111000111000001110110011;
ROM[44557] <= 32'b00000000011100010010000000100011;
ROM[44558] <= 32'b00000000010000010000000100010011;
ROM[44559] <= 32'b00000000001100010010000000100011;
ROM[44560] <= 32'b00000000010000010000000100010011;
ROM[44561] <= 32'b00000000010000010010000000100011;
ROM[44562] <= 32'b00000000010000010000000100010011;
ROM[44563] <= 32'b00000000010100010010000000100011;
ROM[44564] <= 32'b00000000010000010000000100010011;
ROM[44565] <= 32'b00000000011000010010000000100011;
ROM[44566] <= 32'b00000000010000010000000100010011;
ROM[44567] <= 32'b00000001010000000000001110010011;
ROM[44568] <= 32'b00000000110000111000001110010011;
ROM[44569] <= 32'b01000000011100010000001110110011;
ROM[44570] <= 32'b00000000011100000000001000110011;
ROM[44571] <= 32'b00000000001000000000000110110011;
ROM[44572] <= 32'b10010101100111110011000011101111;
ROM[44573] <= 32'b11111111110000010000000100010011;
ROM[44574] <= 32'b00000000000000010010001110000011;
ROM[44575] <= 32'b00000000011101100010000000100011;
ROM[44576] <= 32'b00000011001000000000001110010011;
ROM[44577] <= 32'b00000000011100010010000000100011;
ROM[44578] <= 32'b00000000010000010000000100010011;
ROM[44579] <= 32'b00000110010000000000001110010011;
ROM[44580] <= 32'b00000000011100010010000000100011;
ROM[44581] <= 32'b00000000010000010000000100010011;
ROM[44582] <= 32'b00000110010000000000001110010011;
ROM[44583] <= 32'b00000000011100010010000000100011;
ROM[44584] <= 32'b00000000010000010000000100010011;
ROM[44585] <= 32'b00000000000000101100001110110111;
ROM[44586] <= 32'b10001111000000111000001110010011;
ROM[44587] <= 32'b00000000111000111000001110110011;
ROM[44588] <= 32'b00000000011100010010000000100011;
ROM[44589] <= 32'b00000000010000010000000100010011;
ROM[44590] <= 32'b00000000001100010010000000100011;
ROM[44591] <= 32'b00000000010000010000000100010011;
ROM[44592] <= 32'b00000000010000010010000000100011;
ROM[44593] <= 32'b00000000010000010000000100010011;
ROM[44594] <= 32'b00000000010100010010000000100011;
ROM[44595] <= 32'b00000000010000010000000100010011;
ROM[44596] <= 32'b00000000011000010010000000100011;
ROM[44597] <= 32'b00000000010000010000000100010011;
ROM[44598] <= 32'b00000001010000000000001110010011;
ROM[44599] <= 32'b00000000110000111000001110010011;
ROM[44600] <= 32'b01000000011100010000001110110011;
ROM[44601] <= 32'b00000000011100000000001000110011;
ROM[44602] <= 32'b00000000001000000000000110110011;
ROM[44603] <= 32'b10001101110111110011000011101111;
ROM[44604] <= 32'b11111111110000010000000100010011;
ROM[44605] <= 32'b00000000000000010010001110000011;
ROM[44606] <= 32'b00000000011101100010000000100011;
ROM[44607] <= 32'b00000000000000000000001110010011;
ROM[44608] <= 32'b00000000011100010010000000100011;
ROM[44609] <= 32'b00000000010000010000000100010011;
ROM[44610] <= 32'b00000000000000000000001110010011;
ROM[44611] <= 32'b00000000011100010010000000100011;
ROM[44612] <= 32'b00000000010000010000000100010011;
ROM[44613] <= 32'b00000011001000000000001110010011;
ROM[44614] <= 32'b00000000011100010010000000100011;
ROM[44615] <= 32'b00000000010000010000000100010011;
ROM[44616] <= 32'b00000011001000000000001110010011;
ROM[44617] <= 32'b00000000011100010010000000100011;
ROM[44618] <= 32'b00000000010000010000000100010011;
ROM[44619] <= 32'b00000000000000101100001110110111;
ROM[44620] <= 32'b10010111100000111000001110010011;
ROM[44621] <= 32'b00000000111000111000001110110011;
ROM[44622] <= 32'b00000000011100010010000000100011;
ROM[44623] <= 32'b00000000010000010000000100010011;
ROM[44624] <= 32'b00000000001100010010000000100011;
ROM[44625] <= 32'b00000000010000010000000100010011;
ROM[44626] <= 32'b00000000010000010010000000100011;
ROM[44627] <= 32'b00000000010000010000000100010011;
ROM[44628] <= 32'b00000000010100010010000000100011;
ROM[44629] <= 32'b00000000010000010000000100010011;
ROM[44630] <= 32'b00000000011000010010000000100011;
ROM[44631] <= 32'b00000000010000010000000100010011;
ROM[44632] <= 32'b00000001010000000000001110010011;
ROM[44633] <= 32'b00000001000000111000001110010011;
ROM[44634] <= 32'b01000000011100010000001110110011;
ROM[44635] <= 32'b00000000011100000000001000110011;
ROM[44636] <= 32'b00000000001000000000000110110011;
ROM[44637] <= 32'b10111101010111110010000011101111;
ROM[44638] <= 32'b11111111110000010000000100010011;
ROM[44639] <= 32'b00000000000000010010001110000011;
ROM[44640] <= 32'b00000000011101100010000000100011;
ROM[44641] <= 32'b00010011111100000000001110010011;
ROM[44642] <= 32'b00000000011100010010000000100011;
ROM[44643] <= 32'b00000000010000010000000100010011;
ROM[44644] <= 32'b00001110111100000000001110010011;
ROM[44645] <= 32'b00000000011100010010000000100011;
ROM[44646] <= 32'b00000000010000010000000100010011;
ROM[44647] <= 32'b00000110010000000000001110010011;
ROM[44648] <= 32'b00000000011100010010000000100011;
ROM[44649] <= 32'b00000000010000010000000100010011;
ROM[44650] <= 32'b00000110010000000000001110010011;
ROM[44651] <= 32'b00000000011100010010000000100011;
ROM[44652] <= 32'b00000000010000010000000100010011;
ROM[44653] <= 32'b00000000000000101100001110110111;
ROM[44654] <= 32'b10100000000000111000001110010011;
ROM[44655] <= 32'b00000000111000111000001110110011;
ROM[44656] <= 32'b00000000011100010010000000100011;
ROM[44657] <= 32'b00000000010000010000000100010011;
ROM[44658] <= 32'b00000000001100010010000000100011;
ROM[44659] <= 32'b00000000010000010000000100010011;
ROM[44660] <= 32'b00000000010000010010000000100011;
ROM[44661] <= 32'b00000000010000010000000100010011;
ROM[44662] <= 32'b00000000010100010010000000100011;
ROM[44663] <= 32'b00000000010000010000000100010011;
ROM[44664] <= 32'b00000000011000010010000000100011;
ROM[44665] <= 32'b00000000010000010000000100010011;
ROM[44666] <= 32'b00000001010000000000001110010011;
ROM[44667] <= 32'b00000001000000111000001110010011;
ROM[44668] <= 32'b01000000011100010000001110110011;
ROM[44669] <= 32'b00000000011100000000001000110011;
ROM[44670] <= 32'b00000000001000000000000110110011;
ROM[44671] <= 32'b10110100110111110010000011101111;
ROM[44672] <= 32'b11111111110000010000000100010011;
ROM[44673] <= 32'b00000000000000010010001110000011;
ROM[44674] <= 32'b00000000011101100010000000100011;
ROM[44675] <= 32'b00000000001000000000001110010011;
ROM[44676] <= 32'b00000000011100010010000000100011;
ROM[44677] <= 32'b00000000010000010000000100010011;
ROM[44678] <= 32'b00000000001000000000001110010011;
ROM[44679] <= 32'b00000000011100010010000000100011;
ROM[44680] <= 32'b00000000010000010000000100010011;
ROM[44681] <= 32'b00000000010000000000001110010011;
ROM[44682] <= 32'b00000000011100010010000000100011;
ROM[44683] <= 32'b00000000010000010000000100010011;
ROM[44684] <= 32'b00000000010000000000001110010011;
ROM[44685] <= 32'b00000000011100010010000000100011;
ROM[44686] <= 32'b00000000010000010000000100010011;
ROM[44687] <= 32'b00000000000000101100001110110111;
ROM[44688] <= 32'b10101000100000111000001110010011;
ROM[44689] <= 32'b00000000111000111000001110110011;
ROM[44690] <= 32'b00000000011100010010000000100011;
ROM[44691] <= 32'b00000000010000010000000100010011;
ROM[44692] <= 32'b00000000001100010010000000100011;
ROM[44693] <= 32'b00000000010000010000000100010011;
ROM[44694] <= 32'b00000000010000010010000000100011;
ROM[44695] <= 32'b00000000010000010000000100010011;
ROM[44696] <= 32'b00000000010100010010000000100011;
ROM[44697] <= 32'b00000000010000010000000100010011;
ROM[44698] <= 32'b00000000011000010010000000100011;
ROM[44699] <= 32'b00000000010000010000000100010011;
ROM[44700] <= 32'b00000001010000000000001110010011;
ROM[44701] <= 32'b00000001000000111000001110010011;
ROM[44702] <= 32'b01000000011100010000001110110011;
ROM[44703] <= 32'b00000000011100000000001000110011;
ROM[44704] <= 32'b00000000001000000000000110110011;
ROM[44705] <= 32'b10010110000111110011000011101111;
ROM[44706] <= 32'b11111111110000010000000100010011;
ROM[44707] <= 32'b00000000000000010010001110000011;
ROM[44708] <= 32'b00000000011101100010000000100011;
ROM[44709] <= 32'b00000000000000000000001110010011;
ROM[44710] <= 32'b00000000011100010010000000100011;
ROM[44711] <= 32'b00000000010000010000000100010011;
ROM[44712] <= 32'b00000001010000000000001110010011;
ROM[44713] <= 32'b01000000011100011000001110110011;
ROM[44714] <= 32'b00000000000000111010000010000011;
ROM[44715] <= 32'b11111111110000010000000100010011;
ROM[44716] <= 32'b00000000000000010010001110000011;
ROM[44717] <= 32'b00000000011100100010000000100011;
ROM[44718] <= 32'b00000000010000100000000100010011;
ROM[44719] <= 32'b00000001010000000000001110010011;
ROM[44720] <= 32'b01000000011100011000001110110011;
ROM[44721] <= 32'b00000000010000111010000110000011;
ROM[44722] <= 32'b00000000100000111010001000000011;
ROM[44723] <= 32'b00000000110000111010001010000011;
ROM[44724] <= 32'b00000001000000111010001100000011;
ROM[44725] <= 32'b00000000000000001000000011100111;
ROM[44726] <= 32'b00000000001100000000001110010011;
ROM[44727] <= 32'b00000000011100010010000000100011;
ROM[44728] <= 32'b00000000010000010000000100010011;
ROM[44729] <= 32'b00000000000000101100001110110111;
ROM[44730] <= 32'b10110011000000111000001110010011;
ROM[44731] <= 32'b00000000111000111000001110110011;
ROM[44732] <= 32'b00000000011100010010000000100011;
ROM[44733] <= 32'b00000000010000010000000100010011;
ROM[44734] <= 32'b00000000001100010010000000100011;
ROM[44735] <= 32'b00000000010000010000000100010011;
ROM[44736] <= 32'b00000000010000010010000000100011;
ROM[44737] <= 32'b00000000010000010000000100010011;
ROM[44738] <= 32'b00000000010100010010000000100011;
ROM[44739] <= 32'b00000000010000010000000100010011;
ROM[44740] <= 32'b00000000011000010010000000100011;
ROM[44741] <= 32'b00000000010000010000000100010011;
ROM[44742] <= 32'b00000001010000000000001110010011;
ROM[44743] <= 32'b00000000010000111000001110010011;
ROM[44744] <= 32'b01000000011100010000001110110011;
ROM[44745] <= 32'b00000000011100000000001000110011;
ROM[44746] <= 32'b00000000001000000000000110110011;
ROM[44747] <= 32'b11000001000111111101000011101111;
ROM[44748] <= 32'b00000100010100000000001110010011;
ROM[44749] <= 32'b00000000011100010010000000100011;
ROM[44750] <= 32'b00000000010000010000000100010011;
ROM[44751] <= 32'b00000000000000101100001110110111;
ROM[44752] <= 32'b10111000100000111000001110010011;
ROM[44753] <= 32'b00000000111000111000001110110011;
ROM[44754] <= 32'b00000000011100010010000000100011;
ROM[44755] <= 32'b00000000010000010000000100010011;
ROM[44756] <= 32'b00000000001100010010000000100011;
ROM[44757] <= 32'b00000000010000010000000100010011;
ROM[44758] <= 32'b00000000010000010010000000100011;
ROM[44759] <= 32'b00000000010000010000000100010011;
ROM[44760] <= 32'b00000000010100010010000000100011;
ROM[44761] <= 32'b00000000010000010000000100010011;
ROM[44762] <= 32'b00000000011000010010000000100011;
ROM[44763] <= 32'b00000000010000010000000100010011;
ROM[44764] <= 32'b00000001010000000000001110010011;
ROM[44765] <= 32'b00000000100000111000001110010011;
ROM[44766] <= 32'b01000000011100010000001110110011;
ROM[44767] <= 32'b00000000011100000000001000110011;
ROM[44768] <= 32'b00000000001000000000000110110011;
ROM[44769] <= 32'b10000010100011111110000011101111;
ROM[44770] <= 32'b00000111001000000000001110010011;
ROM[44771] <= 32'b00000000011100010010000000100011;
ROM[44772] <= 32'b00000000010000010000000100010011;
ROM[44773] <= 32'b00000000000000101100001110110111;
ROM[44774] <= 32'b10111110000000111000001110010011;
ROM[44775] <= 32'b00000000111000111000001110110011;
ROM[44776] <= 32'b00000000011100010010000000100011;
ROM[44777] <= 32'b00000000010000010000000100010011;
ROM[44778] <= 32'b00000000001100010010000000100011;
ROM[44779] <= 32'b00000000010000010000000100010011;
ROM[44780] <= 32'b00000000010000010010000000100011;
ROM[44781] <= 32'b00000000010000010000000100010011;
ROM[44782] <= 32'b00000000010100010010000000100011;
ROM[44783] <= 32'b00000000010000010000000100010011;
ROM[44784] <= 32'b00000000011000010010000000100011;
ROM[44785] <= 32'b00000000010000010000000100010011;
ROM[44786] <= 32'b00000001010000000000001110010011;
ROM[44787] <= 32'b00000000100000111000001110010011;
ROM[44788] <= 32'b01000000011100010000001110110011;
ROM[44789] <= 32'b00000000011100000000001000110011;
ROM[44790] <= 32'b00000000001000000000000110110011;
ROM[44791] <= 32'b11111101000111111101000011101111;
ROM[44792] <= 32'b00000111001000000000001110010011;
ROM[44793] <= 32'b00000000011100010010000000100011;
ROM[44794] <= 32'b00000000010000010000000100010011;
ROM[44795] <= 32'b00000000000000101100001110110111;
ROM[44796] <= 32'b11000011100000111000001110010011;
ROM[44797] <= 32'b00000000111000111000001110110011;
ROM[44798] <= 32'b00000000011100010010000000100011;
ROM[44799] <= 32'b00000000010000010000000100010011;
ROM[44800] <= 32'b00000000001100010010000000100011;
ROM[44801] <= 32'b00000000010000010000000100010011;
ROM[44802] <= 32'b00000000010000010010000000100011;
ROM[44803] <= 32'b00000000010000010000000100010011;
ROM[44804] <= 32'b00000000010100010010000000100011;
ROM[44805] <= 32'b00000000010000010000000100010011;
ROM[44806] <= 32'b00000000011000010010000000100011;
ROM[44807] <= 32'b00000000010000010000000100010011;
ROM[44808] <= 32'b00000001010000000000001110010011;
ROM[44809] <= 32'b00000000100000111000001110010011;
ROM[44810] <= 32'b01000000011100010000001110110011;
ROM[44811] <= 32'b00000000011100000000001000110011;
ROM[44812] <= 32'b00000000001000000000000110110011;
ROM[44813] <= 32'b11110111100111111101000011101111;
ROM[44814] <= 32'b00000000000000101100001110110111;
ROM[44815] <= 32'b11001000010000111000001110010011;
ROM[44816] <= 32'b00000000111000111000001110110011;
ROM[44817] <= 32'b00000000011100010010000000100011;
ROM[44818] <= 32'b00000000010000010000000100010011;
ROM[44819] <= 32'b00000000001100010010000000100011;
ROM[44820] <= 32'b00000000010000010000000100010011;
ROM[44821] <= 32'b00000000010000010010000000100011;
ROM[44822] <= 32'b00000000010000010000000100010011;
ROM[44823] <= 32'b00000000010100010010000000100011;
ROM[44824] <= 32'b00000000010000010000000100010011;
ROM[44825] <= 32'b00000000011000010010000000100011;
ROM[44826] <= 32'b00000000010000010000000100010011;
ROM[44827] <= 32'b00000001010000000000001110010011;
ROM[44828] <= 32'b00000000010000111000001110010011;
ROM[44829] <= 32'b01000000011100010000001110110011;
ROM[44830] <= 32'b00000000011100000000001000110011;
ROM[44831] <= 32'b00000000001000000000000110110011;
ROM[44832] <= 32'b10101110100011101011000011101111;
ROM[44833] <= 32'b11111111110000010000000100010011;
ROM[44834] <= 32'b00000000000000010010001110000011;
ROM[44835] <= 32'b00000000011101100010000000100011;
ROM[44836] <= 32'b00000000000000100010001110000011;
ROM[44837] <= 32'b00000000011100010010000000100011;
ROM[44838] <= 32'b00000000010000010000000100010011;
ROM[44839] <= 32'b00000000000000101100001110110111;
ROM[44840] <= 32'b11001110100000111000001110010011;
ROM[44841] <= 32'b00000000111000111000001110110011;
ROM[44842] <= 32'b00000000011100010010000000100011;
ROM[44843] <= 32'b00000000010000010000000100010011;
ROM[44844] <= 32'b00000000001100010010000000100011;
ROM[44845] <= 32'b00000000010000010000000100010011;
ROM[44846] <= 32'b00000000010000010010000000100011;
ROM[44847] <= 32'b00000000010000010000000100010011;
ROM[44848] <= 32'b00000000010100010010000000100011;
ROM[44849] <= 32'b00000000010000010000000100010011;
ROM[44850] <= 32'b00000000011000010010000000100011;
ROM[44851] <= 32'b00000000010000010000000100010011;
ROM[44852] <= 32'b00000001010000000000001110010011;
ROM[44853] <= 32'b00000000010000111000001110010011;
ROM[44854] <= 32'b01000000011100010000001110110011;
ROM[44855] <= 32'b00000000011100000000001000110011;
ROM[44856] <= 32'b00000000001000000000000110110011;
ROM[44857] <= 32'b10101000010011101011000011101111;
ROM[44858] <= 32'b11111111110000010000000100010011;
ROM[44859] <= 32'b00000000000000010010001110000011;
ROM[44860] <= 32'b00000000011101100010000000100011;
ROM[44861] <= 32'b00000000000000101100001110110111;
ROM[44862] <= 32'b11010100000000111000001110010011;
ROM[44863] <= 32'b00000000111000111000001110110011;
ROM[44864] <= 32'b00000000011100010010000000100011;
ROM[44865] <= 32'b00000000010000010000000100010011;
ROM[44866] <= 32'b00000000001100010010000000100011;
ROM[44867] <= 32'b00000000010000010000000100010011;
ROM[44868] <= 32'b00000000010000010010000000100011;
ROM[44869] <= 32'b00000000010000010000000100010011;
ROM[44870] <= 32'b00000000010100010010000000100011;
ROM[44871] <= 32'b00000000010000010000000100010011;
ROM[44872] <= 32'b00000000011000010010000000100011;
ROM[44873] <= 32'b00000000010000010000000100010011;
ROM[44874] <= 32'b00000001010000000000001110010011;
ROM[44875] <= 32'b00000000000000111000001110010011;
ROM[44876] <= 32'b01000000011100010000001110110011;
ROM[44877] <= 32'b00000000011100000000001000110011;
ROM[44878] <= 32'b00000000001000000000000110110011;
ROM[44879] <= 32'b10101110110011111111000011101111;
ROM[44880] <= 32'b11111111110000010000000100010011;
ROM[44881] <= 32'b00000000000000010010001110000011;
ROM[44882] <= 32'b00000000011101100010000000100011;
ROM[44883] <= 32'b00000000000000000000001110010011;
ROM[44884] <= 32'b00000000011100010010000000100011;
ROM[44885] <= 32'b00000000010000010000000100010011;
ROM[44886] <= 32'b00000001010000000000001110010011;
ROM[44887] <= 32'b01000000011100011000001110110011;
ROM[44888] <= 32'b00000000000000111010000010000011;
ROM[44889] <= 32'b11111111110000010000000100010011;
ROM[44890] <= 32'b00000000000000010010001110000011;
ROM[44891] <= 32'b00000000011100100010000000100011;
ROM[44892] <= 32'b00000000010000100000000100010011;
ROM[44893] <= 32'b00000001010000000000001110010011;
ROM[44894] <= 32'b01000000011100011000001110110011;
ROM[44895] <= 32'b00000000010000111010000110000011;
ROM[44896] <= 32'b00000000100000111010001000000011;
ROM[44897] <= 32'b00000000110000111010001010000011;
ROM[44898] <= 32'b00000001000000111010001100000011;
ROM[44899] <= 32'b00000000000000001000000011100111;
ROM[44900] <= 32'b00000000000000111000000010010011;
        end
    assign address = addr[16:2];
    assign Inst = ROM[address];
        
endmodule