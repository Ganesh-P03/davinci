module ROM ( //Instruction Memory
    input [16:0] addr,
    input clock,
    output [31:0] Inst
    );
    wire [14:0] address;
    
    (* ram_style="block" *)
    reg [31:0] ROM[32767:0];

    initial
        begin
    ROM[0] <= 32'b00000000000000000010011100110111;
ROM[1] <= 32'b01011000000001110000011100010011;
ROM[2] <= 32'b00000000000000100010011010110111;
ROM[3] <= 32'b01011000000001101000011010010011;
ROM[4] <= 32'b00000100000001101010000000100011;
ROM[5] <= 32'b00000100000001101010001000100011;
ROM[6] <= 32'b00000100000001101010010000100011;
ROM[7] <= 32'b00000100000001101010011000100011;
ROM[8] <= 32'b00000100000001101010100000100011;
ROM[9] <= 32'b00000100000001101010101000100011;
ROM[10] <= 32'b00000100000001101010110000100011;
ROM[11] <= 32'b00000100000001101010111000100011;
ROM[12] <= 32'b00000110000001101010000000100011;
ROM[13] <= 32'b00000110000001101010001000100011;
ROM[14] <= 32'b00000110000001101010010000100011;
ROM[15] <= 32'b00000110000001101010011000100011;
ROM[16] <= 32'b00000110000001101010100000100011;
ROM[17] <= 32'b00000110000001101010101000100011;
ROM[18] <= 32'b00000110000001101010110000100011;
ROM[19] <= 32'b00000110000001101010111000100011;
ROM[20] <= 32'b00001000000001101010000000100011;
ROM[21] <= 32'b00001000000001101010001000100011;
ROM[22] <= 32'b00001000000001101010010000100011;
ROM[23] <= 32'b00001000000001101010011000100011;
ROM[24] <= 32'b00001000000001101010100000100011;
ROM[25] <= 32'b00001000000001101010101000100011;
ROM[26] <= 32'b00001000000001101010110000100011;
ROM[27] <= 32'b00001000000001101010111000100011;
ROM[28] <= 32'b00001010000001101010000000100011;
ROM[29] <= 32'b00001010000001101010001000100011;
ROM[30] <= 32'b00001010000001101010010000100011;
ROM[31] <= 32'b00001010000001101010011000100011;
ROM[32] <= 32'b00001010000001101010100000100011;
ROM[33] <= 32'b00001010000001101010101000100011;
ROM[34] <= 32'b00001010000001101010110000100011;
ROM[35] <= 32'b00001010000001101010111000100011;
ROM[36] <= 32'b00001100000001101010000000100011;
ROM[37] <= 32'b00001100000001101010001000100011;
ROM[38] <= 32'b00001100000001101010010000100011;
ROM[39] <= 32'b00001100000001101010011000100011;
ROM[40] <= 32'b00001100000001101010100000100011;
ROM[41] <= 32'b00001100000001101010101000100011;
ROM[42] <= 32'b00001100000001101010110000100011;
ROM[43] <= 32'b00001100000001101010111000100011;
ROM[44] <= 32'b00001110000001101010000000100011;
ROM[45] <= 32'b00001110000001101010001000100011;
ROM[46] <= 32'b00001110000001101010010000100011;
ROM[47] <= 32'b00001110000001101010011000100011;
ROM[48] <= 32'b00001110000001101010100000100011;
ROM[49] <= 32'b00001110000001101010101000100011;
ROM[50] <= 32'b00001110000001101010110000100011;
ROM[51] <= 32'b00001110000001101010111000100011;
ROM[52] <= 32'b00010000000001101010000000100011;
ROM[53] <= 32'b00010000000001101010001000100011;
ROM[54] <= 32'b00010000000001101010010000100011;
ROM[55] <= 32'b00010000000001101010011000100011;
ROM[56] <= 32'b00010000000001101010100000100011;
ROM[57] <= 32'b00010000000001101010101000100011;
ROM[58] <= 32'b00010000000001101010110000100011;
ROM[59] <= 32'b00010000000001101010111000100011;
ROM[60] <= 32'b00010010000001101010000000100011;
ROM[61] <= 32'b00010010000001101010001000100011;
ROM[62] <= 32'b00010010000001101010010000100011;
ROM[63] <= 32'b00010010000001101010011000100011;
ROM[64] <= 32'b00010010000001101010100000100011;
ROM[65] <= 32'b00010010000001101010101000100011;
ROM[66] <= 32'b00010010000001101010110000100011;
ROM[67] <= 32'b00010010000001101010111000100011;
ROM[68] <= 32'b00010100000001101010000000100011;
ROM[69] <= 32'b00010100000001101010001000100011;
ROM[70] <= 32'b00010100000001101010010000100011;
ROM[71] <= 32'b00010100000001101010011000100011;
ROM[72] <= 32'b00010100000001101010100000100011;
ROM[73] <= 32'b00010100000001101010101000100011;
ROM[74] <= 32'b00010100000001101010110000100011;
ROM[75] <= 32'b00010100000001101010111000100011;
ROM[76] <= 32'b00010110000001101010000000100011;
ROM[77] <= 32'b00010110000001101010001000100011;
ROM[78] <= 32'b00010110000001101010010000100011;
ROM[79] <= 32'b00010110000001101010011000100011;
ROM[80] <= 32'b00010110000001101010100000100011;
ROM[81] <= 32'b00010110000001101010101000100011;
ROM[82] <= 32'b00010110000001101010110000100011;
ROM[83] <= 32'b00010110000001101010111000100011;
ROM[84] <= 32'b00011000000001101010000000100011;
ROM[85] <= 32'b00011000000001101010001000100011;
ROM[86] <= 32'b00011000000001101010010000100011;
ROM[87] <= 32'b00011000000001101010011000100011;
ROM[88] <= 32'b00011000000001101010100000100011;
ROM[89] <= 32'b00011000000001101010101000100011;
ROM[90] <= 32'b00011000000001101010110000100011;
ROM[91] <= 32'b00011000000001101010111000100011;
ROM[92] <= 32'b00011010000001101010000000100011;
ROM[93] <= 32'b00011010000001101010001000100011;
ROM[94] <= 32'b00011010000001101010010000100011;
ROM[95] <= 32'b00011010000001101010011000100011;
ROM[96] <= 32'b00011010000001101010100000100011;
ROM[97] <= 32'b00011010000001101010101000100011;
ROM[98] <= 32'b00011010000001101010110000100011;
ROM[99] <= 32'b00011010000001101010111000100011;
ROM[100] <= 32'b00011100000001101010000000100011;
ROM[101] <= 32'b00011100000001101010001000100011;
ROM[102] <= 32'b00011100000001101010010000100011;
ROM[103] <= 32'b00011100000001101010011000100011;
ROM[104] <= 32'b00011100000001101010100000100011;
ROM[105] <= 32'b00011100000001101010101000100011;
ROM[106] <= 32'b00011100000001101010110000100011;
ROM[107] <= 32'b00011100000001101010111000100011;
ROM[108] <= 32'b00011110000001101010000000100011;
ROM[109] <= 32'b00011110000001101010001000100011;
ROM[110] <= 32'b00011110000001101010010000100011;
ROM[111] <= 32'b00011110000001101010011000100011;
ROM[112] <= 32'b00011110000001101010100000100011;
ROM[113] <= 32'b00011110000001101010101000100011;
ROM[114] <= 32'b00011110000001101010110000100011;
ROM[115] <= 32'b00011110000001101010111000100011;
ROM[116] <= 32'b00100000000001101010000000100011;
ROM[117] <= 32'b00100000000001101010001000100011;
ROM[118] <= 32'b00100000000001101010010000100011;
ROM[119] <= 32'b00100000000001101010011000100011;
ROM[120] <= 32'b00100000000001101010100000100011;
ROM[121] <= 32'b00100000000001101010101000100011;
ROM[122] <= 32'b00100000000001101010110000100011;
ROM[123] <= 32'b00100000000001101010111000100011;
ROM[124] <= 32'b00100010000001101010000000100011;
ROM[125] <= 32'b00100010000001101010001000100011;
ROM[126] <= 32'b00100010000001101010010000100011;
ROM[127] <= 32'b00100010000001101010011000100011;
ROM[128] <= 32'b00100010000001101010100000100011;
ROM[129] <= 32'b00100010000001101010101000100011;
ROM[130] <= 32'b00100010000001101010110000100011;
ROM[131] <= 32'b00100010000001101010111000100011;
ROM[132] <= 32'b00100100000001101010000000100011;
ROM[133] <= 32'b00100100000001101010001000100011;
ROM[134] <= 32'b00100100000001101010010000100011;
ROM[135] <= 32'b00100100000001101010011000100011;
ROM[136] <= 32'b00100100000001101010100000100011;
ROM[137] <= 32'b00100100000001101010101000100011;
ROM[138] <= 32'b00100100000001101010110000100011;
ROM[139] <= 32'b00100100000001101010111000100011;
ROM[140] <= 32'b00100110000001101010000000100011;
ROM[141] <= 32'b00100110000001101010001000100011;
ROM[142] <= 32'b00100110000001101010010000100011;
ROM[143] <= 32'b00100110000001101010011000100011;
ROM[144] <= 32'b00100110000001101010100000100011;
ROM[145] <= 32'b00100110000001101010101000100011;
ROM[146] <= 32'b00100110000001101010110000100011;
ROM[147] <= 32'b00100110000001101010111000100011;
ROM[148] <= 32'b00101000000001101010000000100011;
ROM[149] <= 32'b00101000000001101010001000100011;
ROM[150] <= 32'b00101000000001101010010000100011;
ROM[151] <= 32'b00101000000001101010011000100011;
ROM[152] <= 32'b00101000000001101010100000100011;
ROM[153] <= 32'b00101000000001101010101000100011;
ROM[154] <= 32'b00101000000001101010110000100011;
ROM[155] <= 32'b00101000000001101010111000100011;
ROM[156] <= 32'b00101010000001101010000000100011;
ROM[157] <= 32'b00101010000001101010001000100011;
ROM[158] <= 32'b00101010000001101010010000100011;
ROM[159] <= 32'b00101010000001101010011000100011;
ROM[160] <= 32'b00101010000001101010100000100011;
ROM[161] <= 32'b00101010000001101010101000100011;
ROM[162] <= 32'b00101010000001101010110000100011;
ROM[163] <= 32'b00101010000001101010111000100011;
ROM[164] <= 32'b00101100000001101010000000100011;
ROM[165] <= 32'b00101100000001101010001000100011;
ROM[166] <= 32'b00101100000001101010010000100011;
ROM[167] <= 32'b00101100000001101010011000100011;
ROM[168] <= 32'b00101100000001101010100000100011;
ROM[169] <= 32'b00101100000001101010101000100011;
ROM[170] <= 32'b00101100000001101010110000100011;
ROM[171] <= 32'b00101100000001101010111000100011;
ROM[172] <= 32'b00101110000001101010000000100011;
ROM[173] <= 32'b00101110000001101010001000100011;
ROM[174] <= 32'b00101110000001101010010000100011;
ROM[175] <= 32'b00101110000001101010011000100011;
ROM[176] <= 32'b00101110000001101010100000100011;
ROM[177] <= 32'b00101110000001101010101000100011;
ROM[178] <= 32'b00101110000001101010110000100011;
ROM[179] <= 32'b00101110000001101010111000100011;
ROM[180] <= 32'b00110000000001101010000000100011;
ROM[181] <= 32'b00110000000001101010001000100011;
ROM[182] <= 32'b00110000000001101010010000100011;
ROM[183] <= 32'b00110000000001101010011000100011;
ROM[184] <= 32'b00110000000001101010100000100011;
ROM[185] <= 32'b00110000000001101010101000100011;
ROM[186] <= 32'b00110000000001101010110000100011;
ROM[187] <= 32'b00110000000001101010111000100011;
ROM[188] <= 32'b00110010000001101010000000100011;
ROM[189] <= 32'b00110010000001101010001000100011;
ROM[190] <= 32'b00110010000001101010010000100011;
ROM[191] <= 32'b00110010000001101010011000100011;
ROM[192] <= 32'b00110010000001101010100000100011;
ROM[193] <= 32'b00110010000001101010101000100011;
ROM[194] <= 32'b00110010000001101010110000100011;
ROM[195] <= 32'b00110010000001101010111000100011;
ROM[196] <= 32'b00110100000001101010000000100011;
ROM[197] <= 32'b00110100000001101010001000100011;
ROM[198] <= 32'b00110100000001101010010000100011;
ROM[199] <= 32'b00110100000001101010011000100011;
ROM[200] <= 32'b00110100000001101010100000100011;
ROM[201] <= 32'b00110100000001101010101000100011;
ROM[202] <= 32'b00110100000001101010110000100011;
ROM[203] <= 32'b00110100000001101010111000100011;
ROM[204] <= 32'b00110110000001101010000000100011;
ROM[205] <= 32'b00110110000001101010001000100011;
ROM[206] <= 32'b00110110000001101010010000100011;
ROM[207] <= 32'b00110110000001101010011000100011;
ROM[208] <= 32'b00110110000001101010100000100011;
ROM[209] <= 32'b00110110000001101010101000100011;
ROM[210] <= 32'b00110110000001101010110000100011;
ROM[211] <= 32'b00110110000001101010111000100011;
ROM[212] <= 32'b00111000000001101010000000100011;
ROM[213] <= 32'b00111000000001101010001000100011;
ROM[214] <= 32'b00111000000001101010010000100011;
ROM[215] <= 32'b00111000000001101010011000100011;
ROM[216] <= 32'b00111000000001101010100000100011;
ROM[217] <= 32'b00111000000001101010101000100011;
ROM[218] <= 32'b00111000000001101010110000100011;
ROM[219] <= 32'b00111000000001101010111000100011;
ROM[220] <= 32'b00111010000001101010000000100011;
ROM[221] <= 32'b00111010000001101010001000100011;
ROM[222] <= 32'b00111010000001101010010000100011;
ROM[223] <= 32'b00111010000001101010011000100011;
ROM[224] <= 32'b00111010000001101010100000100011;
ROM[225] <= 32'b00111010000001101010101000100011;
ROM[226] <= 32'b00111010000001101010110000100011;
ROM[227] <= 32'b00111010000001101010111000100011;
ROM[228] <= 32'b00111100000001101010000000100011;
ROM[229] <= 32'b00111100000001101010001000100011;
ROM[230] <= 32'b00111100000001101010010000100011;
ROM[231] <= 32'b00111100000001101010011000100011;
ROM[232] <= 32'b00111100000001101010100000100011;
ROM[233] <= 32'b00111100000001101010101000100011;
ROM[234] <= 32'b00111100000001101010110000100011;
ROM[235] <= 32'b00111100000001101010111000100011;
ROM[236] <= 32'b00111110000001101010000000100011;
ROM[237] <= 32'b00111110000001101010001000100011;
ROM[238] <= 32'b00111110000001101010010000100011;
ROM[239] <= 32'b00111110000001101010011000100011;
ROM[240] <= 32'b00111110000001101010100000100011;
ROM[241] <= 32'b00111110000001101010101000100011;
ROM[242] <= 32'b00111110000001101010110000100011;
ROM[243] <= 32'b00111110000001101010111000100011;
ROM[244] <= 32'b00000000000001101000011000010011;
ROM[245] <= 32'b01000000000001101000000100010011;
ROM[246] <= 32'b00000000000000010000000110010011;
ROM[247] <= 32'b00000000000000010000001000010011;
ROM[248] <= 32'b00000000000000010000001010010011;
ROM[249] <= 32'b00000000000000010000001100010011;
ROM[250] <= 32'b00000000000000000000001110110111;
ROM[251] <= 32'b01000011010000111000001110010011;
ROM[252] <= 32'b00000000111000111000001110110011;
ROM[253] <= 32'b00000000011100010010000000100011;
ROM[254] <= 32'b00000000010000010000000100010011;
ROM[255] <= 32'b00000000001100010010000000100011;
ROM[256] <= 32'b00000000010000010000000100010011;
ROM[257] <= 32'b00000000010000010010000000100011;
ROM[258] <= 32'b00000000010000010000000100010011;
ROM[259] <= 32'b00000000010100010010000000100011;
ROM[260] <= 32'b00000000010000010000000100010011;
ROM[261] <= 32'b00000000011000010010000000100011;
ROM[262] <= 32'b00000000010000010000000100010011;
ROM[263] <= 32'b00000001010000000000001110010011;
ROM[264] <= 32'b00000000000000111000001110010011;
ROM[265] <= 32'b01000000011100010000001110110011;
ROM[266] <= 32'b00000000011100000000001000110011;
ROM[267] <= 32'b00000000001000000000000110110011;
ROM[268] <= 32'b01110010010000000111000011101111;
ROM[269] <= 32'b11111111110000010000000100010011;
ROM[270] <= 32'b00000000000000010010001110000011;
ROM[271] <= 32'b00101100100100000111000011101111;
ROM[272] <= 32'b00000000000000100010001110000011;
ROM[273] <= 32'b00000000011100010010000000100011;
ROM[274] <= 32'b00000000010000010000000100010011;
ROM[275] <= 32'b00000000000000000000001110110111;
ROM[276] <= 32'b01001001100000111000001110010011;
ROM[277] <= 32'b00000000111000111000001110110011;
ROM[278] <= 32'b00000000011100010010000000100011;
ROM[279] <= 32'b00000000010000010000000100010011;
ROM[280] <= 32'b00000000001100010010000000100011;
ROM[281] <= 32'b00000000010000010000000100010011;
ROM[282] <= 32'b00000000010000010010000000100011;
ROM[283] <= 32'b00000000010000010000000100010011;
ROM[284] <= 32'b00000000010100010010000000100011;
ROM[285] <= 32'b00000000010000010000000100010011;
ROM[286] <= 32'b00000000011000010010000000100011;
ROM[287] <= 32'b00000000010000010000000100010011;
ROM[288] <= 32'b00000001010000000000001110010011;
ROM[289] <= 32'b00000000010000111000001110010011;
ROM[290] <= 32'b01000000011100010000001110110011;
ROM[291] <= 32'b00000000011100000000001000110011;
ROM[292] <= 32'b00000000001000000000000110110011;
ROM[293] <= 32'b01110100100100000010000011101111;
ROM[294] <= 32'b00000001010000000000001110010011;
ROM[295] <= 32'b01000000011100011000001110110011;
ROM[296] <= 32'b00000000000000111010000010000011;
ROM[297] <= 32'b11111111110000010000000100010011;
ROM[298] <= 32'b00000000000000010010001110000011;
ROM[299] <= 32'b00000000011100100010000000100011;
ROM[300] <= 32'b00000000010000100000000100010011;
ROM[301] <= 32'b00000001010000000000001110010011;
ROM[302] <= 32'b01000000011100011000001110110011;
ROM[303] <= 32'b00000000010000111010000110000011;
ROM[304] <= 32'b00000000100000111010001000000011;
ROM[305] <= 32'b00000000110000111010001010000011;
ROM[306] <= 32'b00000001000000111010001100000011;
ROM[307] <= 32'b00000000000000001000000011100111;
ROM[308] <= 32'b00000000000000010010000000100011;
ROM[309] <= 32'b00000000010000010000000100010011;
ROM[310] <= 32'b00000000000000010010000000100011;
ROM[311] <= 32'b00000000010000010000000100010011;
ROM[312] <= 32'b00000000011000000000001110010011;
ROM[313] <= 32'b00000000011100010010000000100011;
ROM[314] <= 32'b00000000010000010000000100010011;
ROM[315] <= 32'b00000000000000000000001110110111;
ROM[316] <= 32'b01010011100000111000001110010011;
ROM[317] <= 32'b00000000111000111000001110110011;
ROM[318] <= 32'b00000000011100010010000000100011;
ROM[319] <= 32'b00000000010000010000000100010011;
ROM[320] <= 32'b00000000001100010010000000100011;
ROM[321] <= 32'b00000000010000010000000100010011;
ROM[322] <= 32'b00000000010000010010000000100011;
ROM[323] <= 32'b00000000010000010000000100010011;
ROM[324] <= 32'b00000000010100010010000000100011;
ROM[325] <= 32'b00000000010000010000000100010011;
ROM[326] <= 32'b00000000011000010010000000100011;
ROM[327] <= 32'b00000000010000010000000100010011;
ROM[328] <= 32'b00000001010000000000001110010011;
ROM[329] <= 32'b00000000010000111000001110010011;
ROM[330] <= 32'b01000000011100010000001110110011;
ROM[331] <= 32'b00000000011100000000001000110011;
ROM[332] <= 32'b00000000001000000000000110110011;
ROM[333] <= 32'b00101110110000000110000011101111;
ROM[334] <= 32'b11111111110000010000000100010011;
ROM[335] <= 32'b00000000000000010010001110000011;
ROM[336] <= 32'b00000000011100011010000000100011;
ROM[337] <= 32'b00000000000000011010001110000011;
ROM[338] <= 32'b00000000011100010010000000100011;
ROM[339] <= 32'b00000000010000010000000100010011;
ROM[340] <= 32'b00000110000100000000001110010011;
ROM[341] <= 32'b00000000011100010010000000100011;
ROM[342] <= 32'b00000000010000010000000100010011;
ROM[343] <= 32'b00000000000000000000001110110111;
ROM[344] <= 32'b01011010100000111000001110010011;
ROM[345] <= 32'b00000000111000111000001110110011;
ROM[346] <= 32'b00000000011100010010000000100011;
ROM[347] <= 32'b00000000010000010000000100010011;
ROM[348] <= 32'b00000000001100010010000000100011;
ROM[349] <= 32'b00000000010000010000000100010011;
ROM[350] <= 32'b00000000010000010010000000100011;
ROM[351] <= 32'b00000000010000010000000100010011;
ROM[352] <= 32'b00000000010100010010000000100011;
ROM[353] <= 32'b00000000010000010000000100010011;
ROM[354] <= 32'b00000000011000010010000000100011;
ROM[355] <= 32'b00000000010000010000000100010011;
ROM[356] <= 32'b00000001010000000000001110010011;
ROM[357] <= 32'b00000000100000111000001110010011;
ROM[358] <= 32'b01000000011100010000001110110011;
ROM[359] <= 32'b00000000011100000000001000110011;
ROM[360] <= 32'b00000000001000000000000110110011;
ROM[361] <= 32'b01100001100000000110000011101111;
ROM[362] <= 32'b11111111110000010000000100010011;
ROM[363] <= 32'b00000000000000010010001110000011;
ROM[364] <= 32'b00000000011100011010001000100011;
ROM[365] <= 32'b00000000010000011010001110000011;
ROM[366] <= 32'b00000000011100010010000000100011;
ROM[367] <= 32'b00000000010000010000000100010011;
ROM[368] <= 32'b00000110111100000000001110010011;
ROM[369] <= 32'b00000000011100010010000000100011;
ROM[370] <= 32'b00000000010000010000000100010011;
ROM[371] <= 32'b00000001010000000000001110010011;
ROM[372] <= 32'b01000000011100011000001110110011;
ROM[373] <= 32'b00000000000000111010000010000011;
ROM[374] <= 32'b11111111110000010000000100010011;
ROM[375] <= 32'b00000000000000010010001110000011;
ROM[376] <= 32'b00000000011100100010000000100011;
ROM[377] <= 32'b00000000010000100000000100010011;
ROM[378] <= 32'b00000001010000000000001110010011;
ROM[379] <= 32'b01000000011100011000001110110011;
ROM[380] <= 32'b00000000010000111010000110000011;
ROM[381] <= 32'b00000000100000111010001000000011;
ROM[382] <= 32'b00000000110000111010001010000011;
ROM[383] <= 32'b00000001000000111010001100000011;
ROM[384] <= 32'b00000000000000001000000011100111;
ROM[385] <= 32'b00000001111100000000001110010011;
ROM[386] <= 32'b00000000011100010010000000100011;
ROM[387] <= 32'b00000000010000010000000100010011;
ROM[388] <= 32'b00000000000000000000001110110111;
ROM[389] <= 32'b01100101110000111000001110010011;
ROM[390] <= 32'b00000000111000111000001110110011;
ROM[391] <= 32'b00000000011100010010000000100011;
ROM[392] <= 32'b00000000010000010000000100010011;
ROM[393] <= 32'b00000000001100010010000000100011;
ROM[394] <= 32'b00000000010000010000000100010011;
ROM[395] <= 32'b00000000010000010010000000100011;
ROM[396] <= 32'b00000000010000010000000100010011;
ROM[397] <= 32'b00000000010100010010000000100011;
ROM[398] <= 32'b00000000010000010000000100010011;
ROM[399] <= 32'b00000000011000010010000000100011;
ROM[400] <= 32'b00000000010000010000000100010011;
ROM[401] <= 32'b00000001010000000000001110010011;
ROM[402] <= 32'b00000000010000111000001110010011;
ROM[403] <= 32'b01000000011100010000001110110011;
ROM[404] <= 32'b00000000011100000000001000110011;
ROM[405] <= 32'b00000000001000000000000110110011;
ROM[406] <= 32'b11011110100111111111000011101111;
ROM[407] <= 32'b11111111110000010000000100010011;
ROM[408] <= 32'b00000000000000010010001110000011;
ROM[409] <= 32'b00000100011101101010000000100011;
ROM[410] <= 32'b00000000000000000000001110010011;
ROM[411] <= 32'b00000000011100010010000000100011;
ROM[412] <= 32'b00000000010000010000000100010011;
ROM[413] <= 32'b00000100000001101010001110000011;
ROM[414] <= 32'b00000000011100010010000000100011;
ROM[415] <= 32'b00000000010000010000000100010011;
ROM[416] <= 32'b11111111110000010000000100010011;
ROM[417] <= 32'b00000000000000010010001110000011;
ROM[418] <= 32'b11111111110000010000000100010011;
ROM[419] <= 32'b00000000000000010010010000000011;
ROM[420] <= 32'b00000000011101000000001110110011;
ROM[421] <= 32'b00000000011100010010000000100011;
ROM[422] <= 32'b00000000010000010000000100010011;
ROM[423] <= 32'b00000000000100000000001110010011;
ROM[424] <= 32'b00000000011100010010000000100011;
ROM[425] <= 32'b00000000010000010000000100010011;
ROM[426] <= 32'b11111111110000010000000100010011;
ROM[427] <= 32'b00000000000000010010001110000011;
ROM[428] <= 32'b00000000011101100010000000100011;
ROM[429] <= 32'b11111111110000010000000100010011;
ROM[430] <= 32'b00000000000000010010001110000011;
ROM[431] <= 32'b00000000000000111000001100010011;
ROM[432] <= 32'b00000000000001100010001110000011;
ROM[433] <= 32'b00000000011100010010000000100011;
ROM[434] <= 32'b00000000010000010000000100010011;
ROM[435] <= 32'b11111111110000010000000100010011;
ROM[436] <= 32'b00000000000000010010001110000011;
ROM[437] <= 32'b00000000110100110000010000110011;
ROM[438] <= 32'b00000000011101000010000000100011;
ROM[439] <= 32'b00000000010000000000001110010011;
ROM[440] <= 32'b00000000011100010010000000100011;
ROM[441] <= 32'b00000000010000010000000100010011;
ROM[442] <= 32'b00000100000001101010001110000011;
ROM[443] <= 32'b00000000011100010010000000100011;
ROM[444] <= 32'b00000000010000010000000100010011;
ROM[445] <= 32'b11111111110000010000000100010011;
ROM[446] <= 32'b00000000000000010010001110000011;
ROM[447] <= 32'b11111111110000010000000100010011;
ROM[448] <= 32'b00000000000000010010010000000011;
ROM[449] <= 32'b00000000011101000000001110110011;
ROM[450] <= 32'b00000000011100010010000000100011;
ROM[451] <= 32'b00000000010000010000000100010011;
ROM[452] <= 32'b00000000001000000000001110010011;
ROM[453] <= 32'b00000000011100010010000000100011;
ROM[454] <= 32'b00000000010000010000000100010011;
ROM[455] <= 32'b11111111110000010000000100010011;
ROM[456] <= 32'b00000000000000010010001110000011;
ROM[457] <= 32'b00000000011101100010000000100011;
ROM[458] <= 32'b11111111110000010000000100010011;
ROM[459] <= 32'b00000000000000010010001110000011;
ROM[460] <= 32'b00000000000000111000001100010011;
ROM[461] <= 32'b00000000000001100010001110000011;
ROM[462] <= 32'b00000000011100010010000000100011;
ROM[463] <= 32'b00000000010000010000000100010011;
ROM[464] <= 32'b11111111110000010000000100010011;
ROM[465] <= 32'b00000000000000010010001110000011;
ROM[466] <= 32'b00000000110100110000010000110011;
ROM[467] <= 32'b00000000011101000010000000100011;
ROM[468] <= 32'b00000000100000000000001110010011;
ROM[469] <= 32'b00000000011100010010000000100011;
ROM[470] <= 32'b00000000010000010000000100010011;
ROM[471] <= 32'b00000100000001101010001110000011;
ROM[472] <= 32'b00000000011100010010000000100011;
ROM[473] <= 32'b00000000010000010000000100010011;
ROM[474] <= 32'b11111111110000010000000100010011;
ROM[475] <= 32'b00000000000000010010001110000011;
ROM[476] <= 32'b11111111110000010000000100010011;
ROM[477] <= 32'b00000000000000010010010000000011;
ROM[478] <= 32'b00000000011101000000001110110011;
ROM[479] <= 32'b00000000011100010010000000100011;
ROM[480] <= 32'b00000000010000010000000100010011;
ROM[481] <= 32'b00000000010000000000001110010011;
ROM[482] <= 32'b00000000011100010010000000100011;
ROM[483] <= 32'b00000000010000010000000100010011;
ROM[484] <= 32'b11111111110000010000000100010011;
ROM[485] <= 32'b00000000000000010010001110000011;
ROM[486] <= 32'b00000000011101100010000000100011;
ROM[487] <= 32'b11111111110000010000000100010011;
ROM[488] <= 32'b00000000000000010010001110000011;
ROM[489] <= 32'b00000000000000111000001100010011;
ROM[490] <= 32'b00000000000001100010001110000011;
ROM[491] <= 32'b00000000011100010010000000100011;
ROM[492] <= 32'b00000000010000010000000100010011;
ROM[493] <= 32'b11111111110000010000000100010011;
ROM[494] <= 32'b00000000000000010010001110000011;
ROM[495] <= 32'b00000000110100110000010000110011;
ROM[496] <= 32'b00000000011101000010000000100011;
ROM[497] <= 32'b00000000110000000000001110010011;
ROM[498] <= 32'b00000000011100010010000000100011;
ROM[499] <= 32'b00000000010000010000000100010011;
ROM[500] <= 32'b00000100000001101010001110000011;
ROM[501] <= 32'b00000000011100010010000000100011;
ROM[502] <= 32'b00000000010000010000000100010011;
ROM[503] <= 32'b11111111110000010000000100010011;
ROM[504] <= 32'b00000000000000010010001110000011;
ROM[505] <= 32'b11111111110000010000000100010011;
ROM[506] <= 32'b00000000000000010010010000000011;
ROM[507] <= 32'b00000000011101000000001110110011;
ROM[508] <= 32'b00000000011100010010000000100011;
ROM[509] <= 32'b00000000010000010000000100010011;
ROM[510] <= 32'b00000000100000000000001110010011;
ROM[511] <= 32'b00000000011100010010000000100011;
ROM[512] <= 32'b00000000010000010000000100010011;
ROM[513] <= 32'b11111111110000010000000100010011;
ROM[514] <= 32'b00000000000000010010001110000011;
ROM[515] <= 32'b00000000011101100010000000100011;
ROM[516] <= 32'b11111111110000010000000100010011;
ROM[517] <= 32'b00000000000000010010001110000011;
ROM[518] <= 32'b00000000000000111000001100010011;
ROM[519] <= 32'b00000000000001100010001110000011;
ROM[520] <= 32'b00000000011100010010000000100011;
ROM[521] <= 32'b00000000010000010000000100010011;
ROM[522] <= 32'b11111111110000010000000100010011;
ROM[523] <= 32'b00000000000000010010001110000011;
ROM[524] <= 32'b00000000110100110000010000110011;
ROM[525] <= 32'b00000000011101000010000000100011;
ROM[526] <= 32'b00000001000000000000001110010011;
ROM[527] <= 32'b00000000011100010010000000100011;
ROM[528] <= 32'b00000000010000010000000100010011;
ROM[529] <= 32'b00000100000001101010001110000011;
ROM[530] <= 32'b00000000011100010010000000100011;
ROM[531] <= 32'b00000000010000010000000100010011;
ROM[532] <= 32'b11111111110000010000000100010011;
ROM[533] <= 32'b00000000000000010010001110000011;
ROM[534] <= 32'b11111111110000010000000100010011;
ROM[535] <= 32'b00000000000000010010010000000011;
ROM[536] <= 32'b00000000011101000000001110110011;
ROM[537] <= 32'b00000000011100010010000000100011;
ROM[538] <= 32'b00000000010000010000000100010011;
ROM[539] <= 32'b00000001000000000000001110010011;
ROM[540] <= 32'b00000000011100010010000000100011;
ROM[541] <= 32'b00000000010000010000000100010011;
ROM[542] <= 32'b11111111110000010000000100010011;
ROM[543] <= 32'b00000000000000010010001110000011;
ROM[544] <= 32'b00000000011101100010000000100011;
ROM[545] <= 32'b11111111110000010000000100010011;
ROM[546] <= 32'b00000000000000010010001110000011;
ROM[547] <= 32'b00000000000000111000001100010011;
ROM[548] <= 32'b00000000000001100010001110000011;
ROM[549] <= 32'b00000000011100010010000000100011;
ROM[550] <= 32'b00000000010000010000000100010011;
ROM[551] <= 32'b11111111110000010000000100010011;
ROM[552] <= 32'b00000000000000010010001110000011;
ROM[553] <= 32'b00000000110100110000010000110011;
ROM[554] <= 32'b00000000011101000010000000100011;
ROM[555] <= 32'b00000001010000000000001110010011;
ROM[556] <= 32'b00000000011100010010000000100011;
ROM[557] <= 32'b00000000010000010000000100010011;
ROM[558] <= 32'b00000100000001101010001110000011;
ROM[559] <= 32'b00000000011100010010000000100011;
ROM[560] <= 32'b00000000010000010000000100010011;
ROM[561] <= 32'b11111111110000010000000100010011;
ROM[562] <= 32'b00000000000000010010001110000011;
ROM[563] <= 32'b11111111110000010000000100010011;
ROM[564] <= 32'b00000000000000010010010000000011;
ROM[565] <= 32'b00000000011101000000001110110011;
ROM[566] <= 32'b00000000011100010010000000100011;
ROM[567] <= 32'b00000000010000010000000100010011;
ROM[568] <= 32'b00000010000000000000001110010011;
ROM[569] <= 32'b00000000011100010010000000100011;
ROM[570] <= 32'b00000000010000010000000100010011;
ROM[571] <= 32'b11111111110000010000000100010011;
ROM[572] <= 32'b00000000000000010010001110000011;
ROM[573] <= 32'b00000000011101100010000000100011;
ROM[574] <= 32'b11111111110000010000000100010011;
ROM[575] <= 32'b00000000000000010010001110000011;
ROM[576] <= 32'b00000000000000111000001100010011;
ROM[577] <= 32'b00000000000001100010001110000011;
ROM[578] <= 32'b00000000011100010010000000100011;
ROM[579] <= 32'b00000000010000010000000100010011;
ROM[580] <= 32'b11111111110000010000000100010011;
ROM[581] <= 32'b00000000000000010010001110000011;
ROM[582] <= 32'b00000000110100110000010000110011;
ROM[583] <= 32'b00000000011101000010000000100011;
ROM[584] <= 32'b00000001100000000000001110010011;
ROM[585] <= 32'b00000000011100010010000000100011;
ROM[586] <= 32'b00000000010000010000000100010011;
ROM[587] <= 32'b00000100000001101010001110000011;
ROM[588] <= 32'b00000000011100010010000000100011;
ROM[589] <= 32'b00000000010000010000000100010011;
ROM[590] <= 32'b11111111110000010000000100010011;
ROM[591] <= 32'b00000000000000010010001110000011;
ROM[592] <= 32'b11111111110000010000000100010011;
ROM[593] <= 32'b00000000000000010010010000000011;
ROM[594] <= 32'b00000000011101000000001110110011;
ROM[595] <= 32'b00000000011100010010000000100011;
ROM[596] <= 32'b00000000010000010000000100010011;
ROM[597] <= 32'b00000100000000000000001110010011;
ROM[598] <= 32'b00000000011100010010000000100011;
ROM[599] <= 32'b00000000010000010000000100010011;
ROM[600] <= 32'b11111111110000010000000100010011;
ROM[601] <= 32'b00000000000000010010001110000011;
ROM[602] <= 32'b00000000011101100010000000100011;
ROM[603] <= 32'b11111111110000010000000100010011;
ROM[604] <= 32'b00000000000000010010001110000011;
ROM[605] <= 32'b00000000000000111000001100010011;
ROM[606] <= 32'b00000000000001100010001110000011;
ROM[607] <= 32'b00000000011100010010000000100011;
ROM[608] <= 32'b00000000010000010000000100010011;
ROM[609] <= 32'b11111111110000010000000100010011;
ROM[610] <= 32'b00000000000000010010001110000011;
ROM[611] <= 32'b00000000110100110000010000110011;
ROM[612] <= 32'b00000000011101000010000000100011;
ROM[613] <= 32'b00000001110000000000001110010011;
ROM[614] <= 32'b00000000011100010010000000100011;
ROM[615] <= 32'b00000000010000010000000100010011;
ROM[616] <= 32'b00000100000001101010001110000011;
ROM[617] <= 32'b00000000011100010010000000100011;
ROM[618] <= 32'b00000000010000010000000100010011;
ROM[619] <= 32'b11111111110000010000000100010011;
ROM[620] <= 32'b00000000000000010010001110000011;
ROM[621] <= 32'b11111111110000010000000100010011;
ROM[622] <= 32'b00000000000000010010010000000011;
ROM[623] <= 32'b00000000011101000000001110110011;
ROM[624] <= 32'b00000000011100010010000000100011;
ROM[625] <= 32'b00000000010000010000000100010011;
ROM[626] <= 32'b00001000000000000000001110010011;
ROM[627] <= 32'b00000000011100010010000000100011;
ROM[628] <= 32'b00000000010000010000000100010011;
ROM[629] <= 32'b11111111110000010000000100010011;
ROM[630] <= 32'b00000000000000010010001110000011;
ROM[631] <= 32'b00000000011101100010000000100011;
ROM[632] <= 32'b11111111110000010000000100010011;
ROM[633] <= 32'b00000000000000010010001110000011;
ROM[634] <= 32'b00000000000000111000001100010011;
ROM[635] <= 32'b00000000000001100010001110000011;
ROM[636] <= 32'b00000000011100010010000000100011;
ROM[637] <= 32'b00000000010000010000000100010011;
ROM[638] <= 32'b11111111110000010000000100010011;
ROM[639] <= 32'b00000000000000010010001110000011;
ROM[640] <= 32'b00000000110100110000010000110011;
ROM[641] <= 32'b00000000011101000010000000100011;
ROM[642] <= 32'b00000010000000000000001110010011;
ROM[643] <= 32'b00000000011100010010000000100011;
ROM[644] <= 32'b00000000010000010000000100010011;
ROM[645] <= 32'b00000100000001101010001110000011;
ROM[646] <= 32'b00000000011100010010000000100011;
ROM[647] <= 32'b00000000010000010000000100010011;
ROM[648] <= 32'b11111111110000010000000100010011;
ROM[649] <= 32'b00000000000000010010001110000011;
ROM[650] <= 32'b11111111110000010000000100010011;
ROM[651] <= 32'b00000000000000010010010000000011;
ROM[652] <= 32'b00000000011101000000001110110011;
ROM[653] <= 32'b00000000011100010010000000100011;
ROM[654] <= 32'b00000000010000010000000100010011;
ROM[655] <= 32'b00010000000000000000001110010011;
ROM[656] <= 32'b00000000011100010010000000100011;
ROM[657] <= 32'b00000000010000010000000100010011;
ROM[658] <= 32'b11111111110000010000000100010011;
ROM[659] <= 32'b00000000000000010010001110000011;
ROM[660] <= 32'b00000000011101100010000000100011;
ROM[661] <= 32'b11111111110000010000000100010011;
ROM[662] <= 32'b00000000000000010010001110000011;
ROM[663] <= 32'b00000000000000111000001100010011;
ROM[664] <= 32'b00000000000001100010001110000011;
ROM[665] <= 32'b00000000011100010010000000100011;
ROM[666] <= 32'b00000000010000010000000100010011;
ROM[667] <= 32'b11111111110000010000000100010011;
ROM[668] <= 32'b00000000000000010010001110000011;
ROM[669] <= 32'b00000000110100110000010000110011;
ROM[670] <= 32'b00000000011101000010000000100011;
ROM[671] <= 32'b00000010010000000000001110010011;
ROM[672] <= 32'b00000000011100010010000000100011;
ROM[673] <= 32'b00000000010000010000000100010011;
ROM[674] <= 32'b00000100000001101010001110000011;
ROM[675] <= 32'b00000000011100010010000000100011;
ROM[676] <= 32'b00000000010000010000000100010011;
ROM[677] <= 32'b11111111110000010000000100010011;
ROM[678] <= 32'b00000000000000010010001110000011;
ROM[679] <= 32'b11111111110000010000000100010011;
ROM[680] <= 32'b00000000000000010010010000000011;
ROM[681] <= 32'b00000000011101000000001110110011;
ROM[682] <= 32'b00000000011100010010000000100011;
ROM[683] <= 32'b00000000010000010000000100010011;
ROM[684] <= 32'b00100000000000000000001110010011;
ROM[685] <= 32'b00000000011100010010000000100011;
ROM[686] <= 32'b00000000010000010000000100010011;
ROM[687] <= 32'b11111111110000010000000100010011;
ROM[688] <= 32'b00000000000000010010001110000011;
ROM[689] <= 32'b00000000011101100010000000100011;
ROM[690] <= 32'b11111111110000010000000100010011;
ROM[691] <= 32'b00000000000000010010001110000011;
ROM[692] <= 32'b00000000000000111000001100010011;
ROM[693] <= 32'b00000000000001100010001110000011;
ROM[694] <= 32'b00000000011100010010000000100011;
ROM[695] <= 32'b00000000010000010000000100010011;
ROM[696] <= 32'b11111111110000010000000100010011;
ROM[697] <= 32'b00000000000000010010001110000011;
ROM[698] <= 32'b00000000110100110000010000110011;
ROM[699] <= 32'b00000000011101000010000000100011;
ROM[700] <= 32'b00000010100000000000001110010011;
ROM[701] <= 32'b00000000011100010010000000100011;
ROM[702] <= 32'b00000000010000010000000100010011;
ROM[703] <= 32'b00000100000001101010001110000011;
ROM[704] <= 32'b00000000011100010010000000100011;
ROM[705] <= 32'b00000000010000010000000100010011;
ROM[706] <= 32'b11111111110000010000000100010011;
ROM[707] <= 32'b00000000000000010010001110000011;
ROM[708] <= 32'b11111111110000010000000100010011;
ROM[709] <= 32'b00000000000000010010010000000011;
ROM[710] <= 32'b00000000011101000000001110110011;
ROM[711] <= 32'b00000000011100010010000000100011;
ROM[712] <= 32'b00000000010000010000000100010011;
ROM[713] <= 32'b01000000000000000000001110010011;
ROM[714] <= 32'b00000000011100010010000000100011;
ROM[715] <= 32'b00000000010000010000000100010011;
ROM[716] <= 32'b11111111110000010000000100010011;
ROM[717] <= 32'b00000000000000010010001110000011;
ROM[718] <= 32'b00000000011101100010000000100011;
ROM[719] <= 32'b11111111110000010000000100010011;
ROM[720] <= 32'b00000000000000010010001110000011;
ROM[721] <= 32'b00000000000000111000001100010011;
ROM[722] <= 32'b00000000000001100010001110000011;
ROM[723] <= 32'b00000000011100010010000000100011;
ROM[724] <= 32'b00000000010000010000000100010011;
ROM[725] <= 32'b11111111110000010000000100010011;
ROM[726] <= 32'b00000000000000010010001110000011;
ROM[727] <= 32'b00000000110100110000010000110011;
ROM[728] <= 32'b00000000011101000010000000100011;
ROM[729] <= 32'b00000010110000000000001110010011;
ROM[730] <= 32'b00000000011100010010000000100011;
ROM[731] <= 32'b00000000010000010000000100010011;
ROM[732] <= 32'b00000100000001101010001110000011;
ROM[733] <= 32'b00000000011100010010000000100011;
ROM[734] <= 32'b00000000010000010000000100010011;
ROM[735] <= 32'b11111111110000010000000100010011;
ROM[736] <= 32'b00000000000000010010001110000011;
ROM[737] <= 32'b11111111110000010000000100010011;
ROM[738] <= 32'b00000000000000010010010000000011;
ROM[739] <= 32'b00000000011101000000001110110011;
ROM[740] <= 32'b00000000011100010010000000100011;
ROM[741] <= 32'b00000000010000010000000100010011;
ROM[742] <= 32'b00000000000000000001001110110111;
ROM[743] <= 32'b10000000000000111000001110010011;
ROM[744] <= 32'b00000000011100010010000000100011;
ROM[745] <= 32'b00000000010000010000000100010011;
ROM[746] <= 32'b11111111110000010000000100010011;
ROM[747] <= 32'b00000000000000010010001110000011;
ROM[748] <= 32'b00000000011101100010000000100011;
ROM[749] <= 32'b11111111110000010000000100010011;
ROM[750] <= 32'b00000000000000010010001110000011;
ROM[751] <= 32'b00000000000000111000001100010011;
ROM[752] <= 32'b00000000000001100010001110000011;
ROM[753] <= 32'b00000000011100010010000000100011;
ROM[754] <= 32'b00000000010000010000000100010011;
ROM[755] <= 32'b11111111110000010000000100010011;
ROM[756] <= 32'b00000000000000010010001110000011;
ROM[757] <= 32'b00000000110100110000010000110011;
ROM[758] <= 32'b00000000011101000010000000100011;
ROM[759] <= 32'b00000011000000000000001110010011;
ROM[760] <= 32'b00000000011100010010000000100011;
ROM[761] <= 32'b00000000010000010000000100010011;
ROM[762] <= 32'b00000100000001101010001110000011;
ROM[763] <= 32'b00000000011100010010000000100011;
ROM[764] <= 32'b00000000010000010000000100010011;
ROM[765] <= 32'b11111111110000010000000100010011;
ROM[766] <= 32'b00000000000000010010001110000011;
ROM[767] <= 32'b11111111110000010000000100010011;
ROM[768] <= 32'b00000000000000010010010000000011;
ROM[769] <= 32'b00000000011101000000001110110011;
ROM[770] <= 32'b00000000011100010010000000100011;
ROM[771] <= 32'b00000000010000010000000100010011;
ROM[772] <= 32'b00000000000000000001001110110111;
ROM[773] <= 32'b00000000000000111000001110010011;
ROM[774] <= 32'b00000000011100010010000000100011;
ROM[775] <= 32'b00000000010000010000000100010011;
ROM[776] <= 32'b11111111110000010000000100010011;
ROM[777] <= 32'b00000000000000010010001110000011;
ROM[778] <= 32'b00000000011101100010000000100011;
ROM[779] <= 32'b11111111110000010000000100010011;
ROM[780] <= 32'b00000000000000010010001110000011;
ROM[781] <= 32'b00000000000000111000001100010011;
ROM[782] <= 32'b00000000000001100010001110000011;
ROM[783] <= 32'b00000000011100010010000000100011;
ROM[784] <= 32'b00000000010000010000000100010011;
ROM[785] <= 32'b11111111110000010000000100010011;
ROM[786] <= 32'b00000000000000010010001110000011;
ROM[787] <= 32'b00000000110100110000010000110011;
ROM[788] <= 32'b00000000011101000010000000100011;
ROM[789] <= 32'b00000011010000000000001110010011;
ROM[790] <= 32'b00000000011100010010000000100011;
ROM[791] <= 32'b00000000010000010000000100010011;
ROM[792] <= 32'b00000100000001101010001110000011;
ROM[793] <= 32'b00000000011100010010000000100011;
ROM[794] <= 32'b00000000010000010000000100010011;
ROM[795] <= 32'b11111111110000010000000100010011;
ROM[796] <= 32'b00000000000000010010001110000011;
ROM[797] <= 32'b11111111110000010000000100010011;
ROM[798] <= 32'b00000000000000010010010000000011;
ROM[799] <= 32'b00000000011101000000001110110011;
ROM[800] <= 32'b00000000011100010010000000100011;
ROM[801] <= 32'b00000000010000010000000100010011;
ROM[802] <= 32'b00000000000000000010001110110111;
ROM[803] <= 32'b00000000000000111000001110010011;
ROM[804] <= 32'b00000000011100010010000000100011;
ROM[805] <= 32'b00000000010000010000000100010011;
ROM[806] <= 32'b11111111110000010000000100010011;
ROM[807] <= 32'b00000000000000010010001110000011;
ROM[808] <= 32'b00000000011101100010000000100011;
ROM[809] <= 32'b11111111110000010000000100010011;
ROM[810] <= 32'b00000000000000010010001110000011;
ROM[811] <= 32'b00000000000000111000001100010011;
ROM[812] <= 32'b00000000000001100010001110000011;
ROM[813] <= 32'b00000000011100010010000000100011;
ROM[814] <= 32'b00000000010000010000000100010011;
ROM[815] <= 32'b11111111110000010000000100010011;
ROM[816] <= 32'b00000000000000010010001110000011;
ROM[817] <= 32'b00000000110100110000010000110011;
ROM[818] <= 32'b00000000011101000010000000100011;
ROM[819] <= 32'b00000011100000000000001110010011;
ROM[820] <= 32'b00000000011100010010000000100011;
ROM[821] <= 32'b00000000010000010000000100010011;
ROM[822] <= 32'b00000100000001101010001110000011;
ROM[823] <= 32'b00000000011100010010000000100011;
ROM[824] <= 32'b00000000010000010000000100010011;
ROM[825] <= 32'b11111111110000010000000100010011;
ROM[826] <= 32'b00000000000000010010001110000011;
ROM[827] <= 32'b11111111110000010000000100010011;
ROM[828] <= 32'b00000000000000010010010000000011;
ROM[829] <= 32'b00000000011101000000001110110011;
ROM[830] <= 32'b00000000011100010010000000100011;
ROM[831] <= 32'b00000000010000010000000100010011;
ROM[832] <= 32'b00000000000000000100001110110111;
ROM[833] <= 32'b00000000000000111000001110010011;
ROM[834] <= 32'b00000000011100010010000000100011;
ROM[835] <= 32'b00000000010000010000000100010011;
ROM[836] <= 32'b11111111110000010000000100010011;
ROM[837] <= 32'b00000000000000010010001110000011;
ROM[838] <= 32'b00000000011101100010000000100011;
ROM[839] <= 32'b11111111110000010000000100010011;
ROM[840] <= 32'b00000000000000010010001110000011;
ROM[841] <= 32'b00000000000000111000001100010011;
ROM[842] <= 32'b00000000000001100010001110000011;
ROM[843] <= 32'b00000000011100010010000000100011;
ROM[844] <= 32'b00000000010000010000000100010011;
ROM[845] <= 32'b11111111110000010000000100010011;
ROM[846] <= 32'b00000000000000010010001110000011;
ROM[847] <= 32'b00000000110100110000010000110011;
ROM[848] <= 32'b00000000011101000010000000100011;
ROM[849] <= 32'b00000011110000000000001110010011;
ROM[850] <= 32'b00000000011100010010000000100011;
ROM[851] <= 32'b00000000010000010000000100010011;
ROM[852] <= 32'b00000100000001101010001110000011;
ROM[853] <= 32'b00000000011100010010000000100011;
ROM[854] <= 32'b00000000010000010000000100010011;
ROM[855] <= 32'b11111111110000010000000100010011;
ROM[856] <= 32'b00000000000000010010001110000011;
ROM[857] <= 32'b11111111110000010000000100010011;
ROM[858] <= 32'b00000000000000010010010000000011;
ROM[859] <= 32'b00000000011101000000001110110011;
ROM[860] <= 32'b00000000011100010010000000100011;
ROM[861] <= 32'b00000000010000010000000100010011;
ROM[862] <= 32'b00000000000000000100001110110111;
ROM[863] <= 32'b00000000000000111000001110010011;
ROM[864] <= 32'b00000000011100010010000000100011;
ROM[865] <= 32'b00000000010000010000000100010011;
ROM[866] <= 32'b00000000000000000100001110110111;
ROM[867] <= 32'b00000000000000111000001110010011;
ROM[868] <= 32'b00000000011100010010000000100011;
ROM[869] <= 32'b00000000010000010000000100010011;
ROM[870] <= 32'b11111111110000010000000100010011;
ROM[871] <= 32'b00000000000000010010001110000011;
ROM[872] <= 32'b11111111110000010000000100010011;
ROM[873] <= 32'b00000000000000010010010000000011;
ROM[874] <= 32'b00000000011101000000001110110011;
ROM[875] <= 32'b00000000011100010010000000100011;
ROM[876] <= 32'b00000000010000010000000100010011;
ROM[877] <= 32'b11111111110000010000000100010011;
ROM[878] <= 32'b00000000000000010010001110000011;
ROM[879] <= 32'b00000000011101100010000000100011;
ROM[880] <= 32'b11111111110000010000000100010011;
ROM[881] <= 32'b00000000000000010010001110000011;
ROM[882] <= 32'b00000000000000111000001100010011;
ROM[883] <= 32'b00000000000001100010001110000011;
ROM[884] <= 32'b00000000011100010010000000100011;
ROM[885] <= 32'b00000000010000010000000100010011;
ROM[886] <= 32'b11111111110000010000000100010011;
ROM[887] <= 32'b00000000000000010010001110000011;
ROM[888] <= 32'b00000000110100110000010000110011;
ROM[889] <= 32'b00000000011101000010000000100011;
ROM[890] <= 32'b00000100000000000000001110010011;
ROM[891] <= 32'b00000000011100010010000000100011;
ROM[892] <= 32'b00000000010000010000000100010011;
ROM[893] <= 32'b00000100000001101010001110000011;
ROM[894] <= 32'b00000000011100010010000000100011;
ROM[895] <= 32'b00000000010000010000000100010011;
ROM[896] <= 32'b11111111110000010000000100010011;
ROM[897] <= 32'b00000000000000010010001110000011;
ROM[898] <= 32'b11111111110000010000000100010011;
ROM[899] <= 32'b00000000000000010010010000000011;
ROM[900] <= 32'b00000000011101000000001110110011;
ROM[901] <= 32'b00000000011100010010000000100011;
ROM[902] <= 32'b00000000010000010000000100010011;
ROM[903] <= 32'b00000011110000000000001110010011;
ROM[904] <= 32'b00000000011100010010000000100011;
ROM[905] <= 32'b00000000010000010000000100010011;
ROM[906] <= 32'b00000100000001101010001110000011;
ROM[907] <= 32'b00000000011100010010000000100011;
ROM[908] <= 32'b00000000010000010000000100010011;
ROM[909] <= 32'b11111111110000010000000100010011;
ROM[910] <= 32'b00000000000000010010001110000011;
ROM[911] <= 32'b11111111110000010000000100010011;
ROM[912] <= 32'b00000000000000010010010000000011;
ROM[913] <= 32'b00000000011101000000001110110011;
ROM[914] <= 32'b00000000011100010010000000100011;
ROM[915] <= 32'b00000000010000010000000100010011;
ROM[916] <= 32'b11111111110000010000000100010011;
ROM[917] <= 32'b00000000000000010010001110000011;
ROM[918] <= 32'b00000000000000111000001100010011;
ROM[919] <= 32'b00000000110100110000010000110011;
ROM[920] <= 32'b00000000000001000010001110000011;
ROM[921] <= 32'b00000000011100010010000000100011;
ROM[922] <= 32'b00000000010000010000000100010011;
ROM[923] <= 32'b00000011110000000000001110010011;
ROM[924] <= 32'b00000000011100010010000000100011;
ROM[925] <= 32'b00000000010000010000000100010011;
ROM[926] <= 32'b00000100000001101010001110000011;
ROM[927] <= 32'b00000000011100010010000000100011;
ROM[928] <= 32'b00000000010000010000000100010011;
ROM[929] <= 32'b11111111110000010000000100010011;
ROM[930] <= 32'b00000000000000010010001110000011;
ROM[931] <= 32'b11111111110000010000000100010011;
ROM[932] <= 32'b00000000000000010010010000000011;
ROM[933] <= 32'b00000000011101000000001110110011;
ROM[934] <= 32'b00000000011100010010000000100011;
ROM[935] <= 32'b00000000010000010000000100010011;
ROM[936] <= 32'b11111111110000010000000100010011;
ROM[937] <= 32'b00000000000000010010001110000011;
ROM[938] <= 32'b00000000000000111000001100010011;
ROM[939] <= 32'b00000000110100110000010000110011;
ROM[940] <= 32'b00000000000001000010001110000011;
ROM[941] <= 32'b00000000011100010010000000100011;
ROM[942] <= 32'b00000000010000010000000100010011;
ROM[943] <= 32'b11111111110000010000000100010011;
ROM[944] <= 32'b00000000000000010010001110000011;
ROM[945] <= 32'b11111111110000010000000100010011;
ROM[946] <= 32'b00000000000000010010010000000011;
ROM[947] <= 32'b00000000011101000000001110110011;
ROM[948] <= 32'b00000000011100010010000000100011;
ROM[949] <= 32'b00000000010000010000000100010011;
ROM[950] <= 32'b11111111110000010000000100010011;
ROM[951] <= 32'b00000000000000010010001110000011;
ROM[952] <= 32'b00000000011101100010000000100011;
ROM[953] <= 32'b11111111110000010000000100010011;
ROM[954] <= 32'b00000000000000010010001110000011;
ROM[955] <= 32'b00000000000000111000001100010011;
ROM[956] <= 32'b00000000000001100010001110000011;
ROM[957] <= 32'b00000000011100010010000000100011;
ROM[958] <= 32'b00000000010000010000000100010011;
ROM[959] <= 32'b11111111110000010000000100010011;
ROM[960] <= 32'b00000000000000010010001110000011;
ROM[961] <= 32'b00000000110100110000010000110011;
ROM[962] <= 32'b00000000011101000010000000100011;
ROM[963] <= 32'b00000100010000000000001110010011;
ROM[964] <= 32'b00000000011100010010000000100011;
ROM[965] <= 32'b00000000010000010000000100010011;
ROM[966] <= 32'b00000100000001101010001110000011;
ROM[967] <= 32'b00000000011100010010000000100011;
ROM[968] <= 32'b00000000010000010000000100010011;
ROM[969] <= 32'b11111111110000010000000100010011;
ROM[970] <= 32'b00000000000000010010001110000011;
ROM[971] <= 32'b11111111110000010000000100010011;
ROM[972] <= 32'b00000000000000010010010000000011;
ROM[973] <= 32'b00000000011101000000001110110011;
ROM[974] <= 32'b00000000011100010010000000100011;
ROM[975] <= 32'b00000000010000010000000100010011;
ROM[976] <= 32'b00000100000000000000001110010011;
ROM[977] <= 32'b00000000011100010010000000100011;
ROM[978] <= 32'b00000000010000010000000100010011;
ROM[979] <= 32'b00000100000001101010001110000011;
ROM[980] <= 32'b00000000011100010010000000100011;
ROM[981] <= 32'b00000000010000010000000100010011;
ROM[982] <= 32'b11111111110000010000000100010011;
ROM[983] <= 32'b00000000000000010010001110000011;
ROM[984] <= 32'b11111111110000010000000100010011;
ROM[985] <= 32'b00000000000000010010010000000011;
ROM[986] <= 32'b00000000011101000000001110110011;
ROM[987] <= 32'b00000000011100010010000000100011;
ROM[988] <= 32'b00000000010000010000000100010011;
ROM[989] <= 32'b11111111110000010000000100010011;
ROM[990] <= 32'b00000000000000010010001110000011;
ROM[991] <= 32'b00000000000000111000001100010011;
ROM[992] <= 32'b00000000110100110000010000110011;
ROM[993] <= 32'b00000000000001000010001110000011;
ROM[994] <= 32'b00000000011100010010000000100011;
ROM[995] <= 32'b00000000010000010000000100010011;
ROM[996] <= 32'b00000100000000000000001110010011;
ROM[997] <= 32'b00000000011100010010000000100011;
ROM[998] <= 32'b00000000010000010000000100010011;
ROM[999] <= 32'b00000100000001101010001110000011;
ROM[1000] <= 32'b00000000011100010010000000100011;
ROM[1001] <= 32'b00000000010000010000000100010011;
ROM[1002] <= 32'b11111111110000010000000100010011;
ROM[1003] <= 32'b00000000000000010010001110000011;
ROM[1004] <= 32'b11111111110000010000000100010011;
ROM[1005] <= 32'b00000000000000010010010000000011;
ROM[1006] <= 32'b00000000011101000000001110110011;
ROM[1007] <= 32'b00000000011100010010000000100011;
ROM[1008] <= 32'b00000000010000010000000100010011;
ROM[1009] <= 32'b11111111110000010000000100010011;
ROM[1010] <= 32'b00000000000000010010001110000011;
ROM[1011] <= 32'b00000000000000111000001100010011;
ROM[1012] <= 32'b00000000110100110000010000110011;
ROM[1013] <= 32'b00000000000001000010001110000011;
ROM[1014] <= 32'b00000000011100010010000000100011;
ROM[1015] <= 32'b00000000010000010000000100010011;
ROM[1016] <= 32'b11111111110000010000000100010011;
ROM[1017] <= 32'b00000000000000010010001110000011;
ROM[1018] <= 32'b11111111110000010000000100010011;
ROM[1019] <= 32'b00000000000000010010010000000011;
ROM[1020] <= 32'b00000000011101000000001110110011;
ROM[1021] <= 32'b00000000011100010010000000100011;
ROM[1022] <= 32'b00000000010000010000000100010011;
ROM[1023] <= 32'b11111111110000010000000100010011;
ROM[1024] <= 32'b00000000000000010010001110000011;
ROM[1025] <= 32'b00000000011101100010000000100011;
ROM[1026] <= 32'b11111111110000010000000100010011;
ROM[1027] <= 32'b00000000000000010010001110000011;
ROM[1028] <= 32'b00000000000000111000001100010011;
ROM[1029] <= 32'b00000000000001100010001110000011;
ROM[1030] <= 32'b00000000011100010010000000100011;
ROM[1031] <= 32'b00000000010000010000000100010011;
ROM[1032] <= 32'b11111111110000010000000100010011;
ROM[1033] <= 32'b00000000000000010010001110000011;
ROM[1034] <= 32'b00000000110100110000010000110011;
ROM[1035] <= 32'b00000000011101000010000000100011;
ROM[1036] <= 32'b00000100100000000000001110010011;
ROM[1037] <= 32'b00000000011100010010000000100011;
ROM[1038] <= 32'b00000000010000010000000100010011;
ROM[1039] <= 32'b00000100000001101010001110000011;
ROM[1040] <= 32'b00000000011100010010000000100011;
ROM[1041] <= 32'b00000000010000010000000100010011;
ROM[1042] <= 32'b11111111110000010000000100010011;
ROM[1043] <= 32'b00000000000000010010001110000011;
ROM[1044] <= 32'b11111111110000010000000100010011;
ROM[1045] <= 32'b00000000000000010010010000000011;
ROM[1046] <= 32'b00000000011101000000001110110011;
ROM[1047] <= 32'b00000000011100010010000000100011;
ROM[1048] <= 32'b00000000010000010000000100010011;
ROM[1049] <= 32'b00000100010000000000001110010011;
ROM[1050] <= 32'b00000000011100010010000000100011;
ROM[1051] <= 32'b00000000010000010000000100010011;
ROM[1052] <= 32'b00000100000001101010001110000011;
ROM[1053] <= 32'b00000000011100010010000000100011;
ROM[1054] <= 32'b00000000010000010000000100010011;
ROM[1055] <= 32'b11111111110000010000000100010011;
ROM[1056] <= 32'b00000000000000010010001110000011;
ROM[1057] <= 32'b11111111110000010000000100010011;
ROM[1058] <= 32'b00000000000000010010010000000011;
ROM[1059] <= 32'b00000000011101000000001110110011;
ROM[1060] <= 32'b00000000011100010010000000100011;
ROM[1061] <= 32'b00000000010000010000000100010011;
ROM[1062] <= 32'b11111111110000010000000100010011;
ROM[1063] <= 32'b00000000000000010010001110000011;
ROM[1064] <= 32'b00000000000000111000001100010011;
ROM[1065] <= 32'b00000000110100110000010000110011;
ROM[1066] <= 32'b00000000000001000010001110000011;
ROM[1067] <= 32'b00000000011100010010000000100011;
ROM[1068] <= 32'b00000000010000010000000100010011;
ROM[1069] <= 32'b00000100010000000000001110010011;
ROM[1070] <= 32'b00000000011100010010000000100011;
ROM[1071] <= 32'b00000000010000010000000100010011;
ROM[1072] <= 32'b00000100000001101010001110000011;
ROM[1073] <= 32'b00000000011100010010000000100011;
ROM[1074] <= 32'b00000000010000010000000100010011;
ROM[1075] <= 32'b11111111110000010000000100010011;
ROM[1076] <= 32'b00000000000000010010001110000011;
ROM[1077] <= 32'b11111111110000010000000100010011;
ROM[1078] <= 32'b00000000000000010010010000000011;
ROM[1079] <= 32'b00000000011101000000001110110011;
ROM[1080] <= 32'b00000000011100010010000000100011;
ROM[1081] <= 32'b00000000010000010000000100010011;
ROM[1082] <= 32'b11111111110000010000000100010011;
ROM[1083] <= 32'b00000000000000010010001110000011;
ROM[1084] <= 32'b00000000000000111000001100010011;
ROM[1085] <= 32'b00000000110100110000010000110011;
ROM[1086] <= 32'b00000000000001000010001110000011;
ROM[1087] <= 32'b00000000011100010010000000100011;
ROM[1088] <= 32'b00000000010000010000000100010011;
ROM[1089] <= 32'b11111111110000010000000100010011;
ROM[1090] <= 32'b00000000000000010010001110000011;
ROM[1091] <= 32'b11111111110000010000000100010011;
ROM[1092] <= 32'b00000000000000010010010000000011;
ROM[1093] <= 32'b00000000011101000000001110110011;
ROM[1094] <= 32'b00000000011100010010000000100011;
ROM[1095] <= 32'b00000000010000010000000100010011;
ROM[1096] <= 32'b11111111110000010000000100010011;
ROM[1097] <= 32'b00000000000000010010001110000011;
ROM[1098] <= 32'b00000000011101100010000000100011;
ROM[1099] <= 32'b11111111110000010000000100010011;
ROM[1100] <= 32'b00000000000000010010001110000011;
ROM[1101] <= 32'b00000000000000111000001100010011;
ROM[1102] <= 32'b00000000000001100010001110000011;
ROM[1103] <= 32'b00000000011100010010000000100011;
ROM[1104] <= 32'b00000000010000010000000100010011;
ROM[1105] <= 32'b11111111110000010000000100010011;
ROM[1106] <= 32'b00000000000000010010001110000011;
ROM[1107] <= 32'b00000000110100110000010000110011;
ROM[1108] <= 32'b00000000011101000010000000100011;
ROM[1109] <= 32'b00000100110000000000001110010011;
ROM[1110] <= 32'b00000000011100010010000000100011;
ROM[1111] <= 32'b00000000010000010000000100010011;
ROM[1112] <= 32'b00000100000001101010001110000011;
ROM[1113] <= 32'b00000000011100010010000000100011;
ROM[1114] <= 32'b00000000010000010000000100010011;
ROM[1115] <= 32'b11111111110000010000000100010011;
ROM[1116] <= 32'b00000000000000010010001110000011;
ROM[1117] <= 32'b11111111110000010000000100010011;
ROM[1118] <= 32'b00000000000000010010010000000011;
ROM[1119] <= 32'b00000000011101000000001110110011;
ROM[1120] <= 32'b00000000011100010010000000100011;
ROM[1121] <= 32'b00000000010000010000000100010011;
ROM[1122] <= 32'b00000100100000000000001110010011;
ROM[1123] <= 32'b00000000011100010010000000100011;
ROM[1124] <= 32'b00000000010000010000000100010011;
ROM[1125] <= 32'b00000100000001101010001110000011;
ROM[1126] <= 32'b00000000011100010010000000100011;
ROM[1127] <= 32'b00000000010000010000000100010011;
ROM[1128] <= 32'b11111111110000010000000100010011;
ROM[1129] <= 32'b00000000000000010010001110000011;
ROM[1130] <= 32'b11111111110000010000000100010011;
ROM[1131] <= 32'b00000000000000010010010000000011;
ROM[1132] <= 32'b00000000011101000000001110110011;
ROM[1133] <= 32'b00000000011100010010000000100011;
ROM[1134] <= 32'b00000000010000010000000100010011;
ROM[1135] <= 32'b11111111110000010000000100010011;
ROM[1136] <= 32'b00000000000000010010001110000011;
ROM[1137] <= 32'b00000000000000111000001100010011;
ROM[1138] <= 32'b00000000110100110000010000110011;
ROM[1139] <= 32'b00000000000001000010001110000011;
ROM[1140] <= 32'b00000000011100010010000000100011;
ROM[1141] <= 32'b00000000010000010000000100010011;
ROM[1142] <= 32'b00000100100000000000001110010011;
ROM[1143] <= 32'b00000000011100010010000000100011;
ROM[1144] <= 32'b00000000010000010000000100010011;
ROM[1145] <= 32'b00000100000001101010001110000011;
ROM[1146] <= 32'b00000000011100010010000000100011;
ROM[1147] <= 32'b00000000010000010000000100010011;
ROM[1148] <= 32'b11111111110000010000000100010011;
ROM[1149] <= 32'b00000000000000010010001110000011;
ROM[1150] <= 32'b11111111110000010000000100010011;
ROM[1151] <= 32'b00000000000000010010010000000011;
ROM[1152] <= 32'b00000000011101000000001110110011;
ROM[1153] <= 32'b00000000011100010010000000100011;
ROM[1154] <= 32'b00000000010000010000000100010011;
ROM[1155] <= 32'b11111111110000010000000100010011;
ROM[1156] <= 32'b00000000000000010010001110000011;
ROM[1157] <= 32'b00000000000000111000001100010011;
ROM[1158] <= 32'b00000000110100110000010000110011;
ROM[1159] <= 32'b00000000000001000010001110000011;
ROM[1160] <= 32'b00000000011100010010000000100011;
ROM[1161] <= 32'b00000000010000010000000100010011;
ROM[1162] <= 32'b11111111110000010000000100010011;
ROM[1163] <= 32'b00000000000000010010001110000011;
ROM[1164] <= 32'b11111111110000010000000100010011;
ROM[1165] <= 32'b00000000000000010010010000000011;
ROM[1166] <= 32'b00000000011101000000001110110011;
ROM[1167] <= 32'b00000000011100010010000000100011;
ROM[1168] <= 32'b00000000010000010000000100010011;
ROM[1169] <= 32'b11111111110000010000000100010011;
ROM[1170] <= 32'b00000000000000010010001110000011;
ROM[1171] <= 32'b00000000011101100010000000100011;
ROM[1172] <= 32'b11111111110000010000000100010011;
ROM[1173] <= 32'b00000000000000010010001110000011;
ROM[1174] <= 32'b00000000000000111000001100010011;
ROM[1175] <= 32'b00000000000001100010001110000011;
ROM[1176] <= 32'b00000000011100010010000000100011;
ROM[1177] <= 32'b00000000010000010000000100010011;
ROM[1178] <= 32'b11111111110000010000000100010011;
ROM[1179] <= 32'b00000000000000010010001110000011;
ROM[1180] <= 32'b00000000110100110000010000110011;
ROM[1181] <= 32'b00000000011101000010000000100011;
ROM[1182] <= 32'b00000101000000000000001110010011;
ROM[1183] <= 32'b00000000011100010010000000100011;
ROM[1184] <= 32'b00000000010000010000000100010011;
ROM[1185] <= 32'b00000100000001101010001110000011;
ROM[1186] <= 32'b00000000011100010010000000100011;
ROM[1187] <= 32'b00000000010000010000000100010011;
ROM[1188] <= 32'b11111111110000010000000100010011;
ROM[1189] <= 32'b00000000000000010010001110000011;
ROM[1190] <= 32'b11111111110000010000000100010011;
ROM[1191] <= 32'b00000000000000010010010000000011;
ROM[1192] <= 32'b00000000011101000000001110110011;
ROM[1193] <= 32'b00000000011100010010000000100011;
ROM[1194] <= 32'b00000000010000010000000100010011;
ROM[1195] <= 32'b00000100110000000000001110010011;
ROM[1196] <= 32'b00000000011100010010000000100011;
ROM[1197] <= 32'b00000000010000010000000100010011;
ROM[1198] <= 32'b00000100000001101010001110000011;
ROM[1199] <= 32'b00000000011100010010000000100011;
ROM[1200] <= 32'b00000000010000010000000100010011;
ROM[1201] <= 32'b11111111110000010000000100010011;
ROM[1202] <= 32'b00000000000000010010001110000011;
ROM[1203] <= 32'b11111111110000010000000100010011;
ROM[1204] <= 32'b00000000000000010010010000000011;
ROM[1205] <= 32'b00000000011101000000001110110011;
ROM[1206] <= 32'b00000000011100010010000000100011;
ROM[1207] <= 32'b00000000010000010000000100010011;
ROM[1208] <= 32'b11111111110000010000000100010011;
ROM[1209] <= 32'b00000000000000010010001110000011;
ROM[1210] <= 32'b00000000000000111000001100010011;
ROM[1211] <= 32'b00000000110100110000010000110011;
ROM[1212] <= 32'b00000000000001000010001110000011;
ROM[1213] <= 32'b00000000011100010010000000100011;
ROM[1214] <= 32'b00000000010000010000000100010011;
ROM[1215] <= 32'b00000100110000000000001110010011;
ROM[1216] <= 32'b00000000011100010010000000100011;
ROM[1217] <= 32'b00000000010000010000000100010011;
ROM[1218] <= 32'b00000100000001101010001110000011;
ROM[1219] <= 32'b00000000011100010010000000100011;
ROM[1220] <= 32'b00000000010000010000000100010011;
ROM[1221] <= 32'b11111111110000010000000100010011;
ROM[1222] <= 32'b00000000000000010010001110000011;
ROM[1223] <= 32'b11111111110000010000000100010011;
ROM[1224] <= 32'b00000000000000010010010000000011;
ROM[1225] <= 32'b00000000011101000000001110110011;
ROM[1226] <= 32'b00000000011100010010000000100011;
ROM[1227] <= 32'b00000000010000010000000100010011;
ROM[1228] <= 32'b11111111110000010000000100010011;
ROM[1229] <= 32'b00000000000000010010001110000011;
ROM[1230] <= 32'b00000000000000111000001100010011;
ROM[1231] <= 32'b00000000110100110000010000110011;
ROM[1232] <= 32'b00000000000001000010001110000011;
ROM[1233] <= 32'b00000000011100010010000000100011;
ROM[1234] <= 32'b00000000010000010000000100010011;
ROM[1235] <= 32'b11111111110000010000000100010011;
ROM[1236] <= 32'b00000000000000010010001110000011;
ROM[1237] <= 32'b11111111110000010000000100010011;
ROM[1238] <= 32'b00000000000000010010010000000011;
ROM[1239] <= 32'b00000000011101000000001110110011;
ROM[1240] <= 32'b00000000011100010010000000100011;
ROM[1241] <= 32'b00000000010000010000000100010011;
ROM[1242] <= 32'b11111111110000010000000100010011;
ROM[1243] <= 32'b00000000000000010010001110000011;
ROM[1244] <= 32'b00000000011101100010000000100011;
ROM[1245] <= 32'b11111111110000010000000100010011;
ROM[1246] <= 32'b00000000000000010010001110000011;
ROM[1247] <= 32'b00000000000000111000001100010011;
ROM[1248] <= 32'b00000000000001100010001110000011;
ROM[1249] <= 32'b00000000011100010010000000100011;
ROM[1250] <= 32'b00000000010000010000000100010011;
ROM[1251] <= 32'b11111111110000010000000100010011;
ROM[1252] <= 32'b00000000000000010010001110000011;
ROM[1253] <= 32'b00000000110100110000010000110011;
ROM[1254] <= 32'b00000000011101000010000000100011;
ROM[1255] <= 32'b00000101010000000000001110010011;
ROM[1256] <= 32'b00000000011100010010000000100011;
ROM[1257] <= 32'b00000000010000010000000100010011;
ROM[1258] <= 32'b00000100000001101010001110000011;
ROM[1259] <= 32'b00000000011100010010000000100011;
ROM[1260] <= 32'b00000000010000010000000100010011;
ROM[1261] <= 32'b11111111110000010000000100010011;
ROM[1262] <= 32'b00000000000000010010001110000011;
ROM[1263] <= 32'b11111111110000010000000100010011;
ROM[1264] <= 32'b00000000000000010010010000000011;
ROM[1265] <= 32'b00000000011101000000001110110011;
ROM[1266] <= 32'b00000000011100010010000000100011;
ROM[1267] <= 32'b00000000010000010000000100010011;
ROM[1268] <= 32'b00000101000000000000001110010011;
ROM[1269] <= 32'b00000000011100010010000000100011;
ROM[1270] <= 32'b00000000010000010000000100010011;
ROM[1271] <= 32'b00000100000001101010001110000011;
ROM[1272] <= 32'b00000000011100010010000000100011;
ROM[1273] <= 32'b00000000010000010000000100010011;
ROM[1274] <= 32'b11111111110000010000000100010011;
ROM[1275] <= 32'b00000000000000010010001110000011;
ROM[1276] <= 32'b11111111110000010000000100010011;
ROM[1277] <= 32'b00000000000000010010010000000011;
ROM[1278] <= 32'b00000000011101000000001110110011;
ROM[1279] <= 32'b00000000011100010010000000100011;
ROM[1280] <= 32'b00000000010000010000000100010011;
ROM[1281] <= 32'b11111111110000010000000100010011;
ROM[1282] <= 32'b00000000000000010010001110000011;
ROM[1283] <= 32'b00000000000000111000001100010011;
ROM[1284] <= 32'b00000000110100110000010000110011;
ROM[1285] <= 32'b00000000000001000010001110000011;
ROM[1286] <= 32'b00000000011100010010000000100011;
ROM[1287] <= 32'b00000000010000010000000100010011;
ROM[1288] <= 32'b00000101000000000000001110010011;
ROM[1289] <= 32'b00000000011100010010000000100011;
ROM[1290] <= 32'b00000000010000010000000100010011;
ROM[1291] <= 32'b00000100000001101010001110000011;
ROM[1292] <= 32'b00000000011100010010000000100011;
ROM[1293] <= 32'b00000000010000010000000100010011;
ROM[1294] <= 32'b11111111110000010000000100010011;
ROM[1295] <= 32'b00000000000000010010001110000011;
ROM[1296] <= 32'b11111111110000010000000100010011;
ROM[1297] <= 32'b00000000000000010010010000000011;
ROM[1298] <= 32'b00000000011101000000001110110011;
ROM[1299] <= 32'b00000000011100010010000000100011;
ROM[1300] <= 32'b00000000010000010000000100010011;
ROM[1301] <= 32'b11111111110000010000000100010011;
ROM[1302] <= 32'b00000000000000010010001110000011;
ROM[1303] <= 32'b00000000000000111000001100010011;
ROM[1304] <= 32'b00000000110100110000010000110011;
ROM[1305] <= 32'b00000000000001000010001110000011;
ROM[1306] <= 32'b00000000011100010010000000100011;
ROM[1307] <= 32'b00000000010000010000000100010011;
ROM[1308] <= 32'b11111111110000010000000100010011;
ROM[1309] <= 32'b00000000000000010010001110000011;
ROM[1310] <= 32'b11111111110000010000000100010011;
ROM[1311] <= 32'b00000000000000010010010000000011;
ROM[1312] <= 32'b00000000011101000000001110110011;
ROM[1313] <= 32'b00000000011100010010000000100011;
ROM[1314] <= 32'b00000000010000010000000100010011;
ROM[1315] <= 32'b11111111110000010000000100010011;
ROM[1316] <= 32'b00000000000000010010001110000011;
ROM[1317] <= 32'b00000000011101100010000000100011;
ROM[1318] <= 32'b11111111110000010000000100010011;
ROM[1319] <= 32'b00000000000000010010001110000011;
ROM[1320] <= 32'b00000000000000111000001100010011;
ROM[1321] <= 32'b00000000000001100010001110000011;
ROM[1322] <= 32'b00000000011100010010000000100011;
ROM[1323] <= 32'b00000000010000010000000100010011;
ROM[1324] <= 32'b11111111110000010000000100010011;
ROM[1325] <= 32'b00000000000000010010001110000011;
ROM[1326] <= 32'b00000000110100110000010000110011;
ROM[1327] <= 32'b00000000011101000010000000100011;
ROM[1328] <= 32'b00000101100000000000001110010011;
ROM[1329] <= 32'b00000000011100010010000000100011;
ROM[1330] <= 32'b00000000010000010000000100010011;
ROM[1331] <= 32'b00000100000001101010001110000011;
ROM[1332] <= 32'b00000000011100010010000000100011;
ROM[1333] <= 32'b00000000010000010000000100010011;
ROM[1334] <= 32'b11111111110000010000000100010011;
ROM[1335] <= 32'b00000000000000010010001110000011;
ROM[1336] <= 32'b11111111110000010000000100010011;
ROM[1337] <= 32'b00000000000000010010010000000011;
ROM[1338] <= 32'b00000000011101000000001110110011;
ROM[1339] <= 32'b00000000011100010010000000100011;
ROM[1340] <= 32'b00000000010000010000000100010011;
ROM[1341] <= 32'b00000101010000000000001110010011;
ROM[1342] <= 32'b00000000011100010010000000100011;
ROM[1343] <= 32'b00000000010000010000000100010011;
ROM[1344] <= 32'b00000100000001101010001110000011;
ROM[1345] <= 32'b00000000011100010010000000100011;
ROM[1346] <= 32'b00000000010000010000000100010011;
ROM[1347] <= 32'b11111111110000010000000100010011;
ROM[1348] <= 32'b00000000000000010010001110000011;
ROM[1349] <= 32'b11111111110000010000000100010011;
ROM[1350] <= 32'b00000000000000010010010000000011;
ROM[1351] <= 32'b00000000011101000000001110110011;
ROM[1352] <= 32'b00000000011100010010000000100011;
ROM[1353] <= 32'b00000000010000010000000100010011;
ROM[1354] <= 32'b11111111110000010000000100010011;
ROM[1355] <= 32'b00000000000000010010001110000011;
ROM[1356] <= 32'b00000000000000111000001100010011;
ROM[1357] <= 32'b00000000110100110000010000110011;
ROM[1358] <= 32'b00000000000001000010001110000011;
ROM[1359] <= 32'b00000000011100010010000000100011;
ROM[1360] <= 32'b00000000010000010000000100010011;
ROM[1361] <= 32'b00000101010000000000001110010011;
ROM[1362] <= 32'b00000000011100010010000000100011;
ROM[1363] <= 32'b00000000010000010000000100010011;
ROM[1364] <= 32'b00000100000001101010001110000011;
ROM[1365] <= 32'b00000000011100010010000000100011;
ROM[1366] <= 32'b00000000010000010000000100010011;
ROM[1367] <= 32'b11111111110000010000000100010011;
ROM[1368] <= 32'b00000000000000010010001110000011;
ROM[1369] <= 32'b11111111110000010000000100010011;
ROM[1370] <= 32'b00000000000000010010010000000011;
ROM[1371] <= 32'b00000000011101000000001110110011;
ROM[1372] <= 32'b00000000011100010010000000100011;
ROM[1373] <= 32'b00000000010000010000000100010011;
ROM[1374] <= 32'b11111111110000010000000100010011;
ROM[1375] <= 32'b00000000000000010010001110000011;
ROM[1376] <= 32'b00000000000000111000001100010011;
ROM[1377] <= 32'b00000000110100110000010000110011;
ROM[1378] <= 32'b00000000000001000010001110000011;
ROM[1379] <= 32'b00000000011100010010000000100011;
ROM[1380] <= 32'b00000000010000010000000100010011;
ROM[1381] <= 32'b11111111110000010000000100010011;
ROM[1382] <= 32'b00000000000000010010001110000011;
ROM[1383] <= 32'b11111111110000010000000100010011;
ROM[1384] <= 32'b00000000000000010010010000000011;
ROM[1385] <= 32'b00000000011101000000001110110011;
ROM[1386] <= 32'b00000000011100010010000000100011;
ROM[1387] <= 32'b00000000010000010000000100010011;
ROM[1388] <= 32'b11111111110000010000000100010011;
ROM[1389] <= 32'b00000000000000010010001110000011;
ROM[1390] <= 32'b00000000011101100010000000100011;
ROM[1391] <= 32'b11111111110000010000000100010011;
ROM[1392] <= 32'b00000000000000010010001110000011;
ROM[1393] <= 32'b00000000000000111000001100010011;
ROM[1394] <= 32'b00000000000001100010001110000011;
ROM[1395] <= 32'b00000000011100010010000000100011;
ROM[1396] <= 32'b00000000010000010000000100010011;
ROM[1397] <= 32'b11111111110000010000000100010011;
ROM[1398] <= 32'b00000000000000010010001110000011;
ROM[1399] <= 32'b00000000110100110000010000110011;
ROM[1400] <= 32'b00000000011101000010000000100011;
ROM[1401] <= 32'b00000101110000000000001110010011;
ROM[1402] <= 32'b00000000011100010010000000100011;
ROM[1403] <= 32'b00000000010000010000000100010011;
ROM[1404] <= 32'b00000100000001101010001110000011;
ROM[1405] <= 32'b00000000011100010010000000100011;
ROM[1406] <= 32'b00000000010000010000000100010011;
ROM[1407] <= 32'b11111111110000010000000100010011;
ROM[1408] <= 32'b00000000000000010010001110000011;
ROM[1409] <= 32'b11111111110000010000000100010011;
ROM[1410] <= 32'b00000000000000010010010000000011;
ROM[1411] <= 32'b00000000011101000000001110110011;
ROM[1412] <= 32'b00000000011100010010000000100011;
ROM[1413] <= 32'b00000000010000010000000100010011;
ROM[1414] <= 32'b00000101100000000000001110010011;
ROM[1415] <= 32'b00000000011100010010000000100011;
ROM[1416] <= 32'b00000000010000010000000100010011;
ROM[1417] <= 32'b00000100000001101010001110000011;
ROM[1418] <= 32'b00000000011100010010000000100011;
ROM[1419] <= 32'b00000000010000010000000100010011;
ROM[1420] <= 32'b11111111110000010000000100010011;
ROM[1421] <= 32'b00000000000000010010001110000011;
ROM[1422] <= 32'b11111111110000010000000100010011;
ROM[1423] <= 32'b00000000000000010010010000000011;
ROM[1424] <= 32'b00000000011101000000001110110011;
ROM[1425] <= 32'b00000000011100010010000000100011;
ROM[1426] <= 32'b00000000010000010000000100010011;
ROM[1427] <= 32'b11111111110000010000000100010011;
ROM[1428] <= 32'b00000000000000010010001110000011;
ROM[1429] <= 32'b00000000000000111000001100010011;
ROM[1430] <= 32'b00000000110100110000010000110011;
ROM[1431] <= 32'b00000000000001000010001110000011;
ROM[1432] <= 32'b00000000011100010010000000100011;
ROM[1433] <= 32'b00000000010000010000000100010011;
ROM[1434] <= 32'b00000101100000000000001110010011;
ROM[1435] <= 32'b00000000011100010010000000100011;
ROM[1436] <= 32'b00000000010000010000000100010011;
ROM[1437] <= 32'b00000100000001101010001110000011;
ROM[1438] <= 32'b00000000011100010010000000100011;
ROM[1439] <= 32'b00000000010000010000000100010011;
ROM[1440] <= 32'b11111111110000010000000100010011;
ROM[1441] <= 32'b00000000000000010010001110000011;
ROM[1442] <= 32'b11111111110000010000000100010011;
ROM[1443] <= 32'b00000000000000010010010000000011;
ROM[1444] <= 32'b00000000011101000000001110110011;
ROM[1445] <= 32'b00000000011100010010000000100011;
ROM[1446] <= 32'b00000000010000010000000100010011;
ROM[1447] <= 32'b11111111110000010000000100010011;
ROM[1448] <= 32'b00000000000000010010001110000011;
ROM[1449] <= 32'b00000000000000111000001100010011;
ROM[1450] <= 32'b00000000110100110000010000110011;
ROM[1451] <= 32'b00000000000001000010001110000011;
ROM[1452] <= 32'b00000000011100010010000000100011;
ROM[1453] <= 32'b00000000010000010000000100010011;
ROM[1454] <= 32'b11111111110000010000000100010011;
ROM[1455] <= 32'b00000000000000010010001110000011;
ROM[1456] <= 32'b11111111110000010000000100010011;
ROM[1457] <= 32'b00000000000000010010010000000011;
ROM[1458] <= 32'b00000000011101000000001110110011;
ROM[1459] <= 32'b00000000011100010010000000100011;
ROM[1460] <= 32'b00000000010000010000000100010011;
ROM[1461] <= 32'b11111111110000010000000100010011;
ROM[1462] <= 32'b00000000000000010010001110000011;
ROM[1463] <= 32'b00000000011101100010000000100011;
ROM[1464] <= 32'b11111111110000010000000100010011;
ROM[1465] <= 32'b00000000000000010010001110000011;
ROM[1466] <= 32'b00000000000000111000001100010011;
ROM[1467] <= 32'b00000000000001100010001110000011;
ROM[1468] <= 32'b00000000011100010010000000100011;
ROM[1469] <= 32'b00000000010000010000000100010011;
ROM[1470] <= 32'b11111111110000010000000100010011;
ROM[1471] <= 32'b00000000000000010010001110000011;
ROM[1472] <= 32'b00000000110100110000010000110011;
ROM[1473] <= 32'b00000000011101000010000000100011;
ROM[1474] <= 32'b00000110000000000000001110010011;
ROM[1475] <= 32'b00000000011100010010000000100011;
ROM[1476] <= 32'b00000000010000010000000100010011;
ROM[1477] <= 32'b00000100000001101010001110000011;
ROM[1478] <= 32'b00000000011100010010000000100011;
ROM[1479] <= 32'b00000000010000010000000100010011;
ROM[1480] <= 32'b11111111110000010000000100010011;
ROM[1481] <= 32'b00000000000000010010001110000011;
ROM[1482] <= 32'b11111111110000010000000100010011;
ROM[1483] <= 32'b00000000000000010010010000000011;
ROM[1484] <= 32'b00000000011101000000001110110011;
ROM[1485] <= 32'b00000000011100010010000000100011;
ROM[1486] <= 32'b00000000010000010000000100010011;
ROM[1487] <= 32'b00000101110000000000001110010011;
ROM[1488] <= 32'b00000000011100010010000000100011;
ROM[1489] <= 32'b00000000010000010000000100010011;
ROM[1490] <= 32'b00000100000001101010001110000011;
ROM[1491] <= 32'b00000000011100010010000000100011;
ROM[1492] <= 32'b00000000010000010000000100010011;
ROM[1493] <= 32'b11111111110000010000000100010011;
ROM[1494] <= 32'b00000000000000010010001110000011;
ROM[1495] <= 32'b11111111110000010000000100010011;
ROM[1496] <= 32'b00000000000000010010010000000011;
ROM[1497] <= 32'b00000000011101000000001110110011;
ROM[1498] <= 32'b00000000011100010010000000100011;
ROM[1499] <= 32'b00000000010000010000000100010011;
ROM[1500] <= 32'b11111111110000010000000100010011;
ROM[1501] <= 32'b00000000000000010010001110000011;
ROM[1502] <= 32'b00000000000000111000001100010011;
ROM[1503] <= 32'b00000000110100110000010000110011;
ROM[1504] <= 32'b00000000000001000010001110000011;
ROM[1505] <= 32'b00000000011100010010000000100011;
ROM[1506] <= 32'b00000000010000010000000100010011;
ROM[1507] <= 32'b00000101110000000000001110010011;
ROM[1508] <= 32'b00000000011100010010000000100011;
ROM[1509] <= 32'b00000000010000010000000100010011;
ROM[1510] <= 32'b00000100000001101010001110000011;
ROM[1511] <= 32'b00000000011100010010000000100011;
ROM[1512] <= 32'b00000000010000010000000100010011;
ROM[1513] <= 32'b11111111110000010000000100010011;
ROM[1514] <= 32'b00000000000000010010001110000011;
ROM[1515] <= 32'b11111111110000010000000100010011;
ROM[1516] <= 32'b00000000000000010010010000000011;
ROM[1517] <= 32'b00000000011101000000001110110011;
ROM[1518] <= 32'b00000000011100010010000000100011;
ROM[1519] <= 32'b00000000010000010000000100010011;
ROM[1520] <= 32'b11111111110000010000000100010011;
ROM[1521] <= 32'b00000000000000010010001110000011;
ROM[1522] <= 32'b00000000000000111000001100010011;
ROM[1523] <= 32'b00000000110100110000010000110011;
ROM[1524] <= 32'b00000000000001000010001110000011;
ROM[1525] <= 32'b00000000011100010010000000100011;
ROM[1526] <= 32'b00000000010000010000000100010011;
ROM[1527] <= 32'b11111111110000010000000100010011;
ROM[1528] <= 32'b00000000000000010010001110000011;
ROM[1529] <= 32'b11111111110000010000000100010011;
ROM[1530] <= 32'b00000000000000010010010000000011;
ROM[1531] <= 32'b00000000011101000000001110110011;
ROM[1532] <= 32'b00000000011100010010000000100011;
ROM[1533] <= 32'b00000000010000010000000100010011;
ROM[1534] <= 32'b11111111110000010000000100010011;
ROM[1535] <= 32'b00000000000000010010001110000011;
ROM[1536] <= 32'b00000000011101100010000000100011;
ROM[1537] <= 32'b11111111110000010000000100010011;
ROM[1538] <= 32'b00000000000000010010001110000011;
ROM[1539] <= 32'b00000000000000111000001100010011;
ROM[1540] <= 32'b00000000000001100010001110000011;
ROM[1541] <= 32'b00000000011100010010000000100011;
ROM[1542] <= 32'b00000000010000010000000100010011;
ROM[1543] <= 32'b11111111110000010000000100010011;
ROM[1544] <= 32'b00000000000000010010001110000011;
ROM[1545] <= 32'b00000000110100110000010000110011;
ROM[1546] <= 32'b00000000011101000010000000100011;
ROM[1547] <= 32'b00000110010000000000001110010011;
ROM[1548] <= 32'b00000000011100010010000000100011;
ROM[1549] <= 32'b00000000010000010000000100010011;
ROM[1550] <= 32'b00000100000001101010001110000011;
ROM[1551] <= 32'b00000000011100010010000000100011;
ROM[1552] <= 32'b00000000010000010000000100010011;
ROM[1553] <= 32'b11111111110000010000000100010011;
ROM[1554] <= 32'b00000000000000010010001110000011;
ROM[1555] <= 32'b11111111110000010000000100010011;
ROM[1556] <= 32'b00000000000000010010010000000011;
ROM[1557] <= 32'b00000000011101000000001110110011;
ROM[1558] <= 32'b00000000011100010010000000100011;
ROM[1559] <= 32'b00000000010000010000000100010011;
ROM[1560] <= 32'b00000110000000000000001110010011;
ROM[1561] <= 32'b00000000011100010010000000100011;
ROM[1562] <= 32'b00000000010000010000000100010011;
ROM[1563] <= 32'b00000100000001101010001110000011;
ROM[1564] <= 32'b00000000011100010010000000100011;
ROM[1565] <= 32'b00000000010000010000000100010011;
ROM[1566] <= 32'b11111111110000010000000100010011;
ROM[1567] <= 32'b00000000000000010010001110000011;
ROM[1568] <= 32'b11111111110000010000000100010011;
ROM[1569] <= 32'b00000000000000010010010000000011;
ROM[1570] <= 32'b00000000011101000000001110110011;
ROM[1571] <= 32'b00000000011100010010000000100011;
ROM[1572] <= 32'b00000000010000010000000100010011;
ROM[1573] <= 32'b11111111110000010000000100010011;
ROM[1574] <= 32'b00000000000000010010001110000011;
ROM[1575] <= 32'b00000000000000111000001100010011;
ROM[1576] <= 32'b00000000110100110000010000110011;
ROM[1577] <= 32'b00000000000001000010001110000011;
ROM[1578] <= 32'b00000000011100010010000000100011;
ROM[1579] <= 32'b00000000010000010000000100010011;
ROM[1580] <= 32'b00000110000000000000001110010011;
ROM[1581] <= 32'b00000000011100010010000000100011;
ROM[1582] <= 32'b00000000010000010000000100010011;
ROM[1583] <= 32'b00000100000001101010001110000011;
ROM[1584] <= 32'b00000000011100010010000000100011;
ROM[1585] <= 32'b00000000010000010000000100010011;
ROM[1586] <= 32'b11111111110000010000000100010011;
ROM[1587] <= 32'b00000000000000010010001110000011;
ROM[1588] <= 32'b11111111110000010000000100010011;
ROM[1589] <= 32'b00000000000000010010010000000011;
ROM[1590] <= 32'b00000000011101000000001110110011;
ROM[1591] <= 32'b00000000011100010010000000100011;
ROM[1592] <= 32'b00000000010000010000000100010011;
ROM[1593] <= 32'b11111111110000010000000100010011;
ROM[1594] <= 32'b00000000000000010010001110000011;
ROM[1595] <= 32'b00000000000000111000001100010011;
ROM[1596] <= 32'b00000000110100110000010000110011;
ROM[1597] <= 32'b00000000000001000010001110000011;
ROM[1598] <= 32'b00000000011100010010000000100011;
ROM[1599] <= 32'b00000000010000010000000100010011;
ROM[1600] <= 32'b11111111110000010000000100010011;
ROM[1601] <= 32'b00000000000000010010001110000011;
ROM[1602] <= 32'b11111111110000010000000100010011;
ROM[1603] <= 32'b00000000000000010010010000000011;
ROM[1604] <= 32'b00000000011101000000001110110011;
ROM[1605] <= 32'b00000000011100010010000000100011;
ROM[1606] <= 32'b00000000010000010000000100010011;
ROM[1607] <= 32'b11111111110000010000000100010011;
ROM[1608] <= 32'b00000000000000010010001110000011;
ROM[1609] <= 32'b00000000011101100010000000100011;
ROM[1610] <= 32'b11111111110000010000000100010011;
ROM[1611] <= 32'b00000000000000010010001110000011;
ROM[1612] <= 32'b00000000000000111000001100010011;
ROM[1613] <= 32'b00000000000001100010001110000011;
ROM[1614] <= 32'b00000000011100010010000000100011;
ROM[1615] <= 32'b00000000010000010000000100010011;
ROM[1616] <= 32'b11111111110000010000000100010011;
ROM[1617] <= 32'b00000000000000010010001110000011;
ROM[1618] <= 32'b00000000110100110000010000110011;
ROM[1619] <= 32'b00000000011101000010000000100011;
ROM[1620] <= 32'b00000110100000000000001110010011;
ROM[1621] <= 32'b00000000011100010010000000100011;
ROM[1622] <= 32'b00000000010000010000000100010011;
ROM[1623] <= 32'b00000100000001101010001110000011;
ROM[1624] <= 32'b00000000011100010010000000100011;
ROM[1625] <= 32'b00000000010000010000000100010011;
ROM[1626] <= 32'b11111111110000010000000100010011;
ROM[1627] <= 32'b00000000000000010010001110000011;
ROM[1628] <= 32'b11111111110000010000000100010011;
ROM[1629] <= 32'b00000000000000010010010000000011;
ROM[1630] <= 32'b00000000011101000000001110110011;
ROM[1631] <= 32'b00000000011100010010000000100011;
ROM[1632] <= 32'b00000000010000010000000100010011;
ROM[1633] <= 32'b00000110010000000000001110010011;
ROM[1634] <= 32'b00000000011100010010000000100011;
ROM[1635] <= 32'b00000000010000010000000100010011;
ROM[1636] <= 32'b00000100000001101010001110000011;
ROM[1637] <= 32'b00000000011100010010000000100011;
ROM[1638] <= 32'b00000000010000010000000100010011;
ROM[1639] <= 32'b11111111110000010000000100010011;
ROM[1640] <= 32'b00000000000000010010001110000011;
ROM[1641] <= 32'b11111111110000010000000100010011;
ROM[1642] <= 32'b00000000000000010010010000000011;
ROM[1643] <= 32'b00000000011101000000001110110011;
ROM[1644] <= 32'b00000000011100010010000000100011;
ROM[1645] <= 32'b00000000010000010000000100010011;
ROM[1646] <= 32'b11111111110000010000000100010011;
ROM[1647] <= 32'b00000000000000010010001110000011;
ROM[1648] <= 32'b00000000000000111000001100010011;
ROM[1649] <= 32'b00000000110100110000010000110011;
ROM[1650] <= 32'b00000000000001000010001110000011;
ROM[1651] <= 32'b00000000011100010010000000100011;
ROM[1652] <= 32'b00000000010000010000000100010011;
ROM[1653] <= 32'b00000110010000000000001110010011;
ROM[1654] <= 32'b00000000011100010010000000100011;
ROM[1655] <= 32'b00000000010000010000000100010011;
ROM[1656] <= 32'b00000100000001101010001110000011;
ROM[1657] <= 32'b00000000011100010010000000100011;
ROM[1658] <= 32'b00000000010000010000000100010011;
ROM[1659] <= 32'b11111111110000010000000100010011;
ROM[1660] <= 32'b00000000000000010010001110000011;
ROM[1661] <= 32'b11111111110000010000000100010011;
ROM[1662] <= 32'b00000000000000010010010000000011;
ROM[1663] <= 32'b00000000011101000000001110110011;
ROM[1664] <= 32'b00000000011100010010000000100011;
ROM[1665] <= 32'b00000000010000010000000100010011;
ROM[1666] <= 32'b11111111110000010000000100010011;
ROM[1667] <= 32'b00000000000000010010001110000011;
ROM[1668] <= 32'b00000000000000111000001100010011;
ROM[1669] <= 32'b00000000110100110000010000110011;
ROM[1670] <= 32'b00000000000001000010001110000011;
ROM[1671] <= 32'b00000000011100010010000000100011;
ROM[1672] <= 32'b00000000010000010000000100010011;
ROM[1673] <= 32'b11111111110000010000000100010011;
ROM[1674] <= 32'b00000000000000010010001110000011;
ROM[1675] <= 32'b11111111110000010000000100010011;
ROM[1676] <= 32'b00000000000000010010010000000011;
ROM[1677] <= 32'b00000000011101000000001110110011;
ROM[1678] <= 32'b00000000011100010010000000100011;
ROM[1679] <= 32'b00000000010000010000000100010011;
ROM[1680] <= 32'b11111111110000010000000100010011;
ROM[1681] <= 32'b00000000000000010010001110000011;
ROM[1682] <= 32'b00000000011101100010000000100011;
ROM[1683] <= 32'b11111111110000010000000100010011;
ROM[1684] <= 32'b00000000000000010010001110000011;
ROM[1685] <= 32'b00000000000000111000001100010011;
ROM[1686] <= 32'b00000000000001100010001110000011;
ROM[1687] <= 32'b00000000011100010010000000100011;
ROM[1688] <= 32'b00000000010000010000000100010011;
ROM[1689] <= 32'b11111111110000010000000100010011;
ROM[1690] <= 32'b00000000000000010010001110000011;
ROM[1691] <= 32'b00000000110100110000010000110011;
ROM[1692] <= 32'b00000000011101000010000000100011;
ROM[1693] <= 32'b00000110110000000000001110010011;
ROM[1694] <= 32'b00000000011100010010000000100011;
ROM[1695] <= 32'b00000000010000010000000100010011;
ROM[1696] <= 32'b00000100000001101010001110000011;
ROM[1697] <= 32'b00000000011100010010000000100011;
ROM[1698] <= 32'b00000000010000010000000100010011;
ROM[1699] <= 32'b11111111110000010000000100010011;
ROM[1700] <= 32'b00000000000000010010001110000011;
ROM[1701] <= 32'b11111111110000010000000100010011;
ROM[1702] <= 32'b00000000000000010010010000000011;
ROM[1703] <= 32'b00000000011101000000001110110011;
ROM[1704] <= 32'b00000000011100010010000000100011;
ROM[1705] <= 32'b00000000010000010000000100010011;
ROM[1706] <= 32'b00000110100000000000001110010011;
ROM[1707] <= 32'b00000000011100010010000000100011;
ROM[1708] <= 32'b00000000010000010000000100010011;
ROM[1709] <= 32'b00000100000001101010001110000011;
ROM[1710] <= 32'b00000000011100010010000000100011;
ROM[1711] <= 32'b00000000010000010000000100010011;
ROM[1712] <= 32'b11111111110000010000000100010011;
ROM[1713] <= 32'b00000000000000010010001110000011;
ROM[1714] <= 32'b11111111110000010000000100010011;
ROM[1715] <= 32'b00000000000000010010010000000011;
ROM[1716] <= 32'b00000000011101000000001110110011;
ROM[1717] <= 32'b00000000011100010010000000100011;
ROM[1718] <= 32'b00000000010000010000000100010011;
ROM[1719] <= 32'b11111111110000010000000100010011;
ROM[1720] <= 32'b00000000000000010010001110000011;
ROM[1721] <= 32'b00000000000000111000001100010011;
ROM[1722] <= 32'b00000000110100110000010000110011;
ROM[1723] <= 32'b00000000000001000010001110000011;
ROM[1724] <= 32'b00000000011100010010000000100011;
ROM[1725] <= 32'b00000000010000010000000100010011;
ROM[1726] <= 32'b00000110100000000000001110010011;
ROM[1727] <= 32'b00000000011100010010000000100011;
ROM[1728] <= 32'b00000000010000010000000100010011;
ROM[1729] <= 32'b00000100000001101010001110000011;
ROM[1730] <= 32'b00000000011100010010000000100011;
ROM[1731] <= 32'b00000000010000010000000100010011;
ROM[1732] <= 32'b11111111110000010000000100010011;
ROM[1733] <= 32'b00000000000000010010001110000011;
ROM[1734] <= 32'b11111111110000010000000100010011;
ROM[1735] <= 32'b00000000000000010010010000000011;
ROM[1736] <= 32'b00000000011101000000001110110011;
ROM[1737] <= 32'b00000000011100010010000000100011;
ROM[1738] <= 32'b00000000010000010000000100010011;
ROM[1739] <= 32'b11111111110000010000000100010011;
ROM[1740] <= 32'b00000000000000010010001110000011;
ROM[1741] <= 32'b00000000000000111000001100010011;
ROM[1742] <= 32'b00000000110100110000010000110011;
ROM[1743] <= 32'b00000000000001000010001110000011;
ROM[1744] <= 32'b00000000011100010010000000100011;
ROM[1745] <= 32'b00000000010000010000000100010011;
ROM[1746] <= 32'b11111111110000010000000100010011;
ROM[1747] <= 32'b00000000000000010010001110000011;
ROM[1748] <= 32'b11111111110000010000000100010011;
ROM[1749] <= 32'b00000000000000010010010000000011;
ROM[1750] <= 32'b00000000011101000000001110110011;
ROM[1751] <= 32'b00000000011100010010000000100011;
ROM[1752] <= 32'b00000000010000010000000100010011;
ROM[1753] <= 32'b11111111110000010000000100010011;
ROM[1754] <= 32'b00000000000000010010001110000011;
ROM[1755] <= 32'b00000000011101100010000000100011;
ROM[1756] <= 32'b11111111110000010000000100010011;
ROM[1757] <= 32'b00000000000000010010001110000011;
ROM[1758] <= 32'b00000000000000111000001100010011;
ROM[1759] <= 32'b00000000000001100010001110000011;
ROM[1760] <= 32'b00000000011100010010000000100011;
ROM[1761] <= 32'b00000000010000010000000100010011;
ROM[1762] <= 32'b11111111110000010000000100010011;
ROM[1763] <= 32'b00000000000000010010001110000011;
ROM[1764] <= 32'b00000000110100110000010000110011;
ROM[1765] <= 32'b00000000011101000010000000100011;
ROM[1766] <= 32'b00000111000000000000001110010011;
ROM[1767] <= 32'b00000000011100010010000000100011;
ROM[1768] <= 32'b00000000010000010000000100010011;
ROM[1769] <= 32'b00000100000001101010001110000011;
ROM[1770] <= 32'b00000000011100010010000000100011;
ROM[1771] <= 32'b00000000010000010000000100010011;
ROM[1772] <= 32'b11111111110000010000000100010011;
ROM[1773] <= 32'b00000000000000010010001110000011;
ROM[1774] <= 32'b11111111110000010000000100010011;
ROM[1775] <= 32'b00000000000000010010010000000011;
ROM[1776] <= 32'b00000000011101000000001110110011;
ROM[1777] <= 32'b00000000011100010010000000100011;
ROM[1778] <= 32'b00000000010000010000000100010011;
ROM[1779] <= 32'b00000110110000000000001110010011;
ROM[1780] <= 32'b00000000011100010010000000100011;
ROM[1781] <= 32'b00000000010000010000000100010011;
ROM[1782] <= 32'b00000100000001101010001110000011;
ROM[1783] <= 32'b00000000011100010010000000100011;
ROM[1784] <= 32'b00000000010000010000000100010011;
ROM[1785] <= 32'b11111111110000010000000100010011;
ROM[1786] <= 32'b00000000000000010010001110000011;
ROM[1787] <= 32'b11111111110000010000000100010011;
ROM[1788] <= 32'b00000000000000010010010000000011;
ROM[1789] <= 32'b00000000011101000000001110110011;
ROM[1790] <= 32'b00000000011100010010000000100011;
ROM[1791] <= 32'b00000000010000010000000100010011;
ROM[1792] <= 32'b11111111110000010000000100010011;
ROM[1793] <= 32'b00000000000000010010001110000011;
ROM[1794] <= 32'b00000000000000111000001100010011;
ROM[1795] <= 32'b00000000110100110000010000110011;
ROM[1796] <= 32'b00000000000001000010001110000011;
ROM[1797] <= 32'b00000000011100010010000000100011;
ROM[1798] <= 32'b00000000010000010000000100010011;
ROM[1799] <= 32'b00000110110000000000001110010011;
ROM[1800] <= 32'b00000000011100010010000000100011;
ROM[1801] <= 32'b00000000010000010000000100010011;
ROM[1802] <= 32'b00000100000001101010001110000011;
ROM[1803] <= 32'b00000000011100010010000000100011;
ROM[1804] <= 32'b00000000010000010000000100010011;
ROM[1805] <= 32'b11111111110000010000000100010011;
ROM[1806] <= 32'b00000000000000010010001110000011;
ROM[1807] <= 32'b11111111110000010000000100010011;
ROM[1808] <= 32'b00000000000000010010010000000011;
ROM[1809] <= 32'b00000000011101000000001110110011;
ROM[1810] <= 32'b00000000011100010010000000100011;
ROM[1811] <= 32'b00000000010000010000000100010011;
ROM[1812] <= 32'b11111111110000010000000100010011;
ROM[1813] <= 32'b00000000000000010010001110000011;
ROM[1814] <= 32'b00000000000000111000001100010011;
ROM[1815] <= 32'b00000000110100110000010000110011;
ROM[1816] <= 32'b00000000000001000010001110000011;
ROM[1817] <= 32'b00000000011100010010000000100011;
ROM[1818] <= 32'b00000000010000010000000100010011;
ROM[1819] <= 32'b11111111110000010000000100010011;
ROM[1820] <= 32'b00000000000000010010001110000011;
ROM[1821] <= 32'b11111111110000010000000100010011;
ROM[1822] <= 32'b00000000000000010010010000000011;
ROM[1823] <= 32'b00000000011101000000001110110011;
ROM[1824] <= 32'b00000000011100010010000000100011;
ROM[1825] <= 32'b00000000010000010000000100010011;
ROM[1826] <= 32'b11111111110000010000000100010011;
ROM[1827] <= 32'b00000000000000010010001110000011;
ROM[1828] <= 32'b00000000011101100010000000100011;
ROM[1829] <= 32'b11111111110000010000000100010011;
ROM[1830] <= 32'b00000000000000010010001110000011;
ROM[1831] <= 32'b00000000000000111000001100010011;
ROM[1832] <= 32'b00000000000001100010001110000011;
ROM[1833] <= 32'b00000000011100010010000000100011;
ROM[1834] <= 32'b00000000010000010000000100010011;
ROM[1835] <= 32'b11111111110000010000000100010011;
ROM[1836] <= 32'b00000000000000010010001110000011;
ROM[1837] <= 32'b00000000110100110000010000110011;
ROM[1838] <= 32'b00000000011101000010000000100011;
ROM[1839] <= 32'b00000111010000000000001110010011;
ROM[1840] <= 32'b00000000011100010010000000100011;
ROM[1841] <= 32'b00000000010000010000000100010011;
ROM[1842] <= 32'b00000100000001101010001110000011;
ROM[1843] <= 32'b00000000011100010010000000100011;
ROM[1844] <= 32'b00000000010000010000000100010011;
ROM[1845] <= 32'b11111111110000010000000100010011;
ROM[1846] <= 32'b00000000000000010010001110000011;
ROM[1847] <= 32'b11111111110000010000000100010011;
ROM[1848] <= 32'b00000000000000010010010000000011;
ROM[1849] <= 32'b00000000011101000000001110110011;
ROM[1850] <= 32'b00000000011100010010000000100011;
ROM[1851] <= 32'b00000000010000010000000100010011;
ROM[1852] <= 32'b00000111000000000000001110010011;
ROM[1853] <= 32'b00000000011100010010000000100011;
ROM[1854] <= 32'b00000000010000010000000100010011;
ROM[1855] <= 32'b00000100000001101010001110000011;
ROM[1856] <= 32'b00000000011100010010000000100011;
ROM[1857] <= 32'b00000000010000010000000100010011;
ROM[1858] <= 32'b11111111110000010000000100010011;
ROM[1859] <= 32'b00000000000000010010001110000011;
ROM[1860] <= 32'b11111111110000010000000100010011;
ROM[1861] <= 32'b00000000000000010010010000000011;
ROM[1862] <= 32'b00000000011101000000001110110011;
ROM[1863] <= 32'b00000000011100010010000000100011;
ROM[1864] <= 32'b00000000010000010000000100010011;
ROM[1865] <= 32'b11111111110000010000000100010011;
ROM[1866] <= 32'b00000000000000010010001110000011;
ROM[1867] <= 32'b00000000000000111000001100010011;
ROM[1868] <= 32'b00000000110100110000010000110011;
ROM[1869] <= 32'b00000000000001000010001110000011;
ROM[1870] <= 32'b00000000011100010010000000100011;
ROM[1871] <= 32'b00000000010000010000000100010011;
ROM[1872] <= 32'b00000111000000000000001110010011;
ROM[1873] <= 32'b00000000011100010010000000100011;
ROM[1874] <= 32'b00000000010000010000000100010011;
ROM[1875] <= 32'b00000100000001101010001110000011;
ROM[1876] <= 32'b00000000011100010010000000100011;
ROM[1877] <= 32'b00000000010000010000000100010011;
ROM[1878] <= 32'b11111111110000010000000100010011;
ROM[1879] <= 32'b00000000000000010010001110000011;
ROM[1880] <= 32'b11111111110000010000000100010011;
ROM[1881] <= 32'b00000000000000010010010000000011;
ROM[1882] <= 32'b00000000011101000000001110110011;
ROM[1883] <= 32'b00000000011100010010000000100011;
ROM[1884] <= 32'b00000000010000010000000100010011;
ROM[1885] <= 32'b11111111110000010000000100010011;
ROM[1886] <= 32'b00000000000000010010001110000011;
ROM[1887] <= 32'b00000000000000111000001100010011;
ROM[1888] <= 32'b00000000110100110000010000110011;
ROM[1889] <= 32'b00000000000001000010001110000011;
ROM[1890] <= 32'b00000000011100010010000000100011;
ROM[1891] <= 32'b00000000010000010000000100010011;
ROM[1892] <= 32'b11111111110000010000000100010011;
ROM[1893] <= 32'b00000000000000010010001110000011;
ROM[1894] <= 32'b11111111110000010000000100010011;
ROM[1895] <= 32'b00000000000000010010010000000011;
ROM[1896] <= 32'b00000000011101000000001110110011;
ROM[1897] <= 32'b00000000011100010010000000100011;
ROM[1898] <= 32'b00000000010000010000000100010011;
ROM[1899] <= 32'b11111111110000010000000100010011;
ROM[1900] <= 32'b00000000000000010010001110000011;
ROM[1901] <= 32'b00000000011101100010000000100011;
ROM[1902] <= 32'b11111111110000010000000100010011;
ROM[1903] <= 32'b00000000000000010010001110000011;
ROM[1904] <= 32'b00000000000000111000001100010011;
ROM[1905] <= 32'b00000000000001100010001110000011;
ROM[1906] <= 32'b00000000011100010010000000100011;
ROM[1907] <= 32'b00000000010000010000000100010011;
ROM[1908] <= 32'b11111111110000010000000100010011;
ROM[1909] <= 32'b00000000000000010010001110000011;
ROM[1910] <= 32'b00000000110100110000010000110011;
ROM[1911] <= 32'b00000000011101000010000000100011;
ROM[1912] <= 32'b00000111100000000000001110010011;
ROM[1913] <= 32'b00000000011100010010000000100011;
ROM[1914] <= 32'b00000000010000010000000100010011;
ROM[1915] <= 32'b00000100000001101010001110000011;
ROM[1916] <= 32'b00000000011100010010000000100011;
ROM[1917] <= 32'b00000000010000010000000100010011;
ROM[1918] <= 32'b11111111110000010000000100010011;
ROM[1919] <= 32'b00000000000000010010001110000011;
ROM[1920] <= 32'b11111111110000010000000100010011;
ROM[1921] <= 32'b00000000000000010010010000000011;
ROM[1922] <= 32'b00000000011101000000001110110011;
ROM[1923] <= 32'b00000000011100010010000000100011;
ROM[1924] <= 32'b00000000010000010000000100010011;
ROM[1925] <= 32'b00000111010000000000001110010011;
ROM[1926] <= 32'b00000000011100010010000000100011;
ROM[1927] <= 32'b00000000010000010000000100010011;
ROM[1928] <= 32'b00000100000001101010001110000011;
ROM[1929] <= 32'b00000000011100010010000000100011;
ROM[1930] <= 32'b00000000010000010000000100010011;
ROM[1931] <= 32'b11111111110000010000000100010011;
ROM[1932] <= 32'b00000000000000010010001110000011;
ROM[1933] <= 32'b11111111110000010000000100010011;
ROM[1934] <= 32'b00000000000000010010010000000011;
ROM[1935] <= 32'b00000000011101000000001110110011;
ROM[1936] <= 32'b00000000011100010010000000100011;
ROM[1937] <= 32'b00000000010000010000000100010011;
ROM[1938] <= 32'b11111111110000010000000100010011;
ROM[1939] <= 32'b00000000000000010010001110000011;
ROM[1940] <= 32'b00000000000000111000001100010011;
ROM[1941] <= 32'b00000000110100110000010000110011;
ROM[1942] <= 32'b00000000000001000010001110000011;
ROM[1943] <= 32'b00000000011100010010000000100011;
ROM[1944] <= 32'b00000000010000010000000100010011;
ROM[1945] <= 32'b00000111010000000000001110010011;
ROM[1946] <= 32'b00000000011100010010000000100011;
ROM[1947] <= 32'b00000000010000010000000100010011;
ROM[1948] <= 32'b00000100000001101010001110000011;
ROM[1949] <= 32'b00000000011100010010000000100011;
ROM[1950] <= 32'b00000000010000010000000100010011;
ROM[1951] <= 32'b11111111110000010000000100010011;
ROM[1952] <= 32'b00000000000000010010001110000011;
ROM[1953] <= 32'b11111111110000010000000100010011;
ROM[1954] <= 32'b00000000000000010010010000000011;
ROM[1955] <= 32'b00000000011101000000001110110011;
ROM[1956] <= 32'b00000000011100010010000000100011;
ROM[1957] <= 32'b00000000010000010000000100010011;
ROM[1958] <= 32'b11111111110000010000000100010011;
ROM[1959] <= 32'b00000000000000010010001110000011;
ROM[1960] <= 32'b00000000000000111000001100010011;
ROM[1961] <= 32'b00000000110100110000010000110011;
ROM[1962] <= 32'b00000000000001000010001110000011;
ROM[1963] <= 32'b00000000011100010010000000100011;
ROM[1964] <= 32'b00000000010000010000000100010011;
ROM[1965] <= 32'b11111111110000010000000100010011;
ROM[1966] <= 32'b00000000000000010010001110000011;
ROM[1967] <= 32'b11111111110000010000000100010011;
ROM[1968] <= 32'b00000000000000010010010000000011;
ROM[1969] <= 32'b00000000011101000000001110110011;
ROM[1970] <= 32'b00000000011100010010000000100011;
ROM[1971] <= 32'b00000000010000010000000100010011;
ROM[1972] <= 32'b11111111110000010000000100010011;
ROM[1973] <= 32'b00000000000000010010001110000011;
ROM[1974] <= 32'b00000000011101100010000000100011;
ROM[1975] <= 32'b11111111110000010000000100010011;
ROM[1976] <= 32'b00000000000000010010001110000011;
ROM[1977] <= 32'b00000000000000111000001100010011;
ROM[1978] <= 32'b00000000000001100010001110000011;
ROM[1979] <= 32'b00000000011100010010000000100011;
ROM[1980] <= 32'b00000000010000010000000100010011;
ROM[1981] <= 32'b11111111110000010000000100010011;
ROM[1982] <= 32'b00000000000000010010001110000011;
ROM[1983] <= 32'b00000000110100110000010000110011;
ROM[1984] <= 32'b00000000011101000010000000100011;
ROM[1985] <= 32'b00000000000000000000001110010011;
ROM[1986] <= 32'b00000000011100010010000000100011;
ROM[1987] <= 32'b00000000010000010000000100010011;
ROM[1988] <= 32'b00000001010000000000001110010011;
ROM[1989] <= 32'b01000000011100011000001110110011;
ROM[1990] <= 32'b00000000000000111010000010000011;
ROM[1991] <= 32'b11111111110000010000000100010011;
ROM[1992] <= 32'b00000000000000010010001110000011;
ROM[1993] <= 32'b00000000011100100010000000100011;
ROM[1994] <= 32'b00000000010000100000000100010011;
ROM[1995] <= 32'b00000001010000000000001110010011;
ROM[1996] <= 32'b01000000011100011000001110110011;
ROM[1997] <= 32'b00000000010000111010000110000011;
ROM[1998] <= 32'b00000000100000111010001000000011;
ROM[1999] <= 32'b00000000110000111010001010000011;
ROM[2000] <= 32'b00000001000000111010001100000011;
ROM[2001] <= 32'b00000000000000001000000011100111;
ROM[2002] <= 32'b00000000000000010010000000100011;
ROM[2003] <= 32'b00000000010000010000000100010011;
ROM[2004] <= 32'b00000000000000010010000000100011;
ROM[2005] <= 32'b00000000010000010000000100010011;
ROM[2006] <= 32'b00000000000000010010000000100011;
ROM[2007] <= 32'b00000000010000010000000100010011;
ROM[2008] <= 32'b00000000000000000000001110010011;
ROM[2009] <= 32'b00000000011100010010000000100011;
ROM[2010] <= 32'b00000000010000010000000100010011;
ROM[2011] <= 32'b11111111110000010000000100010011;
ROM[2012] <= 32'b00000000000000010010001110000011;
ROM[2013] <= 32'b00000000011100011010000000100011;
ROM[2014] <= 32'b00000000000000100010001110000011;
ROM[2015] <= 32'b00000000011100010010000000100011;
ROM[2016] <= 32'b00000000010000010000000100010011;
ROM[2017] <= 32'b11111111110000010000000100010011;
ROM[2018] <= 32'b00000000000000010010001110000011;
ROM[2019] <= 32'b00000000011100011010001000100011;
ROM[2020] <= 32'b00000000000000000000001110010011;
ROM[2021] <= 32'b00000000011100010010000000100011;
ROM[2022] <= 32'b00000000010000010000000100010011;
ROM[2023] <= 32'b11111111110000010000000100010011;
ROM[2024] <= 32'b00000000000000010010001110000011;
ROM[2025] <= 32'b00000000011100011010010000100011;
ROM[2026] <= 32'b00000000100000011010001110000011;
ROM[2027] <= 32'b00000000011100010010000000100011;
ROM[2028] <= 32'b00000000010000010000000100010011;
ROM[2029] <= 32'b00000111110000000000001110010011;
ROM[2030] <= 32'b00000000011100010010000000100011;
ROM[2031] <= 32'b00000000010000010000000100010011;
ROM[2032] <= 32'b11111111110000010000000100010011;
ROM[2033] <= 32'b00000000000000010010001110000011;
ROM[2034] <= 32'b11111111110000010000000100010011;
ROM[2035] <= 32'b00000000000000010010010000000011;
ROM[2036] <= 32'b00000000011101000010001110110011;
ROM[2037] <= 32'b00000000011100010010000000100011;
ROM[2038] <= 32'b00000000010000010000000100010011;
ROM[2039] <= 32'b11111111110000010000000100010011;
ROM[2040] <= 32'b00000000000000010010001110000011;
ROM[2041] <= 32'b01000000011100000000001110110011;
ROM[2042] <= 32'b00000000000100111000001110010011;
ROM[2043] <= 32'b00000000011100010010000000100011;
ROM[2044] <= 32'b00000000010000010000000100010011;
ROM[2045] <= 32'b11111111110000010000000100010011;
ROM[2046] <= 32'b00000000000000010010001110000011;
ROM[2047] <= 32'b00000000000000111000101001100011;
ROM[2048] <= 32'b00000000000000001000001110110111;
ROM[2049] <= 32'b11001110010000111000001110010011;
ROM[2050] <= 32'b00000000111000111000001110110011;
ROM[2051] <= 32'b00000000000000111000000011100111;
ROM[2052] <= 32'b00000000010000100010001110000011;
ROM[2053] <= 32'b00000000011100010010000000100011;
ROM[2054] <= 32'b00000000010000010000000100010011;
ROM[2055] <= 32'b00000000100000011010001110000011;
ROM[2056] <= 32'b00000000011100010010000000100011;
ROM[2057] <= 32'b00000000010000010000000100010011;
ROM[2058] <= 32'b00000100000001101010001110000011;
ROM[2059] <= 32'b00000000011100010010000000100011;
ROM[2060] <= 32'b00000000010000010000000100010011;
ROM[2061] <= 32'b11111111110000010000000100010011;
ROM[2062] <= 32'b00000000000000010010001110000011;
ROM[2063] <= 32'b11111111110000010000000100010011;
ROM[2064] <= 32'b00000000000000010010010000000011;
ROM[2065] <= 32'b00000000011101000000001110110011;
ROM[2066] <= 32'b00000000011100010010000000100011;
ROM[2067] <= 32'b00000000010000010000000100010011;
ROM[2068] <= 32'b11111111110000010000000100010011;
ROM[2069] <= 32'b00000000000000010010001110000011;
ROM[2070] <= 32'b00000000000000111000001100010011;
ROM[2071] <= 32'b00000000110100110000010000110011;
ROM[2072] <= 32'b00000000000001000010001110000011;
ROM[2073] <= 32'b00000000011100010010000000100011;
ROM[2074] <= 32'b00000000010000010000000100010011;
ROM[2075] <= 32'b11111111110000010000000100010011;
ROM[2076] <= 32'b00000000000000010010001110000011;
ROM[2077] <= 32'b11111111110000010000000100010011;
ROM[2078] <= 32'b00000000000000010010010000000011;
ROM[2079] <= 32'b00000000011101000111001110110011;
ROM[2080] <= 32'b00000000011100010010000000100011;
ROM[2081] <= 32'b00000000010000010000000100010011;
ROM[2082] <= 32'b00000000000000000000001110010011;
ROM[2083] <= 32'b00000000011100010010000000100011;
ROM[2084] <= 32'b00000000010000010000000100010011;
ROM[2085] <= 32'b11111111110000010000000100010011;
ROM[2086] <= 32'b00000000000000010010001110000011;
ROM[2087] <= 32'b11111111110000010000000100010011;
ROM[2088] <= 32'b00000000000000010010010000000011;
ROM[2089] <= 32'b00000000011101000010010010110011;
ROM[2090] <= 32'b00000000100000111010010100110011;
ROM[2091] <= 32'b00000000101001001000001110110011;
ROM[2092] <= 32'b00000000000100111000001110010011;
ROM[2093] <= 32'b00000000000100111111001110010011;
ROM[2094] <= 32'b00000000011100010010000000100011;
ROM[2095] <= 32'b00000000010000010000000100010011;
ROM[2096] <= 32'b11111111110000010000000100010011;
ROM[2097] <= 32'b00000000000000010010001110000011;
ROM[2098] <= 32'b01000000011100000000001110110011;
ROM[2099] <= 32'b00000000000100111000001110010011;
ROM[2100] <= 32'b00000000011100010010000000100011;
ROM[2101] <= 32'b00000000010000010000000100010011;
ROM[2102] <= 32'b11111111110000010000000100010011;
ROM[2103] <= 32'b00000000000000010010001110000011;
ROM[2104] <= 32'b00000000000000111000101001100011;
ROM[2105] <= 32'b00000000000000000111001110110111;
ROM[2106] <= 32'b10001110100000111000001110010011;
ROM[2107] <= 32'b00000000111000111000001110110011;
ROM[2108] <= 32'b00000000000000111000000011100111;
ROM[2109] <= 32'b00000001000100000100000011101111;
ROM[2110] <= 32'b00000000000000011010001110000011;
ROM[2111] <= 32'b00000000011100010010000000100011;
ROM[2112] <= 32'b00000000010000010000000100010011;
ROM[2113] <= 32'b00000000010000011010001110000011;
ROM[2114] <= 32'b00000000011100010010000000100011;
ROM[2115] <= 32'b00000000010000010000000100010011;
ROM[2116] <= 32'b11111111110000010000000100010011;
ROM[2117] <= 32'b00000000000000010010001110000011;
ROM[2118] <= 32'b11111111110000010000000100010011;
ROM[2119] <= 32'b00000000000000010010010000000011;
ROM[2120] <= 32'b00000000011101000000001110110011;
ROM[2121] <= 32'b00000000011100010010000000100011;
ROM[2122] <= 32'b00000000010000010000000100010011;
ROM[2123] <= 32'b11111111110000010000000100010011;
ROM[2124] <= 32'b00000000000000010010001110000011;
ROM[2125] <= 32'b00000000011100011010000000100011;
ROM[2126] <= 32'b01111100110000000100000011101111;
ROM[2127] <= 32'b00000000010000011010001110000011;
ROM[2128] <= 32'b00000000011100010010000000100011;
ROM[2129] <= 32'b00000000010000010000000100010011;
ROM[2130] <= 32'b00000000010000011010001110000011;
ROM[2131] <= 32'b00000000011100010010000000100011;
ROM[2132] <= 32'b00000000010000010000000100010011;
ROM[2133] <= 32'b11111111110000010000000100010011;
ROM[2134] <= 32'b00000000000000010010001110000011;
ROM[2135] <= 32'b11111111110000010000000100010011;
ROM[2136] <= 32'b00000000000000010010010000000011;
ROM[2137] <= 32'b00000000011101000000001110110011;
ROM[2138] <= 32'b00000000011100010010000000100011;
ROM[2139] <= 32'b00000000010000010000000100010011;
ROM[2140] <= 32'b11111111110000010000000100010011;
ROM[2141] <= 32'b00000000000000010010001110000011;
ROM[2142] <= 32'b00000000011100011010001000100011;
ROM[2143] <= 32'b00000000100000011010001110000011;
ROM[2144] <= 32'b00000000011100010010000000100011;
ROM[2145] <= 32'b00000000010000010000000100010011;
ROM[2146] <= 32'b00000000010000000000001110010011;
ROM[2147] <= 32'b00000000011100010010000000100011;
ROM[2148] <= 32'b00000000010000010000000100010011;
ROM[2149] <= 32'b11111111110000010000000100010011;
ROM[2150] <= 32'b00000000000000010010001110000011;
ROM[2151] <= 32'b11111111110000010000000100010011;
ROM[2152] <= 32'b00000000000000010010010000000011;
ROM[2153] <= 32'b00000000011101000000001110110011;
ROM[2154] <= 32'b00000000011100010010000000100011;
ROM[2155] <= 32'b00000000010000010000000100010011;
ROM[2156] <= 32'b11111111110000010000000100010011;
ROM[2157] <= 32'b00000000000000010010001110000011;
ROM[2158] <= 32'b00000000011100011010010000100011;
ROM[2159] <= 32'b00101100110100000101000011101111;
ROM[2160] <= 32'b00000000000000011010001110000011;
ROM[2161] <= 32'b00000000011100010010000000100011;
ROM[2162] <= 32'b00000000010000010000000100010011;
ROM[2163] <= 32'b00000001010000000000001110010011;
ROM[2164] <= 32'b01000000011100011000001110110011;
ROM[2165] <= 32'b00000000000000111010000010000011;
ROM[2166] <= 32'b11111111110000010000000100010011;
ROM[2167] <= 32'b00000000000000010010001110000011;
ROM[2168] <= 32'b00000000011100100010000000100011;
ROM[2169] <= 32'b00000000010000100000000100010011;
ROM[2170] <= 32'b00000001010000000000001110010011;
ROM[2171] <= 32'b01000000011100011000001110110011;
ROM[2172] <= 32'b00000000010000111010000110000011;
ROM[2173] <= 32'b00000000100000111010001000000011;
ROM[2174] <= 32'b00000000110000111010001010000011;
ROM[2175] <= 32'b00000001000000111010001100000011;
ROM[2176] <= 32'b00000000000000001000000011100111;
ROM[2177] <= 32'b00000000000000100010001110000011;
ROM[2178] <= 32'b00000000011100010010000000100011;
ROM[2179] <= 32'b00000000010000010000000100010011;
ROM[2180] <= 32'b00000000000000000000001110010011;
ROM[2181] <= 32'b00000000011100010010000000100011;
ROM[2182] <= 32'b00000000010000010000000100010011;
ROM[2183] <= 32'b11111111110000010000000100010011;
ROM[2184] <= 32'b00000000000000010010001110000011;
ROM[2185] <= 32'b11111111110000010000000100010011;
ROM[2186] <= 32'b00000000000000010010010000000011;
ROM[2187] <= 32'b00000000011101000010001110110011;
ROM[2188] <= 32'b00000000011100010010000000100011;
ROM[2189] <= 32'b00000000010000010000000100010011;
ROM[2190] <= 32'b11111111110000010000000100010011;
ROM[2191] <= 32'b00000000000000010010001110000011;
ROM[2192] <= 32'b00000000000000111000101001100011;
ROM[2193] <= 32'b00000000000000000111001110110111;
ROM[2194] <= 32'b11000011000000111000001110010011;
ROM[2195] <= 32'b00000000111000111000001110110011;
ROM[2196] <= 32'b00000000000000111000000011100111;
ROM[2197] <= 32'b00101010010100000100000011101111;
ROM[2198] <= 32'b00000000000000100010001110000011;
ROM[2199] <= 32'b00000000011100010010000000100011;
ROM[2200] <= 32'b00000000010000010000000100010011;
ROM[2201] <= 32'b11111111110000010000000100010011;
ROM[2202] <= 32'b00000000000000010010001110000011;
ROM[2203] <= 32'b01000000011100000000001110110011;
ROM[2204] <= 32'b00000000011100010010000000100011;
ROM[2205] <= 32'b00000000010000010000000100010011;
ROM[2206] <= 32'b11111111110000010000000100010011;
ROM[2207] <= 32'b00000000000000010010001110000011;
ROM[2208] <= 32'b00000000011100100010000000100011;
ROM[2209] <= 32'b00100111010100000100000011101111;
ROM[2210] <= 32'b00000000000000100010001110000011;
ROM[2211] <= 32'b00000000011100010010000000100011;
ROM[2212] <= 32'b00000000010000010000000100010011;
ROM[2213] <= 32'b00000001010000000000001110010011;
ROM[2214] <= 32'b01000000011100011000001110110011;
ROM[2215] <= 32'b00000000000000111010000010000011;
ROM[2216] <= 32'b11111111110000010000000100010011;
ROM[2217] <= 32'b00000000000000010010001110000011;
ROM[2218] <= 32'b00000000011100100010000000100011;
ROM[2219] <= 32'b00000000010000100000000100010011;
ROM[2220] <= 32'b00000001010000000000001110010011;
ROM[2221] <= 32'b01000000011100011000001110110011;
ROM[2222] <= 32'b00000000010000111010000110000011;
ROM[2223] <= 32'b00000000100000111010001000000011;
ROM[2224] <= 32'b00000000110000111010001010000011;
ROM[2225] <= 32'b00000001000000111010001100000011;
ROM[2226] <= 32'b00000000000000001000000011100111;
ROM[2227] <= 32'b00000000000000010010000000100011;
ROM[2228] <= 32'b00000000010000010000000100010011;
ROM[2229] <= 32'b00000000000000010010000000100011;
ROM[2230] <= 32'b00000000010000010000000100010011;
ROM[2231] <= 32'b00000000000000010010000000100011;
ROM[2232] <= 32'b00000000010000010000000100010011;
ROM[2233] <= 32'b00000000010000100010001110000011;
ROM[2234] <= 32'b00000000011100010010000000100011;
ROM[2235] <= 32'b00000000010000010000000100010011;
ROM[2236] <= 32'b00000000000000000000001110010011;
ROM[2237] <= 32'b00000000011100010010000000100011;
ROM[2238] <= 32'b00000000010000010000000100010011;
ROM[2239] <= 32'b11111111110000010000000100010011;
ROM[2240] <= 32'b00000000000000010010001110000011;
ROM[2241] <= 32'b11111111110000010000000100010011;
ROM[2242] <= 32'b00000000000000010010010000000011;
ROM[2243] <= 32'b00000000011101000010010010110011;
ROM[2244] <= 32'b00000000100000111010010100110011;
ROM[2245] <= 32'b00000000101001001000001110110011;
ROM[2246] <= 32'b00000000000100111000001110010011;
ROM[2247] <= 32'b00000000000100111111001110010011;
ROM[2248] <= 32'b00000000011100010010000000100011;
ROM[2249] <= 32'b00000000010000010000000100010011;
ROM[2250] <= 32'b11111111110000010000000100010011;
ROM[2251] <= 32'b00000000000000010010001110000011;
ROM[2252] <= 32'b00000000000000111000101001100011;
ROM[2253] <= 32'b00000000000000000111001110110111;
ROM[2254] <= 32'b11011011000000111000001110010011;
ROM[2255] <= 32'b00000000111000111000001110110011;
ROM[2256] <= 32'b00000000000000111000000011100111;
ROM[2257] <= 32'b00101011100100000100000011101111;
ROM[2258] <= 32'b00000000000100000000001110010011;
ROM[2259] <= 32'b00000000011100010010000000100011;
ROM[2260] <= 32'b00000000010000010000000100010011;
ROM[2261] <= 32'b11111111110000010000000100010011;
ROM[2262] <= 32'b00000000000000010010001110000011;
ROM[2263] <= 32'b01000000011100000000001110110011;
ROM[2264] <= 32'b00000000011100010010000000100011;
ROM[2265] <= 32'b00000000010000010000000100010011;
ROM[2266] <= 32'b00000001010000000000001110010011;
ROM[2267] <= 32'b01000000011100011000001110110011;
ROM[2268] <= 32'b00000000000000111010000010000011;
ROM[2269] <= 32'b11111111110000010000000100010011;
ROM[2270] <= 32'b00000000000000010010001110000011;
ROM[2271] <= 32'b00000000011100100010000000100011;
ROM[2272] <= 32'b00000000010000100000000100010011;
ROM[2273] <= 32'b00000001010000000000001110010011;
ROM[2274] <= 32'b01000000011100011000001110110011;
ROM[2275] <= 32'b00000000010000111010000110000011;
ROM[2276] <= 32'b00000000100000111010001000000011;
ROM[2277] <= 32'b00000000110000111010001010000011;
ROM[2278] <= 32'b00000001000000111010001100000011;
ROM[2279] <= 32'b00000000000000001000000011100111;
ROM[2280] <= 32'b00100101110100000100000011101111;
ROM[2281] <= 32'b00000000000000100010001110000011;
ROM[2282] <= 32'b00000000011100010010000000100011;
ROM[2283] <= 32'b00000000010000010000000100010011;
ROM[2284] <= 32'b00000000000000000000001110010011;
ROM[2285] <= 32'b00000000011100010010000000100011;
ROM[2286] <= 32'b00000000010000010000000100010011;
ROM[2287] <= 32'b11111111110000010000000100010011;
ROM[2288] <= 32'b00000000000000010010001110000011;
ROM[2289] <= 32'b11111111110000010000000100010011;
ROM[2290] <= 32'b00000000000000010010010000000011;
ROM[2291] <= 32'b00000000011101000010001110110011;
ROM[2292] <= 32'b00000000011100010010000000100011;
ROM[2293] <= 32'b00000000010000010000000100010011;
ROM[2294] <= 32'b00000000010000100010001110000011;
ROM[2295] <= 32'b00000000011100010010000000100011;
ROM[2296] <= 32'b00000000010000010000000100010011;
ROM[2297] <= 32'b00000000000000000000001110010011;
ROM[2298] <= 32'b00000000011100010010000000100011;
ROM[2299] <= 32'b00000000010000010000000100010011;
ROM[2300] <= 32'b11111111110000010000000100010011;
ROM[2301] <= 32'b00000000000000010010001110000011;
ROM[2302] <= 32'b11111111110000010000000100010011;
ROM[2303] <= 32'b00000000000000010010010000000011;
ROM[2304] <= 32'b00000000011101000010001110110011;
ROM[2305] <= 32'b00000000011100010010000000100011;
ROM[2306] <= 32'b00000000010000010000000100010011;
ROM[2307] <= 32'b11111111110000010000000100010011;
ROM[2308] <= 32'b00000000000000010010001110000011;
ROM[2309] <= 32'b11111111110000010000000100010011;
ROM[2310] <= 32'b00000000000000010010010000000011;
ROM[2311] <= 32'b00000000011101000010010010110011;
ROM[2312] <= 32'b00000000100000111010010100110011;
ROM[2313] <= 32'b00000000101001001000001110110011;
ROM[2314] <= 32'b00000000000100111000001110010011;
ROM[2315] <= 32'b00000000000100111111001110010011;
ROM[2316] <= 32'b00000000011100010010000000100011;
ROM[2317] <= 32'b00000000010000010000000100010011;
ROM[2318] <= 32'b11111111110000010000000100010011;
ROM[2319] <= 32'b00000000000000010010001110000011;
ROM[2320] <= 32'b01000000011100000000001110110011;
ROM[2321] <= 32'b00000000000100111000001110010011;
ROM[2322] <= 32'b00000000011100010010000000100011;
ROM[2323] <= 32'b00000000010000010000000100010011;
ROM[2324] <= 32'b11111111110000010000000100010011;
ROM[2325] <= 32'b00000000000000010010001110000011;
ROM[2326] <= 32'b00000000011100011010001000100011;
ROM[2327] <= 32'b00000000000000100010001110000011;
ROM[2328] <= 32'b00000000011100010010000000100011;
ROM[2329] <= 32'b00000000010000010000000100010011;
ROM[2330] <= 32'b00000000000000000010001110110111;
ROM[2331] <= 32'b01001011010000111000001110010011;
ROM[2332] <= 32'b00000000111000111000001110110011;
ROM[2333] <= 32'b00000000011100010010000000100011;
ROM[2334] <= 32'b00000000010000010000000100010011;
ROM[2335] <= 32'b00000000001100010010000000100011;
ROM[2336] <= 32'b00000000010000010000000100010011;
ROM[2337] <= 32'b00000000010000010010000000100011;
ROM[2338] <= 32'b00000000010000010000000100010011;
ROM[2339] <= 32'b00000000010100010010000000100011;
ROM[2340] <= 32'b00000000010000010000000100010011;
ROM[2341] <= 32'b00000000011000010010000000100011;
ROM[2342] <= 32'b00000000010000010000000100010011;
ROM[2343] <= 32'b00000001010000000000001110010011;
ROM[2344] <= 32'b00000000010000111000001110010011;
ROM[2345] <= 32'b01000000011100010000001110110011;
ROM[2346] <= 32'b00000000011100000000001000110011;
ROM[2347] <= 32'b00000000001000000000000110110011;
ROM[2348] <= 32'b11010101010111111111000011101111;
ROM[2349] <= 32'b11111111110000010000000100010011;
ROM[2350] <= 32'b00000000000000010010001110000011;
ROM[2351] <= 32'b00000000011100100010000000100011;
ROM[2352] <= 32'b00000000010000100010001110000011;
ROM[2353] <= 32'b00000000011100010010000000100011;
ROM[2354] <= 32'b00000000010000010000000100010011;
ROM[2355] <= 32'b00000000000000000010001110110111;
ROM[2356] <= 32'b01010001100000111000001110010011;
ROM[2357] <= 32'b00000000111000111000001110110011;
ROM[2358] <= 32'b00000000011100010010000000100011;
ROM[2359] <= 32'b00000000010000010000000100010011;
ROM[2360] <= 32'b00000000001100010010000000100011;
ROM[2361] <= 32'b00000000010000010000000100010011;
ROM[2362] <= 32'b00000000010000010010000000100011;
ROM[2363] <= 32'b00000000010000010000000100010011;
ROM[2364] <= 32'b00000000010100010010000000100011;
ROM[2365] <= 32'b00000000010000010000000100010011;
ROM[2366] <= 32'b00000000011000010010000000100011;
ROM[2367] <= 32'b00000000010000010000000100010011;
ROM[2368] <= 32'b00000001010000000000001110010011;
ROM[2369] <= 32'b00000000010000111000001110010011;
ROM[2370] <= 32'b01000000011100010000001110110011;
ROM[2371] <= 32'b00000000011100000000001000110011;
ROM[2372] <= 32'b00000000001000000000000110110011;
ROM[2373] <= 32'b11001111000111111111000011101111;
ROM[2374] <= 32'b11111111110000010000000100010011;
ROM[2375] <= 32'b00000000000000010010001110000011;
ROM[2376] <= 32'b00000000011100100010001000100011;
ROM[2377] <= 32'b00000000000000000000001110010011;
ROM[2378] <= 32'b00000000011100010010000000100011;
ROM[2379] <= 32'b00000000010000010000000100010011;
ROM[2380] <= 32'b11111111110000010000000100010011;
ROM[2381] <= 32'b00000000000000010010001110000011;
ROM[2382] <= 32'b00000000011100011010000000100011;
ROM[2383] <= 32'b00000000010000100010001110000011;
ROM[2384] <= 32'b00000000011100010010000000100011;
ROM[2385] <= 32'b00000000010000010000000100010011;
ROM[2386] <= 32'b00000000000000100010001110000011;
ROM[2387] <= 32'b00000000011100010010000000100011;
ROM[2388] <= 32'b00000000010000010000000100010011;
ROM[2389] <= 32'b11111111110000010000000100010011;
ROM[2390] <= 32'b00000000000000010010001110000011;
ROM[2391] <= 32'b11111111110000010000000100010011;
ROM[2392] <= 32'b00000000000000010010010000000011;
ROM[2393] <= 32'b00000000100000111010001110110011;
ROM[2394] <= 32'b00000000011100010010000000100011;
ROM[2395] <= 32'b00000000010000010000000100010011;
ROM[2396] <= 32'b11111111110000010000000100010011;
ROM[2397] <= 32'b00000000000000010010001110000011;
ROM[2398] <= 32'b01000000011100000000001110110011;
ROM[2399] <= 32'b00000000000100111000001110010011;
ROM[2400] <= 32'b00000000011100010010000000100011;
ROM[2401] <= 32'b00000000010000010000000100010011;
ROM[2402] <= 32'b11111111110000010000000100010011;
ROM[2403] <= 32'b00000000000000010010001110000011;
ROM[2404] <= 32'b00000000011100011010010000100011;
ROM[2405] <= 32'b00000000100000011010001110000011;
ROM[2406] <= 32'b00000000011100010010000000100011;
ROM[2407] <= 32'b00000000010000010000000100010011;
ROM[2408] <= 32'b11111111110000010000000100010011;
ROM[2409] <= 32'b00000000000000010010001110000011;
ROM[2410] <= 32'b01000000011100000000001110110011;
ROM[2411] <= 32'b00000000000100111000001110010011;
ROM[2412] <= 32'b00000000011100010010000000100011;
ROM[2413] <= 32'b00000000010000010000000100010011;
ROM[2414] <= 32'b11111111110000010000000100010011;
ROM[2415] <= 32'b00000000000000010010001110000011;
ROM[2416] <= 32'b00000000000000111000101001100011;
ROM[2417] <= 32'b00000000000000001000001110110111;
ROM[2418] <= 32'b11101100000000111000001110010011;
ROM[2419] <= 32'b00000000111000111000001110110011;
ROM[2420] <= 32'b00000000000000111000000011100111;
ROM[2421] <= 32'b00000000000000100010001110000011;
ROM[2422] <= 32'b00000000011100010010000000100011;
ROM[2423] <= 32'b00000000010000010000000100010011;
ROM[2424] <= 32'b00000000010000100010001110000011;
ROM[2425] <= 32'b00000000011100010010000000100011;
ROM[2426] <= 32'b00000000010000010000000100010011;
ROM[2427] <= 32'b11111111110000010000000100010011;
ROM[2428] <= 32'b00000000000000010010001110000011;
ROM[2429] <= 32'b11111111110000010000000100010011;
ROM[2430] <= 32'b00000000000000010010010000000011;
ROM[2431] <= 32'b01000000011101000000001110110011;
ROM[2432] <= 32'b00000000011100010010000000100011;
ROM[2433] <= 32'b00000000010000010000000100010011;
ROM[2434] <= 32'b11111111110000010000000100010011;
ROM[2435] <= 32'b00000000000000010010001110000011;
ROM[2436] <= 32'b00000000011100100010000000100011;
ROM[2437] <= 32'b00000000000000011010001110000011;
ROM[2438] <= 32'b00000000011100010010000000100011;
ROM[2439] <= 32'b00000000010000010000000100010011;
ROM[2440] <= 32'b00000000000100000000001110010011;
ROM[2441] <= 32'b00000000011100010010000000100011;
ROM[2442] <= 32'b00000000010000010000000100010011;
ROM[2443] <= 32'b11111111110000010000000100010011;
ROM[2444] <= 32'b00000000000000010010001110000011;
ROM[2445] <= 32'b11111111110000010000000100010011;
ROM[2446] <= 32'b00000000000000010010010000000011;
ROM[2447] <= 32'b00000000011101000000001110110011;
ROM[2448] <= 32'b00000000011100010010000000100011;
ROM[2449] <= 32'b00000000010000010000000100010011;
ROM[2450] <= 32'b11111111110000010000000100010011;
ROM[2451] <= 32'b00000000000000010010001110000011;
ROM[2452] <= 32'b00000000011100011010000000100011;
ROM[2453] <= 32'b00000000010000100010001110000011;
ROM[2454] <= 32'b00000000011100010010000000100011;
ROM[2455] <= 32'b00000000010000010000000100010011;
ROM[2456] <= 32'b00000000000000100010001110000011;
ROM[2457] <= 32'b00000000011100010010000000100011;
ROM[2458] <= 32'b00000000010000010000000100010011;
ROM[2459] <= 32'b11111111110000010000000100010011;
ROM[2460] <= 32'b00000000000000010010001110000011;
ROM[2461] <= 32'b11111111110000010000000100010011;
ROM[2462] <= 32'b00000000000000010010010000000011;
ROM[2463] <= 32'b00000000100000111010001110110011;
ROM[2464] <= 32'b00000000011100010010000000100011;
ROM[2465] <= 32'b00000000010000010000000100010011;
ROM[2466] <= 32'b11111111110000010000000100010011;
ROM[2467] <= 32'b00000000000000010010001110000011;
ROM[2468] <= 32'b01000000011100000000001110110011;
ROM[2469] <= 32'b00000000000100111000001110010011;
ROM[2470] <= 32'b00000000011100010010000000100011;
ROM[2471] <= 32'b00000000010000010000000100010011;
ROM[2472] <= 32'b11111111110000010000000100010011;
ROM[2473] <= 32'b00000000000000010010001110000011;
ROM[2474] <= 32'b00000000011100011010010000100011;
ROM[2475] <= 32'b01101010010000000101000011101111;
ROM[2476] <= 32'b00000000010000011010001110000011;
ROM[2477] <= 32'b00000000011100010010000000100011;
ROM[2478] <= 32'b00000000010000010000000100010011;
ROM[2479] <= 32'b11111111110000010000000100010011;
ROM[2480] <= 32'b00000000000000010010001110000011;
ROM[2481] <= 32'b00000000000000111000101001100011;
ROM[2482] <= 32'b00000000000000000111001110110111;
ROM[2483] <= 32'b11111000100000111000001110010011;
ROM[2484] <= 32'b00000000111000111000001110110011;
ROM[2485] <= 32'b00000000000000111000000011100111;
ROM[2486] <= 32'b00001111110100000100000011101111;
ROM[2487] <= 32'b00000000000000011010001110000011;
ROM[2488] <= 32'b00000000011100010010000000100011;
ROM[2489] <= 32'b00000000010000010000000100010011;
ROM[2490] <= 32'b11111111110000010000000100010011;
ROM[2491] <= 32'b00000000000000010010001110000011;
ROM[2492] <= 32'b01000000011100000000001110110011;
ROM[2493] <= 32'b00000000011100010010000000100011;
ROM[2494] <= 32'b00000000010000010000000100010011;
ROM[2495] <= 32'b11111111110000010000000100010011;
ROM[2496] <= 32'b00000000000000010010001110000011;
ROM[2497] <= 32'b00000000011100011010000000100011;
ROM[2498] <= 32'b00001111110100000100000011101111;
ROM[2499] <= 32'b00000000000000011010001110000011;
ROM[2500] <= 32'b00000000011100010010000000100011;
ROM[2501] <= 32'b00000000010000010000000100010011;
ROM[2502] <= 32'b00000001010000000000001110010011;
ROM[2503] <= 32'b01000000011100011000001110110011;
ROM[2504] <= 32'b00000000000000111010000010000011;
ROM[2505] <= 32'b11111111110000010000000100010011;
ROM[2506] <= 32'b00000000000000010010001110000011;
ROM[2507] <= 32'b00000000011100100010000000100011;
ROM[2508] <= 32'b00000000010000100000000100010011;
ROM[2509] <= 32'b00000001010000000000001110010011;
ROM[2510] <= 32'b01000000011100011000001110110011;
ROM[2511] <= 32'b00000000010000111010000110000011;
ROM[2512] <= 32'b00000000100000111010001000000011;
ROM[2513] <= 32'b00000000110000111010001010000011;
ROM[2514] <= 32'b00000001000000111010001100000011;
ROM[2515] <= 32'b00000000000000001000000011100111;
ROM[2516] <= 32'b00000000000000100010001110000011;
ROM[2517] <= 32'b00000000011100010010000000100011;
ROM[2518] <= 32'b00000000010000010000000100010011;
ROM[2519] <= 32'b00000000010000100010001110000011;
ROM[2520] <= 32'b00000000011100010010000000100011;
ROM[2521] <= 32'b00000000010000010000000100010011;
ROM[2522] <= 32'b11111111110000010000000100010011;
ROM[2523] <= 32'b00000000000000010010001110000011;
ROM[2524] <= 32'b11111111110000010000000100010011;
ROM[2525] <= 32'b00000000000000010010010000000011;
ROM[2526] <= 32'b00000000100000111010001110110011;
ROM[2527] <= 32'b00000000011100010010000000100011;
ROM[2528] <= 32'b00000000010000010000000100010011;
ROM[2529] <= 32'b11111111110000010000000100010011;
ROM[2530] <= 32'b00000000000000010010001110000011;
ROM[2531] <= 32'b00000000000000111000101001100011;
ROM[2532] <= 32'b00000000000000000111001110110111;
ROM[2533] <= 32'b00101100100000111000001110010011;
ROM[2534] <= 32'b00000000111000111000001110110011;
ROM[2535] <= 32'b00000000000000111000000011100111;
ROM[2536] <= 32'b00111000010100000100000011101111;
ROM[2537] <= 32'b00000000000000100010001110000011;
ROM[2538] <= 32'b00000000011100010010000000100011;
ROM[2539] <= 32'b00000000010000010000000100010011;
ROM[2540] <= 32'b00000001010000000000001110010011;
ROM[2541] <= 32'b01000000011100011000001110110011;
ROM[2542] <= 32'b00000000000000111010000010000011;
ROM[2543] <= 32'b11111111110000010000000100010011;
ROM[2544] <= 32'b00000000000000010010001110000011;
ROM[2545] <= 32'b00000000011100100010000000100011;
ROM[2546] <= 32'b00000000010000100000000100010011;
ROM[2547] <= 32'b00000001010000000000001110010011;
ROM[2548] <= 32'b01000000011100011000001110110011;
ROM[2549] <= 32'b00000000010000111010000110000011;
ROM[2550] <= 32'b00000000100000111010001000000011;
ROM[2551] <= 32'b00000000110000111010001010000011;
ROM[2552] <= 32'b00000001000000111010001100000011;
ROM[2553] <= 32'b00000000000000001000000011100111;
ROM[2554] <= 32'b00111000000100000100000011101111;
ROM[2555] <= 32'b00000000010000100010001110000011;
ROM[2556] <= 32'b00000000011100010010000000100011;
ROM[2557] <= 32'b00000000010000010000000100010011;
ROM[2558] <= 32'b00000001010000000000001110010011;
ROM[2559] <= 32'b01000000011100011000001110110011;
ROM[2560] <= 32'b00000000000000111010000010000011;
ROM[2561] <= 32'b11111111110000010000000100010011;
ROM[2562] <= 32'b00000000000000010010001110000011;
ROM[2563] <= 32'b00000000011100100010000000100011;
ROM[2564] <= 32'b00000000010000100000000100010011;
ROM[2565] <= 32'b00000001010000000000001110010011;
ROM[2566] <= 32'b01000000011100011000001110110011;
ROM[2567] <= 32'b00000000010000111010000110000011;
ROM[2568] <= 32'b00000000100000111010001000000011;
ROM[2569] <= 32'b00000000110000111010001010000011;
ROM[2570] <= 32'b00000001000000111010001100000011;
ROM[2571] <= 32'b00000000000000001000000011100111;
ROM[2572] <= 32'b00000000000000100010001110000011;
ROM[2573] <= 32'b00000000011100010010000000100011;
ROM[2574] <= 32'b00000000010000010000000100010011;
ROM[2575] <= 32'b00000000010000100010001110000011;
ROM[2576] <= 32'b00000000011100010010000000100011;
ROM[2577] <= 32'b00000000010000010000000100010011;
ROM[2578] <= 32'b11111111110000010000000100010011;
ROM[2579] <= 32'b00000000000000010010001110000011;
ROM[2580] <= 32'b11111111110000010000000100010011;
ROM[2581] <= 32'b00000000000000010010010000000011;
ROM[2582] <= 32'b00000000011101000010001110110011;
ROM[2583] <= 32'b00000000011100010010000000100011;
ROM[2584] <= 32'b00000000010000010000000100010011;
ROM[2585] <= 32'b11111111110000010000000100010011;
ROM[2586] <= 32'b00000000000000010010001110000011;
ROM[2587] <= 32'b00000000000000111000101001100011;
ROM[2588] <= 32'b00000000000000000111001110110111;
ROM[2589] <= 32'b01011011010000111000001110010011;
ROM[2590] <= 32'b00000000111000111000001110110011;
ROM[2591] <= 32'b00000000000000111000000011100111;
ROM[2592] <= 32'b01011101000100000100000011101111;
ROM[2593] <= 32'b00000000000000100010001110000011;
ROM[2594] <= 32'b00000000011100010010000000100011;
ROM[2595] <= 32'b00000000010000010000000100010011;
ROM[2596] <= 32'b00000001010000000000001110010011;
ROM[2597] <= 32'b01000000011100011000001110110011;
ROM[2598] <= 32'b00000000000000111010000010000011;
ROM[2599] <= 32'b11111111110000010000000100010011;
ROM[2600] <= 32'b00000000000000010010001110000011;
ROM[2601] <= 32'b00000000011100100010000000100011;
ROM[2602] <= 32'b00000000010000100000000100010011;
ROM[2603] <= 32'b00000001010000000000001110010011;
ROM[2604] <= 32'b01000000011100011000001110110011;
ROM[2605] <= 32'b00000000010000111010000110000011;
ROM[2606] <= 32'b00000000100000111010001000000011;
ROM[2607] <= 32'b00000000110000111010001010000011;
ROM[2608] <= 32'b00000001000000111010001100000011;
ROM[2609] <= 32'b00000000000000001000000011100111;
ROM[2610] <= 32'b01011000100100000100000011101111;
ROM[2611] <= 32'b00000000010000100010001110000011;
ROM[2612] <= 32'b00000000011100010010000000100011;
ROM[2613] <= 32'b00000000010000010000000100010011;
ROM[2614] <= 32'b00000001010000000000001110010011;
ROM[2615] <= 32'b01000000011100011000001110110011;
ROM[2616] <= 32'b00000000000000111010000010000011;
ROM[2617] <= 32'b11111111110000010000000100010011;
ROM[2618] <= 32'b00000000000000010010001110000011;
ROM[2619] <= 32'b00000000011100100010000000100011;
ROM[2620] <= 32'b00000000010000100000000100010011;
ROM[2621] <= 32'b00000001010000000000001110010011;
ROM[2622] <= 32'b01000000011100011000001110110011;
ROM[2623] <= 32'b00000000010000111010000110000011;
ROM[2624] <= 32'b00000000100000111010001000000011;
ROM[2625] <= 32'b00000000110000111010001010000011;
ROM[2626] <= 32'b00000001000000111010001100000011;
ROM[2627] <= 32'b00000000000000001000000011100111;
ROM[2628] <= 32'b00000000000000100010001110000011;
ROM[2629] <= 32'b00000000011100010010000000100011;
ROM[2630] <= 32'b00000000010000010000000100010011;
ROM[2631] <= 32'b00000000000000100010001110000011;
ROM[2632] <= 32'b00000000011100010010000000100011;
ROM[2633] <= 32'b00000000010000010000000100010011;
ROM[2634] <= 32'b00000000010000100010001110000011;
ROM[2635] <= 32'b00000000011100010010000000100011;
ROM[2636] <= 32'b00000000010000010000000100010011;
ROM[2637] <= 32'b00000000000000000011001110110111;
ROM[2638] <= 32'b10011000000000111000001110010011;
ROM[2639] <= 32'b00000000111000111000001110110011;
ROM[2640] <= 32'b00000000011100010010000000100011;
ROM[2641] <= 32'b00000000010000010000000100010011;
ROM[2642] <= 32'b00000000001100010010000000100011;
ROM[2643] <= 32'b00000000010000010000000100010011;
ROM[2644] <= 32'b00000000010000010010000000100011;
ROM[2645] <= 32'b00000000010000010000000100010011;
ROM[2646] <= 32'b00000000010100010010000000100011;
ROM[2647] <= 32'b00000000010000010000000100010011;
ROM[2648] <= 32'b00000000011000010010000000100011;
ROM[2649] <= 32'b00000000010000010000000100010011;
ROM[2650] <= 32'b00000001010000000000001110010011;
ROM[2651] <= 32'b00000000100000111000001110010011;
ROM[2652] <= 32'b01000000011100010000001110110011;
ROM[2653] <= 32'b00000000011100000000001000110011;
ROM[2654] <= 32'b00000000001000000000000110110011;
ROM[2655] <= 32'b10010101000111111111000011101111;
ROM[2656] <= 32'b00000000010000100010001110000011;
ROM[2657] <= 32'b00000000011100010010000000100011;
ROM[2658] <= 32'b00000000010000010000000100010011;
ROM[2659] <= 32'b00000000000000000011001110110111;
ROM[2660] <= 32'b10011101100000111000001110010011;
ROM[2661] <= 32'b00000000111000111000001110110011;
ROM[2662] <= 32'b00000000011100010010000000100011;
ROM[2663] <= 32'b00000000010000010000000100010011;
ROM[2664] <= 32'b00000000001100010010000000100011;
ROM[2665] <= 32'b00000000010000010000000100010011;
ROM[2666] <= 32'b00000000010000010010000000100011;
ROM[2667] <= 32'b00000000010000010000000100010011;
ROM[2668] <= 32'b00000000010100010010000000100011;
ROM[2669] <= 32'b00000000010000010000000100010011;
ROM[2670] <= 32'b00000000011000010010000000100011;
ROM[2671] <= 32'b00000000010000010000000100010011;
ROM[2672] <= 32'b00000001010000000000001110010011;
ROM[2673] <= 32'b00000000100000111000001110010011;
ROM[2674] <= 32'b01000000011100010000001110110011;
ROM[2675] <= 32'b00000000011100000000001000110011;
ROM[2676] <= 32'b00000000001000000000000110110011;
ROM[2677] <= 32'b11010111010011111111000011101111;
ROM[2678] <= 32'b11111111110000010000000100010011;
ROM[2679] <= 32'b00000000000000010010001110000011;
ROM[2680] <= 32'b11111111110000010000000100010011;
ROM[2681] <= 32'b00000000000000010010010000000011;
ROM[2682] <= 32'b01000000011101000000001110110011;
ROM[2683] <= 32'b00000000011100010010000000100011;
ROM[2684] <= 32'b00000000010000010000000100010011;
ROM[2685] <= 32'b00000001010000000000001110010011;
ROM[2686] <= 32'b01000000011100011000001110110011;
ROM[2687] <= 32'b00000000000000111010000010000011;
ROM[2688] <= 32'b11111111110000010000000100010011;
ROM[2689] <= 32'b00000000000000010010001110000011;
ROM[2690] <= 32'b00000000011100100010000000100011;
ROM[2691] <= 32'b00000000010000100000000100010011;
ROM[2692] <= 32'b00000001010000000000001110010011;
ROM[2693] <= 32'b01000000011100011000001110110011;
ROM[2694] <= 32'b00000000010000111010000110000011;
ROM[2695] <= 32'b00000000100000111010001000000011;
ROM[2696] <= 32'b00000000110000111010001010000011;
ROM[2697] <= 32'b00000001000000111010001100000011;
ROM[2698] <= 32'b00000000000000001000000011100111;
ROM[2699] <= 32'b00000000000000100010001110000011;
ROM[2700] <= 32'b00000000011100010010000000100011;
ROM[2701] <= 32'b00000000010000010000000100010011;
ROM[2702] <= 32'b00000000010000000000001110010011;
ROM[2703] <= 32'b00000000011100010010000000100011;
ROM[2704] <= 32'b00000000010000010000000100010011;
ROM[2705] <= 32'b00000000000000000011001110110111;
ROM[2706] <= 32'b10101001000000111000001110010011;
ROM[2707] <= 32'b00000000111000111000001110110011;
ROM[2708] <= 32'b00000000011100010010000000100011;
ROM[2709] <= 32'b00000000010000010000000100010011;
ROM[2710] <= 32'b00000000001100010010000000100011;
ROM[2711] <= 32'b00000000010000010000000100010011;
ROM[2712] <= 32'b00000000010000010010000000100011;
ROM[2713] <= 32'b00000000010000010000000100010011;
ROM[2714] <= 32'b00000000010100010010000000100011;
ROM[2715] <= 32'b00000000010000010000000100010011;
ROM[2716] <= 32'b00000000011000010010000000100011;
ROM[2717] <= 32'b00000000010000010000000100010011;
ROM[2718] <= 32'b00000001010000000000001110010011;
ROM[2719] <= 32'b00000000100000111000001110010011;
ROM[2720] <= 32'b01000000011100010000001110110011;
ROM[2721] <= 32'b00000000011100000000001000110011;
ROM[2722] <= 32'b00000000001000000000000110110011;
ROM[2723] <= 32'b11001011110011111111000011101111;
ROM[2724] <= 32'b11111111110000010000000100010011;
ROM[2725] <= 32'b00000000000000010010001110000011;
ROM[2726] <= 32'b00000000011100100010000000100011;
ROM[2727] <= 32'b00000000000000100010001110000011;
ROM[2728] <= 32'b00000000011100010010000000100011;
ROM[2729] <= 32'b00000000010000010000000100010011;
ROM[2730] <= 32'b00000100000001101010001110000011;
ROM[2731] <= 32'b00000000011100010010000000100011;
ROM[2732] <= 32'b00000000010000010000000100010011;
ROM[2733] <= 32'b11111111110000010000000100010011;
ROM[2734] <= 32'b00000000000000010010001110000011;
ROM[2735] <= 32'b11111111110000010000000100010011;
ROM[2736] <= 32'b00000000000000010010010000000011;
ROM[2737] <= 32'b00000000011101000000001110110011;
ROM[2738] <= 32'b00000000011100010010000000100011;
ROM[2739] <= 32'b00000000010000010000000100010011;
ROM[2740] <= 32'b11111111110000010000000100010011;
ROM[2741] <= 32'b00000000000000010010001110000011;
ROM[2742] <= 32'b00000000000000111000001100010011;
ROM[2743] <= 32'b00000000110100110000010000110011;
ROM[2744] <= 32'b00000000000001000010001110000011;
ROM[2745] <= 32'b00000000011100010010000000100011;
ROM[2746] <= 32'b00000000010000010000000100010011;
ROM[2747] <= 32'b00000001010000000000001110010011;
ROM[2748] <= 32'b01000000011100011000001110110011;
ROM[2749] <= 32'b00000000000000111010000010000011;
ROM[2750] <= 32'b11111111110000010000000100010011;
ROM[2751] <= 32'b00000000000000010010001110000011;
ROM[2752] <= 32'b00000000011100100010000000100011;
ROM[2753] <= 32'b00000000010000100000000100010011;
ROM[2754] <= 32'b00000001010000000000001110010011;
ROM[2755] <= 32'b01000000011100011000001110110011;
ROM[2756] <= 32'b00000000010000111010000110000011;
ROM[2757] <= 32'b00000000100000111010001000000011;
ROM[2758] <= 32'b00000000110000111010001010000011;
ROM[2759] <= 32'b00000001000000111010001100000011;
ROM[2760] <= 32'b00000000000000001000000011100111;
ROM[2761] <= 32'b00000000000000000010001110110111;
ROM[2762] <= 32'b00000000000000111000001110010011;
ROM[2763] <= 32'b00000000011100010010000000100011;
ROM[2764] <= 32'b00000000010000010000000100010011;
ROM[2765] <= 32'b11111111110000010000000100010011;
ROM[2766] <= 32'b00000000000000010010001110000011;
ROM[2767] <= 32'b00000100011101101010001000100011;
ROM[2768] <= 32'b00000000000000000100001110110111;
ROM[2769] <= 32'b00000000000000111000001110010011;
ROM[2770] <= 32'b00000000011100010010000000100011;
ROM[2771] <= 32'b00000000010000010000000100010011;
ROM[2772] <= 32'b11111111110000010000000100010011;
ROM[2773] <= 32'b00000000000000010010001110000011;
ROM[2774] <= 32'b00000100011101101010010000100011;
ROM[2775] <= 32'b00000000000000000001001110110111;
ROM[2776] <= 32'b10000000000000111000001110010011;
ROM[2777] <= 32'b00000000011100010010000000100011;
ROM[2778] <= 32'b00000000010000010000000100010011;
ROM[2779] <= 32'b11111111110000010000000100010011;
ROM[2780] <= 32'b00000000000000010010001110000011;
ROM[2781] <= 32'b00000100011101101010011000100011;
ROM[2782] <= 32'b00000000000000000100001110110111;
ROM[2783] <= 32'b00000000000000111000001110010011;
ROM[2784] <= 32'b00000000011100010010000000100011;
ROM[2785] <= 32'b00000000010000010000000100010011;
ROM[2786] <= 32'b11111111110000010000000100010011;
ROM[2787] <= 32'b00000000000000010010001110000011;
ROM[2788] <= 32'b00000100011101101010100000100011;
ROM[2789] <= 32'b00000000000000000000001110010011;
ROM[2790] <= 32'b00000000011100010010000000100011;
ROM[2791] <= 32'b00000000010000010000000100010011;
ROM[2792] <= 32'b11111111110000010000000100010011;
ROM[2793] <= 32'b00000000000000010010001110000011;
ROM[2794] <= 32'b00000100011101101010101000100011;
ROM[2795] <= 32'b00000100010001101010001110000011;
ROM[2796] <= 32'b00000000011100010010000000100011;
ROM[2797] <= 32'b00000000010000010000000100010011;
ROM[2798] <= 32'b11111111110000010000000100010011;
ROM[2799] <= 32'b00000000000000010010001110000011;
ROM[2800] <= 32'b00000100011101101010110000100011;
ROM[2801] <= 32'b00000000000000000000001110010011;
ROM[2802] <= 32'b00000000011100010010000000100011;
ROM[2803] <= 32'b00000000010000010000000100010011;
ROM[2804] <= 32'b11111111110000010000000100010011;
ROM[2805] <= 32'b00000000000000010010001110000011;
ROM[2806] <= 32'b00000100011101101010111000100011;
ROM[2807] <= 32'b00000000010000000000001110010011;
ROM[2808] <= 32'b00000000011100010010000000100011;
ROM[2809] <= 32'b00000000010000010000000100010011;
ROM[2810] <= 32'b11111111110000010000000100010011;
ROM[2811] <= 32'b00000000000000010010001110000011;
ROM[2812] <= 32'b00000110011101101010000000100011;
ROM[2813] <= 32'b00000101110001101010001110000011;
ROM[2814] <= 32'b00000000011100010010000000100011;
ROM[2815] <= 32'b00000000010000010000000100010011;
ROM[2816] <= 32'b00000101100001101010001110000011;
ROM[2817] <= 32'b00000000011100010010000000100011;
ROM[2818] <= 32'b00000000010000010000000100010011;
ROM[2819] <= 32'b11111111110000010000000100010011;
ROM[2820] <= 32'b00000000000000010010001110000011;
ROM[2821] <= 32'b11111111110000010000000100010011;
ROM[2822] <= 32'b00000000000000010010010000000011;
ROM[2823] <= 32'b00000000011101000000001110110011;
ROM[2824] <= 32'b00000000011100010010000000100011;
ROM[2825] <= 32'b00000000010000010000000100010011;
ROM[2826] <= 32'b00000101000001101010001110000011;
ROM[2827] <= 32'b00000000011100010010000000100011;
ROM[2828] <= 32'b00000000010000010000000100010011;
ROM[2829] <= 32'b00000100110001101010001110000011;
ROM[2830] <= 32'b00000000011100010010000000100011;
ROM[2831] <= 32'b00000000010000010000000100010011;
ROM[2832] <= 32'b11111111110000010000000100010011;
ROM[2833] <= 32'b00000000000000010010001110000011;
ROM[2834] <= 32'b11111111110000010000000100010011;
ROM[2835] <= 32'b00000000000000010010010000000011;
ROM[2836] <= 32'b01000000011101000000001110110011;
ROM[2837] <= 32'b00000000011100010010000000100011;
ROM[2838] <= 32'b00000000010000010000000100010011;
ROM[2839] <= 32'b11111111110000010000000100010011;
ROM[2840] <= 32'b00000000000000010010001110000011;
ROM[2841] <= 32'b00000000011101100010000000100011;
ROM[2842] <= 32'b11111111110000010000000100010011;
ROM[2843] <= 32'b00000000000000010010001110000011;
ROM[2844] <= 32'b00000000000000111000001100010011;
ROM[2845] <= 32'b00000000000001100010001110000011;
ROM[2846] <= 32'b00000000011100010010000000100011;
ROM[2847] <= 32'b00000000010000010000000100010011;
ROM[2848] <= 32'b11111111110000010000000100010011;
ROM[2849] <= 32'b00000000000000010010001110000011;
ROM[2850] <= 32'b00000000110100110000010000110011;
ROM[2851] <= 32'b00000000011101000010000000100011;
ROM[2852] <= 32'b00000110000001101010001110000011;
ROM[2853] <= 32'b00000000011100010010000000100011;
ROM[2854] <= 32'b00000000010000010000000100010011;
ROM[2855] <= 32'b00000101100001101010001110000011;
ROM[2856] <= 32'b00000000011100010010000000100011;
ROM[2857] <= 32'b00000000010000010000000100010011;
ROM[2858] <= 32'b11111111110000010000000100010011;
ROM[2859] <= 32'b00000000000000010010001110000011;
ROM[2860] <= 32'b11111111110000010000000100010011;
ROM[2861] <= 32'b00000000000000010010010000000011;
ROM[2862] <= 32'b00000000011101000000001110110011;
ROM[2863] <= 32'b00000000011100010010000000100011;
ROM[2864] <= 32'b00000000010000010000000100010011;
ROM[2865] <= 32'b00000000000000000000001110010011;
ROM[2866] <= 32'b00000000011100010010000000100011;
ROM[2867] <= 32'b00000000010000010000000100010011;
ROM[2868] <= 32'b11111111110000010000000100010011;
ROM[2869] <= 32'b00000000000000010010001110000011;
ROM[2870] <= 32'b00000000011101100010000000100011;
ROM[2871] <= 32'b11111111110000010000000100010011;
ROM[2872] <= 32'b00000000000000010010001110000011;
ROM[2873] <= 32'b00000000000000111000001100010011;
ROM[2874] <= 32'b00000000000001100010001110000011;
ROM[2875] <= 32'b00000000011100010010000000100011;
ROM[2876] <= 32'b00000000010000010000000100010011;
ROM[2877] <= 32'b11111111110000010000000100010011;
ROM[2878] <= 32'b00000000000000010010001110000011;
ROM[2879] <= 32'b00000000110100110000010000110011;
ROM[2880] <= 32'b00000000011101000010000000100011;
ROM[2881] <= 32'b00000000010000000000001110010011;
ROM[2882] <= 32'b00000000011100010010000000100011;
ROM[2883] <= 32'b00000000010000010000000100010011;
ROM[2884] <= 32'b11111111110000010000000100010011;
ROM[2885] <= 32'b00000000000000010010001110000011;
ROM[2886] <= 32'b01000000011100000000001110110011;
ROM[2887] <= 32'b00000000011100010010000000100011;
ROM[2888] <= 32'b00000000010000010000000100010011;
ROM[2889] <= 32'b11111111110000010000000100010011;
ROM[2890] <= 32'b00000000000000010010001110000011;
ROM[2891] <= 32'b00000110011101101010001000100011;
ROM[2892] <= 32'b00000000000000000000001110010011;
ROM[2893] <= 32'b00000000011100010010000000100011;
ROM[2894] <= 32'b00000000010000010000000100010011;
ROM[2895] <= 32'b00000001010000000000001110010011;
ROM[2896] <= 32'b01000000011100011000001110110011;
ROM[2897] <= 32'b00000000000000111010000010000011;
ROM[2898] <= 32'b11111111110000010000000100010011;
ROM[2899] <= 32'b00000000000000010010001110000011;
ROM[2900] <= 32'b00000000011100100010000000100011;
ROM[2901] <= 32'b00000000010000100000000100010011;
ROM[2902] <= 32'b00000001010000000000001110010011;
ROM[2903] <= 32'b01000000011100011000001110110011;
ROM[2904] <= 32'b00000000010000111010000110000011;
ROM[2905] <= 32'b00000000100000111010001000000011;
ROM[2906] <= 32'b00000000110000111010001010000011;
ROM[2907] <= 32'b00000001000000111010001100000011;
ROM[2908] <= 32'b00000000000000001000000011100111;
ROM[2909] <= 32'b00000000000000100010001110000011;
ROM[2910] <= 32'b00000000011100010010000000100011;
ROM[2911] <= 32'b00000000010000010000000100010011;
ROM[2912] <= 32'b00000000000000100010001110000011;
ROM[2913] <= 32'b00000000011100010010000000100011;
ROM[2914] <= 32'b00000000010000010000000100010011;
ROM[2915] <= 32'b11111111110000010000000100010011;
ROM[2916] <= 32'b00000000000000010010001110000011;
ROM[2917] <= 32'b11111111110000010000000100010011;
ROM[2918] <= 32'b00000000000000010010010000000011;
ROM[2919] <= 32'b00000000011101000000001110110011;
ROM[2920] <= 32'b00000000011100010010000000100011;
ROM[2921] <= 32'b00000000010000010000000100010011;
ROM[2922] <= 32'b11111111110000010000000100010011;
ROM[2923] <= 32'b00000000000000010010001110000011;
ROM[2924] <= 32'b00000000011100100010000000100011;
ROM[2925] <= 32'b00000000000000100010001110000011;
ROM[2926] <= 32'b00000000011100010010000000100011;
ROM[2927] <= 32'b00000000010000010000000100010011;
ROM[2928] <= 32'b00000000000000100010001110000011;
ROM[2929] <= 32'b00000000011100010010000000100011;
ROM[2930] <= 32'b00000000010000010000000100010011;
ROM[2931] <= 32'b11111111110000010000000100010011;
ROM[2932] <= 32'b00000000000000010010001110000011;
ROM[2933] <= 32'b11111111110000010000000100010011;
ROM[2934] <= 32'b00000000000000010010010000000011;
ROM[2935] <= 32'b00000000011101000000001110110011;
ROM[2936] <= 32'b00000000011100010010000000100011;
ROM[2937] <= 32'b00000000010000010000000100010011;
ROM[2938] <= 32'b11111111110000010000000100010011;
ROM[2939] <= 32'b00000000000000010010001110000011;
ROM[2940] <= 32'b00000000011100100010000000100011;
ROM[2941] <= 32'b00000000000000100010001110000011;
ROM[2942] <= 32'b00000000011100010010000000100011;
ROM[2943] <= 32'b00000000010000010000000100010011;
ROM[2944] <= 32'b00000101010001101010001110000011;
ROM[2945] <= 32'b00000000011100010010000000100011;
ROM[2946] <= 32'b00000000010000010000000100010011;
ROM[2947] <= 32'b11111111110000010000000100010011;
ROM[2948] <= 32'b00000000000000010010001110000011;
ROM[2949] <= 32'b11111111110000010000000100010011;
ROM[2950] <= 32'b00000000000000010010010000000011;
ROM[2951] <= 32'b00000000011101000000001110110011;
ROM[2952] <= 32'b00000000011100010010000000100011;
ROM[2953] <= 32'b00000000010000010000000100010011;
ROM[2954] <= 32'b11111111110000010000000100010011;
ROM[2955] <= 32'b00000000000000010010001110000011;
ROM[2956] <= 32'b00000000000000111000001100010011;
ROM[2957] <= 32'b00000000110100110000010000110011;
ROM[2958] <= 32'b00000000000001000010001110000011;
ROM[2959] <= 32'b00000000011100010010000000100011;
ROM[2960] <= 32'b00000000010000010000000100010011;
ROM[2961] <= 32'b00000001010000000000001110010011;
ROM[2962] <= 32'b01000000011100011000001110110011;
ROM[2963] <= 32'b00000000000000111010000010000011;
ROM[2964] <= 32'b11111111110000010000000100010011;
ROM[2965] <= 32'b00000000000000010010001110000011;
ROM[2966] <= 32'b00000000011100100010000000100011;
ROM[2967] <= 32'b00000000010000100000000100010011;
ROM[2968] <= 32'b00000001010000000000001110010011;
ROM[2969] <= 32'b01000000011100011000001110110011;
ROM[2970] <= 32'b00000000010000111010000110000011;
ROM[2971] <= 32'b00000000100000111010001000000011;
ROM[2972] <= 32'b00000000110000111010001010000011;
ROM[2973] <= 32'b00000001000000111010001100000011;
ROM[2974] <= 32'b00000000000000001000000011100111;
ROM[2975] <= 32'b00000000000000100010001110000011;
ROM[2976] <= 32'b00000000011100010010000000100011;
ROM[2977] <= 32'b00000000010000010000000100010011;
ROM[2978] <= 32'b00000000000000100010001110000011;
ROM[2979] <= 32'b00000000011100010010000000100011;
ROM[2980] <= 32'b00000000010000010000000100010011;
ROM[2981] <= 32'b11111111110000010000000100010011;
ROM[2982] <= 32'b00000000000000010010001110000011;
ROM[2983] <= 32'b11111111110000010000000100010011;
ROM[2984] <= 32'b00000000000000010010010000000011;
ROM[2985] <= 32'b00000000011101000000001110110011;
ROM[2986] <= 32'b00000000011100010010000000100011;
ROM[2987] <= 32'b00000000010000010000000100010011;
ROM[2988] <= 32'b11111111110000010000000100010011;
ROM[2989] <= 32'b00000000000000010010001110000011;
ROM[2990] <= 32'b00000000011100100010000000100011;
ROM[2991] <= 32'b00000000000000100010001110000011;
ROM[2992] <= 32'b00000000011100010010000000100011;
ROM[2993] <= 32'b00000000010000010000000100010011;
ROM[2994] <= 32'b00000000000000100010001110000011;
ROM[2995] <= 32'b00000000011100010010000000100011;
ROM[2996] <= 32'b00000000010000010000000100010011;
ROM[2997] <= 32'b11111111110000010000000100010011;
ROM[2998] <= 32'b00000000000000010010001110000011;
ROM[2999] <= 32'b11111111110000010000000100010011;
ROM[3000] <= 32'b00000000000000010010010000000011;
ROM[3001] <= 32'b00000000011101000000001110110011;
ROM[3002] <= 32'b00000000011100010010000000100011;
ROM[3003] <= 32'b00000000010000010000000100010011;
ROM[3004] <= 32'b11111111110000010000000100010011;
ROM[3005] <= 32'b00000000000000010010001110000011;
ROM[3006] <= 32'b00000000011100100010000000100011;
ROM[3007] <= 32'b00000000000000100010001110000011;
ROM[3008] <= 32'b00000000011100010010000000100011;
ROM[3009] <= 32'b00000000010000010000000100010011;
ROM[3010] <= 32'b00000101010001101010001110000011;
ROM[3011] <= 32'b00000000011100010010000000100011;
ROM[3012] <= 32'b00000000010000010000000100010011;
ROM[3013] <= 32'b11111111110000010000000100010011;
ROM[3014] <= 32'b00000000000000010010001110000011;
ROM[3015] <= 32'b11111111110000010000000100010011;
ROM[3016] <= 32'b00000000000000010010010000000011;
ROM[3017] <= 32'b00000000011101000000001110110011;
ROM[3018] <= 32'b00000000011100010010000000100011;
ROM[3019] <= 32'b00000000010000010000000100010011;
ROM[3020] <= 32'b00000000010000100010001110000011;
ROM[3021] <= 32'b00000000011100010010000000100011;
ROM[3022] <= 32'b00000000010000010000000100010011;
ROM[3023] <= 32'b11111111110000010000000100010011;
ROM[3024] <= 32'b00000000000000010010001110000011;
ROM[3025] <= 32'b00000000011101100010000000100011;
ROM[3026] <= 32'b11111111110000010000000100010011;
ROM[3027] <= 32'b00000000000000010010001110000011;
ROM[3028] <= 32'b00000000000000111000001100010011;
ROM[3029] <= 32'b00000000000001100010001110000011;
ROM[3030] <= 32'b00000000011100010010000000100011;
ROM[3031] <= 32'b00000000010000010000000100010011;
ROM[3032] <= 32'b11111111110000010000000100010011;
ROM[3033] <= 32'b00000000000000010010001110000011;
ROM[3034] <= 32'b00000000110100110000010000110011;
ROM[3035] <= 32'b00000000011101000010000000100011;
ROM[3036] <= 32'b00000000000000000000001110010011;
ROM[3037] <= 32'b00000000011100010010000000100011;
ROM[3038] <= 32'b00000000010000010000000100010011;
ROM[3039] <= 32'b00000001010000000000001110010011;
ROM[3040] <= 32'b01000000011100011000001110110011;
ROM[3041] <= 32'b00000000000000111010000010000011;
ROM[3042] <= 32'b11111111110000010000000100010011;
ROM[3043] <= 32'b00000000000000010010001110000011;
ROM[3044] <= 32'b00000000011100100010000000100011;
ROM[3045] <= 32'b00000000010000100000000100010011;
ROM[3046] <= 32'b00000001010000000000001110010011;
ROM[3047] <= 32'b01000000011100011000001110110011;
ROM[3048] <= 32'b00000000010000111010000110000011;
ROM[3049] <= 32'b00000000100000111010001000000011;
ROM[3050] <= 32'b00000000110000111010001010000011;
ROM[3051] <= 32'b00000001000000111010001100000011;
ROM[3052] <= 32'b00000000000000001000000011100111;
ROM[3053] <= 32'b00000000000000010010000000100011;
ROM[3054] <= 32'b00000000010000010000000100010011;
ROM[3055] <= 32'b00000000000000010010000000100011;
ROM[3056] <= 32'b00000000010000010000000100010011;
ROM[3057] <= 32'b00000000000000010010000000100011;
ROM[3058] <= 32'b00000000010000010000000100010011;
ROM[3059] <= 32'b00000000000000010010000000100011;
ROM[3060] <= 32'b00000000010000010000000100010011;
ROM[3061] <= 32'b00000000000000000000001110010011;
ROM[3062] <= 32'b00000000011100010010000000100011;
ROM[3063] <= 32'b00000000010000010000000100010011;
ROM[3064] <= 32'b11111111110000010000000100010011;
ROM[3065] <= 32'b00000000000000010010001110000011;
ROM[3066] <= 32'b00000000011100011010001000100011;
ROM[3067] <= 32'b00000101000001101010001110000011;
ROM[3068] <= 32'b00000000011100010010000000100011;
ROM[3069] <= 32'b00000000010000010000000100010011;
ROM[3070] <= 32'b00000100110001101010001110000011;
ROM[3071] <= 32'b00000000011100010010000000100011;
ROM[3072] <= 32'b00000000010000010000000100010011;
ROM[3073] <= 32'b11111111110000010000000100010011;
ROM[3074] <= 32'b00000000000000010010001110000011;
ROM[3075] <= 32'b11111111110000010000000100010011;
ROM[3076] <= 32'b00000000000000010010010000000011;
ROM[3077] <= 32'b01000000011101000000001110110011;
ROM[3078] <= 32'b00000000011100010010000000100011;
ROM[3079] <= 32'b00000000010000010000000100010011;
ROM[3080] <= 32'b11111111110000010000000100010011;
ROM[3081] <= 32'b00000000000000010010001110000011;
ROM[3082] <= 32'b00000000011100011010010000100011;
ROM[3083] <= 32'b00000101100001101010001110000011;
ROM[3084] <= 32'b00000000011100010010000000100011;
ROM[3085] <= 32'b00000000010000010000000100010011;
ROM[3086] <= 32'b11111111110000010000000100010011;
ROM[3087] <= 32'b00000000000000010010001110000011;
ROM[3088] <= 32'b00000000011100011010000000100011;
ROM[3089] <= 32'b00000110000001101010001110000011;
ROM[3090] <= 32'b00000000011100010010000000100011;
ROM[3091] <= 32'b00000000010000010000000100010011;
ROM[3092] <= 32'b00000000000000011010001110000011;
ROM[3093] <= 32'b00000000011100010010000000100011;
ROM[3094] <= 32'b00000000010000010000000100010011;
ROM[3095] <= 32'b11111111110000010000000100010011;
ROM[3096] <= 32'b00000000000000010010001110000011;
ROM[3097] <= 32'b11111111110000010000000100010011;
ROM[3098] <= 32'b00000000000000010010010000000011;
ROM[3099] <= 32'b00000000011101000000001110110011;
ROM[3100] <= 32'b00000000011100010010000000100011;
ROM[3101] <= 32'b00000000010000010000000100010011;
ROM[3102] <= 32'b11111111110000010000000100010011;
ROM[3103] <= 32'b00000000000000010010001110000011;
ROM[3104] <= 32'b00000000000000111000001100010011;
ROM[3105] <= 32'b00000000110100110000010000110011;
ROM[3106] <= 32'b00000000000001000010001110000011;
ROM[3107] <= 32'b00000000011100010010000000100011;
ROM[3108] <= 32'b00000000010000010000000100010011;
ROM[3109] <= 32'b00000000000000000000001110010011;
ROM[3110] <= 32'b00000000011100010010000000100011;
ROM[3111] <= 32'b00000000010000010000000100010011;
ROM[3112] <= 32'b11111111110000010000000100010011;
ROM[3113] <= 32'b00000000000000010010001110000011;
ROM[3114] <= 32'b11111111110000010000000100010011;
ROM[3115] <= 32'b00000000000000010010010000000011;
ROM[3116] <= 32'b00000000011101000010010010110011;
ROM[3117] <= 32'b00000000100000111010010100110011;
ROM[3118] <= 32'b00000000101001001000001110110011;
ROM[3119] <= 32'b00000000000100111000001110010011;
ROM[3120] <= 32'b00000000000100111111001110010011;
ROM[3121] <= 32'b00000000011100010010000000100011;
ROM[3122] <= 32'b00000000010000010000000100010011;
ROM[3123] <= 32'b11111111110000010000000100010011;
ROM[3124] <= 32'b00000000000000010010001110000011;
ROM[3125] <= 32'b00000000000000111000101001100011;
ROM[3126] <= 32'b00000000000000000111001110110111;
ROM[3127] <= 32'b10001110100000111000001110010011;
ROM[3128] <= 32'b00000000111000111000001110110011;
ROM[3129] <= 32'b00000000000000111000000011100111;
ROM[3130] <= 32'b00000001110100000011000011101111;
ROM[3131] <= 32'b00000000000000011010001110000011;
ROM[3132] <= 32'b00000000011100010010000000100011;
ROM[3133] <= 32'b00000000010000010000000100010011;
ROM[3134] <= 32'b00000001010000000000001110010011;
ROM[3135] <= 32'b01000000011100011000001110110011;
ROM[3136] <= 32'b00000000000000111010000010000011;
ROM[3137] <= 32'b11111111110000010000000100010011;
ROM[3138] <= 32'b00000000000000010010001110000011;
ROM[3139] <= 32'b00000000011100100010000000100011;
ROM[3140] <= 32'b00000000010000100000000100010011;
ROM[3141] <= 32'b00000001010000000000001110010011;
ROM[3142] <= 32'b01000000011100011000001110110011;
ROM[3143] <= 32'b00000000010000111010000110000011;
ROM[3144] <= 32'b00000000100000111010001000000011;
ROM[3145] <= 32'b00000000110000111010001010000011;
ROM[3146] <= 32'b00000001000000111010001100000011;
ROM[3147] <= 32'b00000000000000001000000011100111;
ROM[3148] <= 32'b01111101010000000011000011101111;
ROM[3149] <= 32'b00000000000000011010001110000011;
ROM[3150] <= 32'b00000000011100010010000000100011;
ROM[3151] <= 32'b00000000010000010000000100010011;
ROM[3152] <= 32'b00000000000000000000001110010011;
ROM[3153] <= 32'b00000000011100010010000000100011;
ROM[3154] <= 32'b00000000010000010000000100010011;
ROM[3155] <= 32'b11111111110000010000000100010011;
ROM[3156] <= 32'b00000000000000010010001110000011;
ROM[3157] <= 32'b11111111110000010000000100010011;
ROM[3158] <= 32'b00000000000000010010010000000011;
ROM[3159] <= 32'b00000000011101000010010010110011;
ROM[3160] <= 32'b00000000100000111010010100110011;
ROM[3161] <= 32'b00000000101001001000001110110011;
ROM[3162] <= 32'b00000000000100111000001110010011;
ROM[3163] <= 32'b00000000000100111111001110010011;
ROM[3164] <= 32'b00000000011100010010000000100011;
ROM[3165] <= 32'b00000000010000010000000100010011;
ROM[3166] <= 32'b11111111110000010000000100010011;
ROM[3167] <= 32'b00000000000000010010001110000011;
ROM[3168] <= 32'b01000000011100000000001110110011;
ROM[3169] <= 32'b00000000000100111000001110010011;
ROM[3170] <= 32'b00000000011100010010000000100011;
ROM[3171] <= 32'b00000000010000010000000100010011;
ROM[3172] <= 32'b11111111110000010000000100010011;
ROM[3173] <= 32'b00000000000000010010001110000011;
ROM[3174] <= 32'b01000000011100000000001110110011;
ROM[3175] <= 32'b00000000000100111000001110010011;
ROM[3176] <= 32'b00000000011100010010000000100011;
ROM[3177] <= 32'b00000000010000010000000100010011;
ROM[3178] <= 32'b11111111110000010000000100010011;
ROM[3179] <= 32'b00000000000000010010001110000011;
ROM[3180] <= 32'b00000000000000111000101001100011;
ROM[3181] <= 32'b00000000000000001000001110110111;
ROM[3182] <= 32'b11001110010000111000001110010011;
ROM[3183] <= 32'b00000000111000111000001110110011;
ROM[3184] <= 32'b00000000000000111000000011100111;
ROM[3185] <= 32'b00000101110001101010001110000011;
ROM[3186] <= 32'b00000000011100010010000000100011;
ROM[3187] <= 32'b00000000010000010000000100010011;
ROM[3188] <= 32'b00000000000000011010001110000011;
ROM[3189] <= 32'b00000000011100010010000000100011;
ROM[3190] <= 32'b00000000010000010000000100010011;
ROM[3191] <= 32'b11111111110000010000000100010011;
ROM[3192] <= 32'b00000000000000010010001110000011;
ROM[3193] <= 32'b11111111110000010000000100010011;
ROM[3194] <= 32'b00000000000000010010010000000011;
ROM[3195] <= 32'b00000000011101000000001110110011;
ROM[3196] <= 32'b00000000011100010010000000100011;
ROM[3197] <= 32'b00000000010000010000000100010011;
ROM[3198] <= 32'b11111111110000010000000100010011;
ROM[3199] <= 32'b00000000000000010010001110000011;
ROM[3200] <= 32'b00000000000000111000001100010011;
ROM[3201] <= 32'b00000000110100110000010000110011;
ROM[3202] <= 32'b00000000000001000010001110000011;
ROM[3203] <= 32'b00000000011100010010000000100011;
ROM[3204] <= 32'b00000000010000010000000100010011;
ROM[3205] <= 32'b00000000000100000000001110010011;
ROM[3206] <= 32'b00000000011100010010000000100011;
ROM[3207] <= 32'b00000000010000010000000100010011;
ROM[3208] <= 32'b11111111110000010000000100010011;
ROM[3209] <= 32'b00000000000000010010001110000011;
ROM[3210] <= 32'b11111111110000010000000100010011;
ROM[3211] <= 32'b00000000000000010010010000000011;
ROM[3212] <= 32'b01000000011101000000001110110011;
ROM[3213] <= 32'b00000000011100010010000000100011;
ROM[3214] <= 32'b00000000010000010000000100010011;
ROM[3215] <= 32'b11111111110000010000000100010011;
ROM[3216] <= 32'b00000000000000010010001110000011;
ROM[3217] <= 32'b00000000011100011010011000100011;
ROM[3218] <= 32'b00000000110000011010001110000011;
ROM[3219] <= 32'b00000000011100010010000000100011;
ROM[3220] <= 32'b00000000010000010000000100010011;
ROM[3221] <= 32'b00000000000000100010001110000011;
ROM[3222] <= 32'b00000000011100010010000000100011;
ROM[3223] <= 32'b00000000010000010000000100010011;
ROM[3224] <= 32'b11111111110000010000000100010011;
ROM[3225] <= 32'b00000000000000010010001110000011;
ROM[3226] <= 32'b11111111110000010000000100010011;
ROM[3227] <= 32'b00000000000000010010010000000011;
ROM[3228] <= 32'b00000000011101000010001110110011;
ROM[3229] <= 32'b00000000011100010010000000100011;
ROM[3230] <= 32'b00000000010000010000000100010011;
ROM[3231] <= 32'b11111111110000010000000100010011;
ROM[3232] <= 32'b00000000000000010010001110000011;
ROM[3233] <= 32'b01000000011100000000001110110011;
ROM[3234] <= 32'b00000000000100111000001110010011;
ROM[3235] <= 32'b00000000011100010010000000100011;
ROM[3236] <= 32'b00000000010000010000000100010011;
ROM[3237] <= 32'b00000000110000011010001110000011;
ROM[3238] <= 32'b00000000011100010010000000100011;
ROM[3239] <= 32'b00000000010000010000000100010011;
ROM[3240] <= 32'b00000000100000011010001110000011;
ROM[3241] <= 32'b00000000011100010010000000100011;
ROM[3242] <= 32'b00000000010000010000000100010011;
ROM[3243] <= 32'b11111111110000010000000100010011;
ROM[3244] <= 32'b00000000000000010010001110000011;
ROM[3245] <= 32'b11111111110000010000000100010011;
ROM[3246] <= 32'b00000000000000010010010000000011;
ROM[3247] <= 32'b00000000011101000010001110110011;
ROM[3248] <= 32'b00000000011100010010000000100011;
ROM[3249] <= 32'b00000000010000010000000100010011;
ROM[3250] <= 32'b11111111110000010000000100010011;
ROM[3251] <= 32'b00000000000000010010001110000011;
ROM[3252] <= 32'b11111111110000010000000100010011;
ROM[3253] <= 32'b00000000000000010010010000000011;
ROM[3254] <= 32'b00000000011101000111001110110011;
ROM[3255] <= 32'b00000000011100010010000000100011;
ROM[3256] <= 32'b00000000010000010000000100010011;
ROM[3257] <= 32'b11111111110000010000000100010011;
ROM[3258] <= 32'b00000000000000010010001110000011;
ROM[3259] <= 32'b00000000000000111000101001100011;
ROM[3260] <= 32'b00000000000000000111001110110111;
ROM[3261] <= 32'b11000011000000111000001110010011;
ROM[3262] <= 32'b00000000111000111000001110110011;
ROM[3263] <= 32'b00000000000000111000000011100111;
ROM[3264] <= 32'b00011111100100000011000011101111;
ROM[3265] <= 32'b00000000000000011010001110000011;
ROM[3266] <= 32'b00000000011100010010000000100011;
ROM[3267] <= 32'b00000000010000010000000100010011;
ROM[3268] <= 32'b11111111110000010000000100010011;
ROM[3269] <= 32'b00000000000000010010001110000011;
ROM[3270] <= 32'b00000000011100011010001000100011;
ROM[3271] <= 32'b00000000110000011010001110000011;
ROM[3272] <= 32'b00000000011100010010000000100011;
ROM[3273] <= 32'b00000000010000010000000100010011;
ROM[3274] <= 32'b11111111110000010000000100010011;
ROM[3275] <= 32'b00000000000000010010001110000011;
ROM[3276] <= 32'b00000000011100011010010000100011;
ROM[3277] <= 32'b00011100010100000011000011101111;
ROM[3278] <= 32'b00000110000001101010001110000011;
ROM[3279] <= 32'b00000000011100010010000000100011;
ROM[3280] <= 32'b00000000010000010000000100010011;
ROM[3281] <= 32'b00000000000000011010001110000011;
ROM[3282] <= 32'b00000000011100010010000000100011;
ROM[3283] <= 32'b00000000010000010000000100010011;
ROM[3284] <= 32'b11111111110000010000000100010011;
ROM[3285] <= 32'b00000000000000010010001110000011;
ROM[3286] <= 32'b11111111110000010000000100010011;
ROM[3287] <= 32'b00000000000000010010010000000011;
ROM[3288] <= 32'b00000000011101000000001110110011;
ROM[3289] <= 32'b00000000011100010010000000100011;
ROM[3290] <= 32'b00000000010000010000000100010011;
ROM[3291] <= 32'b11111111110000010000000100010011;
ROM[3292] <= 32'b00000000000000010010001110000011;
ROM[3293] <= 32'b00000000000000111000001100010011;
ROM[3294] <= 32'b00000000110100110000010000110011;
ROM[3295] <= 32'b00000000000001000010001110000011;
ROM[3296] <= 32'b00000000011100010010000000100011;
ROM[3297] <= 32'b00000000010000010000000100010011;
ROM[3298] <= 32'b11111111110000010000000100010011;
ROM[3299] <= 32'b00000000000000010010001110000011;
ROM[3300] <= 32'b00000000011100011010000000100011;
ROM[3301] <= 32'b00001111010100000100000011101111;
ROM[3302] <= 32'b00000000010000011010001110000011;
ROM[3303] <= 32'b00000000011100010010000000100011;
ROM[3304] <= 32'b00000000010000010000000100010011;
ROM[3305] <= 32'b00000001010000000000001110010011;
ROM[3306] <= 32'b01000000011100011000001110110011;
ROM[3307] <= 32'b00000000000000111010000010000011;
ROM[3308] <= 32'b11111111110000010000000100010011;
ROM[3309] <= 32'b00000000000000010010001110000011;
ROM[3310] <= 32'b00000000011100100010000000100011;
ROM[3311] <= 32'b00000000010000100000000100010011;
ROM[3312] <= 32'b00000001010000000000001110010011;
ROM[3313] <= 32'b01000000011100011000001110110011;
ROM[3314] <= 32'b00000000010000111010000110000011;
ROM[3315] <= 32'b00000000100000111010001000000011;
ROM[3316] <= 32'b00000000110000111010001010000011;
ROM[3317] <= 32'b00000001000000111010001100000011;
ROM[3318] <= 32'b00000000000000001000000011100111;
ROM[3319] <= 32'b00000000000000010010000000100011;
ROM[3320] <= 32'b00000000010000010000000100010011;
ROM[3321] <= 32'b00000000000000010010000000100011;
ROM[3322] <= 32'b00000000010000010000000100010011;
ROM[3323] <= 32'b00000000000000010010000000100011;
ROM[3324] <= 32'b00000000010000010000000100010011;
ROM[3325] <= 32'b00000000000000100010001110000011;
ROM[3326] <= 32'b00000000011100010010000000100011;
ROM[3327] <= 32'b00000000010000010000000100010011;
ROM[3328] <= 32'b00000000000000000011001110110111;
ROM[3329] <= 32'b01000100110000111000001110010011;
ROM[3330] <= 32'b00000000111000111000001110110011;
ROM[3331] <= 32'b00000000011100010010000000100011;
ROM[3332] <= 32'b00000000010000010000000100010011;
ROM[3333] <= 32'b00000000001100010010000000100011;
ROM[3334] <= 32'b00000000010000010000000100010011;
ROM[3335] <= 32'b00000000010000010010000000100011;
ROM[3336] <= 32'b00000000010000010000000100010011;
ROM[3337] <= 32'b00000000010100010010000000100011;
ROM[3338] <= 32'b00000000010000010000000100010011;
ROM[3339] <= 32'b00000000011000010010000000100011;
ROM[3340] <= 32'b00000000010000010000000100010011;
ROM[3341] <= 32'b00000001010000000000001110010011;
ROM[3342] <= 32'b00000000010000111000001110010011;
ROM[3343] <= 32'b01000000011100010000001110110011;
ROM[3344] <= 32'b00000000011100000000001000110011;
ROM[3345] <= 32'b00000000001000000000000110110011;
ROM[3346] <= 32'b10110110110111111111000011101111;
ROM[3347] <= 32'b11111111110000010000000100010011;
ROM[3348] <= 32'b00000000000000010010001110000011;
ROM[3349] <= 32'b00000000011100011010000000100011;
ROM[3350] <= 32'b00000000000000011010001110000011;
ROM[3351] <= 32'b00000000011100010010000000100011;
ROM[3352] <= 32'b00000000010000010000000100010011;
ROM[3353] <= 32'b00000000010000000000001110010011;
ROM[3354] <= 32'b00000000011100010010000000100011;
ROM[3355] <= 32'b00000000010000010000000100010011;
ROM[3356] <= 32'b11111111110000010000000100010011;
ROM[3357] <= 32'b00000000000000010010001110000011;
ROM[3358] <= 32'b11111111110000010000000100010011;
ROM[3359] <= 32'b00000000000000010010010000000011;
ROM[3360] <= 32'b00000000011101000000001110110011;
ROM[3361] <= 32'b00000000011100010010000000100011;
ROM[3362] <= 32'b00000000010000010000000100010011;
ROM[3363] <= 32'b11111111110000010000000100010011;
ROM[3364] <= 32'b00000000000000010010001110000011;
ROM[3365] <= 32'b00000000011100011010010000100011;
ROM[3366] <= 32'b00000000100000011010001110000011;
ROM[3367] <= 32'b00000000011100010010000000100011;
ROM[3368] <= 32'b00000000010000010000000100010011;
ROM[3369] <= 32'b11111111110000010000000100010011;
ROM[3370] <= 32'b00000000000000010010001110000011;
ROM[3371] <= 32'b00000110011101101010010000100011;
ROM[3372] <= 32'b00000000000000011010001110000011;
ROM[3373] <= 32'b00000000011100010010000000100011;
ROM[3374] <= 32'b00000000010000010000000100010011;
ROM[3375] <= 32'b00000000000000000000001110010011;
ROM[3376] <= 32'b00000000011100010010000000100011;
ROM[3377] <= 32'b00000000010000010000000100010011;
ROM[3378] <= 32'b11111111110000010000000100010011;
ROM[3379] <= 32'b00000000000000010010001110000011;
ROM[3380] <= 32'b11111111110000010000000100010011;
ROM[3381] <= 32'b00000000000000010010010000000011;
ROM[3382] <= 32'b00000000011101000010010010110011;
ROM[3383] <= 32'b00000000100000111010010100110011;
ROM[3384] <= 32'b00000000101001001000001110110011;
ROM[3385] <= 32'b00000000000100111000001110010011;
ROM[3386] <= 32'b00000000000100111111001110010011;
ROM[3387] <= 32'b00000000011100010010000000100011;
ROM[3388] <= 32'b00000000010000010000000100010011;
ROM[3389] <= 32'b11111111110000010000000100010011;
ROM[3390] <= 32'b00000000000000010010001110000011;
ROM[3391] <= 32'b01000000011100000000001110110011;
ROM[3392] <= 32'b00000000000100111000001110010011;
ROM[3393] <= 32'b00000000011100010010000000100011;
ROM[3394] <= 32'b00000000010000010000000100010011;
ROM[3395] <= 32'b11111111110000010000000100010011;
ROM[3396] <= 32'b00000000000000010010001110000011;
ROM[3397] <= 32'b00000000000000111000101001100011;
ROM[3398] <= 32'b00000000000000000111001110110111;
ROM[3399] <= 32'b11011011000000111000001110010011;
ROM[3400] <= 32'b00000000111000111000001110110011;
ROM[3401] <= 32'b00000000000000111000000011100111;
ROM[3402] <= 32'b00001101010100000011000011101111;
ROM[3403] <= 32'b00000101110001101010001110000011;
ROM[3404] <= 32'b00000000011100010010000000100011;
ROM[3405] <= 32'b00000000010000010000000100010011;
ROM[3406] <= 32'b00000000000000011010001110000011;
ROM[3407] <= 32'b00000000011100010010000000100011;
ROM[3408] <= 32'b00000000010000010000000100010011;
ROM[3409] <= 32'b11111111110000010000000100010011;
ROM[3410] <= 32'b00000000000000010010001110000011;
ROM[3411] <= 32'b11111111110000010000000100010011;
ROM[3412] <= 32'b00000000000000010010010000000011;
ROM[3413] <= 32'b00000000011101000000001110110011;
ROM[3414] <= 32'b00000000011100010010000000100011;
ROM[3415] <= 32'b00000000010000010000000100010011;
ROM[3416] <= 32'b11111111110000010000000100010011;
ROM[3417] <= 32'b00000000000000010010001110000011;
ROM[3418] <= 32'b00000000000000111000001100010011;
ROM[3419] <= 32'b00000000110100110000010000110011;
ROM[3420] <= 32'b00000000000001000010001110000011;
ROM[3421] <= 32'b00000000011100010010000000100011;
ROM[3422] <= 32'b00000000010000010000000100010011;
ROM[3423] <= 32'b00000000000000100010001110000011;
ROM[3424] <= 32'b00000000011100010010000000100011;
ROM[3425] <= 32'b00000000010000010000000100010011;
ROM[3426] <= 32'b00000000001100000000001110010011;
ROM[3427] <= 32'b00000000011100010010000000100011;
ROM[3428] <= 32'b00000000010000010000000100010011;
ROM[3429] <= 32'b11111111110000010000000100010011;
ROM[3430] <= 32'b00000000000000010010001110000011;
ROM[3431] <= 32'b11111111110000010000000100010011;
ROM[3432] <= 32'b00000000000000010010010000000011;
ROM[3433] <= 32'b00000000011101000000001110110011;
ROM[3434] <= 32'b00000000011100010010000000100011;
ROM[3435] <= 32'b00000000010000010000000100010011;
ROM[3436] <= 32'b11111111110000010000000100010011;
ROM[3437] <= 32'b00000000000000010010001110000011;
ROM[3438] <= 32'b11111111110000010000000100010011;
ROM[3439] <= 32'b00000000000000010010010000000011;
ROM[3440] <= 32'b00000000100000111010001110110011;
ROM[3441] <= 32'b00000000011100010010000000100011;
ROM[3442] <= 32'b00000000010000010000000100010011;
ROM[3443] <= 32'b11111111110000010000000100010011;
ROM[3444] <= 32'b00000000000000010010001110000011;
ROM[3445] <= 32'b00000000000000111000101001100011;
ROM[3446] <= 32'b00000000000000000111001110110111;
ROM[3447] <= 32'b11111000100000111000001110010011;
ROM[3448] <= 32'b00000000111000111000001110110011;
ROM[3449] <= 32'b00000000000000111000000011100111;
ROM[3450] <= 32'b00011110110100000011000011101111;
ROM[3451] <= 32'b00000000000000011010001110000011;
ROM[3452] <= 32'b00000000011100010010000000100011;
ROM[3453] <= 32'b00000000010000010000000100010011;
ROM[3454] <= 32'b00000000000000100010001110000011;
ROM[3455] <= 32'b00000000011100010010000000100011;
ROM[3456] <= 32'b00000000010000010000000100010011;
ROM[3457] <= 32'b11111111110000010000000100010011;
ROM[3458] <= 32'b00000000000000010010001110000011;
ROM[3459] <= 32'b11111111110000010000000100010011;
ROM[3460] <= 32'b00000000000000010010010000000011;
ROM[3461] <= 32'b00000000011101000000001110110011;
ROM[3462] <= 32'b00000000011100010010000000100011;
ROM[3463] <= 32'b00000000010000010000000100010011;
ROM[3464] <= 32'b00000000000000100010001110000011;
ROM[3465] <= 32'b00000000011100010010000000100011;
ROM[3466] <= 32'b00000000010000010000000100010011;
ROM[3467] <= 32'b11111111110000010000000100010011;
ROM[3468] <= 32'b00000000000000010010001110000011;
ROM[3469] <= 32'b11111111110000010000000100010011;
ROM[3470] <= 32'b00000000000000010010010000000011;
ROM[3471] <= 32'b00000000011101000000001110110011;
ROM[3472] <= 32'b00000000011100010010000000100011;
ROM[3473] <= 32'b00000000010000010000000100010011;
ROM[3474] <= 32'b00000000000000100010001110000011;
ROM[3475] <= 32'b00000000011100010010000000100011;
ROM[3476] <= 32'b00000000010000010000000100010011;
ROM[3477] <= 32'b11111111110000010000000100010011;
ROM[3478] <= 32'b00000000000000010010001110000011;
ROM[3479] <= 32'b11111111110000010000000100010011;
ROM[3480] <= 32'b00000000000000010010010000000011;
ROM[3481] <= 32'b00000000011101000000001110110011;
ROM[3482] <= 32'b00000000011100010010000000100011;
ROM[3483] <= 32'b00000000010000010000000100010011;
ROM[3484] <= 32'b00000000000000100010001110000011;
ROM[3485] <= 32'b00000000011100010010000000100011;
ROM[3486] <= 32'b00000000010000010000000100010011;
ROM[3487] <= 32'b11111111110000010000000100010011;
ROM[3488] <= 32'b00000000000000010010001110000011;
ROM[3489] <= 32'b11111111110000010000000100010011;
ROM[3490] <= 32'b00000000000000010010010000000011;
ROM[3491] <= 32'b00000000011101000000001110110011;
ROM[3492] <= 32'b00000000011100010010000000100011;
ROM[3493] <= 32'b00000000010000010000000100010011;
ROM[3494] <= 32'b00000000010000000000001110010011;
ROM[3495] <= 32'b00000000011100010010000000100011;
ROM[3496] <= 32'b00000000010000010000000100010011;
ROM[3497] <= 32'b11111111110000010000000100010011;
ROM[3498] <= 32'b00000000000000010010001110000011;
ROM[3499] <= 32'b11111111110000010000000100010011;
ROM[3500] <= 32'b00000000000000010010010000000011;
ROM[3501] <= 32'b00000000011101000000001110110011;
ROM[3502] <= 32'b00000000011100010010000000100011;
ROM[3503] <= 32'b00000000010000010000000100010011;
ROM[3504] <= 32'b11111111110000010000000100010011;
ROM[3505] <= 32'b00000000000000010010001110000011;
ROM[3506] <= 32'b00000000011100011010001000100011;
ROM[3507] <= 32'b00000110000001101010001110000011;
ROM[3508] <= 32'b00000000011100010010000000100011;
ROM[3509] <= 32'b00000000010000010000000100010011;
ROM[3510] <= 32'b00000000010000011010001110000011;
ROM[3511] <= 32'b00000000011100010010000000100011;
ROM[3512] <= 32'b00000000010000010000000100010011;
ROM[3513] <= 32'b11111111110000010000000100010011;
ROM[3514] <= 32'b00000000000000010010001110000011;
ROM[3515] <= 32'b11111111110000010000000100010011;
ROM[3516] <= 32'b00000000000000010010010000000011;
ROM[3517] <= 32'b00000000011101000000001110110011;
ROM[3518] <= 32'b00000000011100010010000000100011;
ROM[3519] <= 32'b00000000010000010000000100010011;
ROM[3520] <= 32'b00000110000001101010001110000011;
ROM[3521] <= 32'b00000000011100010010000000100011;
ROM[3522] <= 32'b00000000010000010000000100010011;
ROM[3523] <= 32'b00000000000000011010001110000011;
ROM[3524] <= 32'b00000000011100010010000000100011;
ROM[3525] <= 32'b00000000010000010000000100010011;
ROM[3526] <= 32'b11111111110000010000000100010011;
ROM[3527] <= 32'b00000000000000010010001110000011;
ROM[3528] <= 32'b11111111110000010000000100010011;
ROM[3529] <= 32'b00000000000000010010010000000011;
ROM[3530] <= 32'b00000000011101000000001110110011;
ROM[3531] <= 32'b00000000011100010010000000100011;
ROM[3532] <= 32'b00000000010000010000000100010011;
ROM[3533] <= 32'b11111111110000010000000100010011;
ROM[3534] <= 32'b00000000000000010010001110000011;
ROM[3535] <= 32'b00000000000000111000001100010011;
ROM[3536] <= 32'b00000000110100110000010000110011;
ROM[3537] <= 32'b00000000000001000010001110000011;
ROM[3538] <= 32'b00000000011100010010000000100011;
ROM[3539] <= 32'b00000000010000010000000100010011;
ROM[3540] <= 32'b11111111110000010000000100010011;
ROM[3541] <= 32'b00000000000000010010001110000011;
ROM[3542] <= 32'b00000000011101100010000000100011;
ROM[3543] <= 32'b11111111110000010000000100010011;
ROM[3544] <= 32'b00000000000000010010001110000011;
ROM[3545] <= 32'b00000000000000111000001100010011;
ROM[3546] <= 32'b00000000000001100010001110000011;
ROM[3547] <= 32'b00000000011100010010000000100011;
ROM[3548] <= 32'b00000000010000010000000100010011;
ROM[3549] <= 32'b11111111110000010000000100010011;
ROM[3550] <= 32'b00000000000000010010001110000011;
ROM[3551] <= 32'b00000000110100110000010000110011;
ROM[3552] <= 32'b00000000011101000010000000100011;
ROM[3553] <= 32'b00000101110001101010001110000011;
ROM[3554] <= 32'b00000000011100010010000000100011;
ROM[3555] <= 32'b00000000010000010000000100010011;
ROM[3556] <= 32'b00000000010000011010001110000011;
ROM[3557] <= 32'b00000000011100010010000000100011;
ROM[3558] <= 32'b00000000010000010000000100010011;
ROM[3559] <= 32'b11111111110000010000000100010011;
ROM[3560] <= 32'b00000000000000010010001110000011;
ROM[3561] <= 32'b11111111110000010000000100010011;
ROM[3562] <= 32'b00000000000000010010010000000011;
ROM[3563] <= 32'b00000000011101000000001110110011;
ROM[3564] <= 32'b00000000011100010010000000100011;
ROM[3565] <= 32'b00000000010000010000000100010011;
ROM[3566] <= 32'b00000101110001101010001110000011;
ROM[3567] <= 32'b00000000011100010010000000100011;
ROM[3568] <= 32'b00000000010000010000000100010011;
ROM[3569] <= 32'b00000000000000011010001110000011;
ROM[3570] <= 32'b00000000011100010010000000100011;
ROM[3571] <= 32'b00000000010000010000000100010011;
ROM[3572] <= 32'b11111111110000010000000100010011;
ROM[3573] <= 32'b00000000000000010010001110000011;
ROM[3574] <= 32'b11111111110000010000000100010011;
ROM[3575] <= 32'b00000000000000010010010000000011;
ROM[3576] <= 32'b00000000011101000000001110110011;
ROM[3577] <= 32'b00000000011100010010000000100011;
ROM[3578] <= 32'b00000000010000010000000100010011;
ROM[3579] <= 32'b11111111110000010000000100010011;
ROM[3580] <= 32'b00000000000000010010001110000011;
ROM[3581] <= 32'b00000000000000111000001100010011;
ROM[3582] <= 32'b00000000110100110000010000110011;
ROM[3583] <= 32'b00000000000001000010001110000011;
ROM[3584] <= 32'b00000000011100010010000000100011;
ROM[3585] <= 32'b00000000010000010000000100010011;
ROM[3586] <= 32'b00000000000000100010001110000011;
ROM[3587] <= 32'b00000000011100010010000000100011;
ROM[3588] <= 32'b00000000010000010000000100010011;
ROM[3589] <= 32'b11111111110000010000000100010011;
ROM[3590] <= 32'b00000000000000010010001110000011;
ROM[3591] <= 32'b11111111110000010000000100010011;
ROM[3592] <= 32'b00000000000000010010010000000011;
ROM[3593] <= 32'b01000000011101000000001110110011;
ROM[3594] <= 32'b00000000011100010010000000100011;
ROM[3595] <= 32'b00000000010000010000000100010011;
ROM[3596] <= 32'b00000000000100000000001110010011;
ROM[3597] <= 32'b00000000011100010010000000100011;
ROM[3598] <= 32'b00000000010000010000000100010011;
ROM[3599] <= 32'b11111111110000010000000100010011;
ROM[3600] <= 32'b00000000000000010010001110000011;
ROM[3601] <= 32'b11111111110000010000000100010011;
ROM[3602] <= 32'b00000000000000010010010000000011;
ROM[3603] <= 32'b01000000011101000000001110110011;
ROM[3604] <= 32'b00000000011100010010000000100011;
ROM[3605] <= 32'b00000000010000010000000100010011;
ROM[3606] <= 32'b11111111110000010000000100010011;
ROM[3607] <= 32'b00000000000000010010001110000011;
ROM[3608] <= 32'b00000000011101100010000000100011;
ROM[3609] <= 32'b11111111110000010000000100010011;
ROM[3610] <= 32'b00000000000000010010001110000011;
ROM[3611] <= 32'b00000000000000111000001100010011;
ROM[3612] <= 32'b00000000000001100010001110000011;
ROM[3613] <= 32'b00000000011100010010000000100011;
ROM[3614] <= 32'b00000000010000010000000100010011;
ROM[3615] <= 32'b11111111110000010000000100010011;
ROM[3616] <= 32'b00000000000000010010001110000011;
ROM[3617] <= 32'b00000000110100110000010000110011;
ROM[3618] <= 32'b00000000011101000010000000100011;
ROM[3619] <= 32'b00000110010001101010001110000011;
ROM[3620] <= 32'b00000000011100010010000000100011;
ROM[3621] <= 32'b00000000010000010000000100010011;
ROM[3622] <= 32'b00000000100000011010001110000011;
ROM[3623] <= 32'b00000000011100010010000000100011;
ROM[3624] <= 32'b00000000010000010000000100010011;
ROM[3625] <= 32'b11111111110000010000000100010011;
ROM[3626] <= 32'b00000000000000010010001110000011;
ROM[3627] <= 32'b11111111110000010000000100010011;
ROM[3628] <= 32'b00000000000000010010010000000011;
ROM[3629] <= 32'b00000000011101000000001110110011;
ROM[3630] <= 32'b00000000011100010010000000100011;
ROM[3631] <= 32'b00000000010000010000000100010011;
ROM[3632] <= 32'b00000000000000100010001110000011;
ROM[3633] <= 32'b00000000011100010010000000100011;
ROM[3634] <= 32'b00000000010000010000000100010011;
ROM[3635] <= 32'b00000000000100000000001110010011;
ROM[3636] <= 32'b00000000011100010010000000100011;
ROM[3637] <= 32'b00000000010000010000000100010011;
ROM[3638] <= 32'b11111111110000010000000100010011;
ROM[3639] <= 32'b00000000000000010010001110000011;
ROM[3640] <= 32'b11111111110000010000000100010011;
ROM[3641] <= 32'b00000000000000010010010000000011;
ROM[3642] <= 32'b00000000011101000000001110110011;
ROM[3643] <= 32'b00000000011100010010000000100011;
ROM[3644] <= 32'b00000000010000010000000100010011;
ROM[3645] <= 32'b11111111110000010000000100010011;
ROM[3646] <= 32'b00000000000000010010001110000011;
ROM[3647] <= 32'b00000000011101100010000000100011;
ROM[3648] <= 32'b11111111110000010000000100010011;
ROM[3649] <= 32'b00000000000000010010001110000011;
ROM[3650] <= 32'b00000000000000111000001100010011;
ROM[3651] <= 32'b00000000000001100010001110000011;
ROM[3652] <= 32'b00000000011100010010000000100011;
ROM[3653] <= 32'b00000000010000010000000100010011;
ROM[3654] <= 32'b11111111110000010000000100010011;
ROM[3655] <= 32'b00000000000000010010001110000011;
ROM[3656] <= 32'b00000000110100110000010000110011;
ROM[3657] <= 32'b00000000011101000010000000100011;
ROM[3658] <= 32'b00000000100000011010001110000011;
ROM[3659] <= 32'b00000000011100010010000000100011;
ROM[3660] <= 32'b00000000010000010000000100010011;
ROM[3661] <= 32'b11111111110000010000000100010011;
ROM[3662] <= 32'b00000000000000010010001110000011;
ROM[3663] <= 32'b00000110011101101010011000100011;
ROM[3664] <= 32'b00000000010000011010001110000011;
ROM[3665] <= 32'b00000000011100010010000000100011;
ROM[3666] <= 32'b00000000010000010000000100010011;
ROM[3667] <= 32'b11111111110000010000000100010011;
ROM[3668] <= 32'b00000000000000010010001110000011;
ROM[3669] <= 32'b00000100011101101010110000100011;
ROM[3670] <= 32'b00000000000100000000001110010011;
ROM[3671] <= 32'b00000000011100010010000000100011;
ROM[3672] <= 32'b00000000010000010000000100010011;
ROM[3673] <= 32'b11111111110000010000000100010011;
ROM[3674] <= 32'b00000000000000010010001110000011;
ROM[3675] <= 32'b00000110011101101010100000100011;
ROM[3676] <= 32'b01101001010000000011000011101111;
ROM[3677] <= 32'b00000110000001101010001110000011;
ROM[3678] <= 32'b00000000011100010010000000100011;
ROM[3679] <= 32'b00000000010000010000000100010011;
ROM[3680] <= 32'b00000000000000011010001110000011;
ROM[3681] <= 32'b00000000011100010010000000100011;
ROM[3682] <= 32'b00000000010000010000000100010011;
ROM[3683] <= 32'b11111111110000010000000100010011;
ROM[3684] <= 32'b00000000000000010010001110000011;
ROM[3685] <= 32'b11111111110000010000000100010011;
ROM[3686] <= 32'b00000000000000010010010000000011;
ROM[3687] <= 32'b00000000011101000000001110110011;
ROM[3688] <= 32'b00000000011100010010000000100011;
ROM[3689] <= 32'b00000000010000010000000100010011;
ROM[3690] <= 32'b11111111110000010000000100010011;
ROM[3691] <= 32'b00000000000000010010001110000011;
ROM[3692] <= 32'b00000000000000111000001100010011;
ROM[3693] <= 32'b00000000110100110000010000110011;
ROM[3694] <= 32'b00000000000001000010001110000011;
ROM[3695] <= 32'b00000000011100010010000000100011;
ROM[3696] <= 32'b00000000010000010000000100010011;
ROM[3697] <= 32'b11111111110000010000000100010011;
ROM[3698] <= 32'b00000000000000010010001110000011;
ROM[3699] <= 32'b00000000011100011010001000100011;
ROM[3700] <= 32'b00000110010001101010001110000011;
ROM[3701] <= 32'b00000000011100010010000000100011;
ROM[3702] <= 32'b00000000010000010000000100010011;
ROM[3703] <= 32'b00000000100000011010001110000011;
ROM[3704] <= 32'b00000000011100010010000000100011;
ROM[3705] <= 32'b00000000010000010000000100010011;
ROM[3706] <= 32'b11111111110000010000000100010011;
ROM[3707] <= 32'b00000000000000010010001110000011;
ROM[3708] <= 32'b11111111110000010000000100010011;
ROM[3709] <= 32'b00000000000000010010010000000011;
ROM[3710] <= 32'b00000000011101000000001110110011;
ROM[3711] <= 32'b00000000011100010010000000100011;
ROM[3712] <= 32'b00000000010000010000000100010011;
ROM[3713] <= 32'b00000101110001101010001110000011;
ROM[3714] <= 32'b00000000011100010010000000100011;
ROM[3715] <= 32'b00000000010000010000000100010011;
ROM[3716] <= 32'b00000000000000011010001110000011;
ROM[3717] <= 32'b00000000011100010010000000100011;
ROM[3718] <= 32'b00000000010000010000000100010011;
ROM[3719] <= 32'b11111111110000010000000100010011;
ROM[3720] <= 32'b00000000000000010010001110000011;
ROM[3721] <= 32'b11111111110000010000000100010011;
ROM[3722] <= 32'b00000000000000010010010000000011;
ROM[3723] <= 32'b00000000011101000000001110110011;
ROM[3724] <= 32'b00000000011100010010000000100011;
ROM[3725] <= 32'b00000000010000010000000100010011;
ROM[3726] <= 32'b11111111110000010000000100010011;
ROM[3727] <= 32'b00000000000000010010001110000011;
ROM[3728] <= 32'b00000000000000111000001100010011;
ROM[3729] <= 32'b00000000110100110000010000110011;
ROM[3730] <= 32'b00000000000001000010001110000011;
ROM[3731] <= 32'b00000000011100010010000000100011;
ROM[3732] <= 32'b00000000010000010000000100010011;
ROM[3733] <= 32'b11111111110000010000000100010011;
ROM[3734] <= 32'b00000000000000010010001110000011;
ROM[3735] <= 32'b00000000011101100010000000100011;
ROM[3736] <= 32'b11111111110000010000000100010011;
ROM[3737] <= 32'b00000000000000010010001110000011;
ROM[3738] <= 32'b00000000000000111000001100010011;
ROM[3739] <= 32'b00000000000001100010001110000011;
ROM[3740] <= 32'b00000000011100010010000000100011;
ROM[3741] <= 32'b00000000010000010000000100010011;
ROM[3742] <= 32'b11111111110000010000000100010011;
ROM[3743] <= 32'b00000000000000010010001110000011;
ROM[3744] <= 32'b00000000110100110000010000110011;
ROM[3745] <= 32'b00000000011101000010000000100011;
ROM[3746] <= 32'b00000000001000000000001110010011;
ROM[3747] <= 32'b00000000011100010010000000100011;
ROM[3748] <= 32'b00000000010000010000000100010011;
ROM[3749] <= 32'b11111111110000010000000100010011;
ROM[3750] <= 32'b00000000000000010010001110000011;
ROM[3751] <= 32'b00000110011101101010100000100011;
ROM[3752] <= 32'b00110101110000000011000011101111;
ROM[3753] <= 32'b00000000100000011010001110000011;
ROM[3754] <= 32'b00000000011100010010000000100011;
ROM[3755] <= 32'b00000000010000010000000100010011;
ROM[3756] <= 32'b00000001010000000000001110010011;
ROM[3757] <= 32'b01000000011100011000001110110011;
ROM[3758] <= 32'b00000000000000111010000010000011;
ROM[3759] <= 32'b11111111110000010000000100010011;
ROM[3760] <= 32'b00000000000000010010001110000011;
ROM[3761] <= 32'b00000000011100100010000000100011;
ROM[3762] <= 32'b00000000010000100000000100010011;
ROM[3763] <= 32'b00000001010000000000001110010011;
ROM[3764] <= 32'b01000000011100011000001110110011;
ROM[3765] <= 32'b00000000010000111010000110000011;
ROM[3766] <= 32'b00000000100000111010001000000011;
ROM[3767] <= 32'b00000000110000111010001010000011;
ROM[3768] <= 32'b00000001000000111010001100000011;
ROM[3769] <= 32'b00000000000000001000000011100111;
ROM[3770] <= 32'b00000000000000000100001110110111;
ROM[3771] <= 32'b00000000000000111000001110010011;
ROM[3772] <= 32'b00000000011100010010000000100011;
ROM[3773] <= 32'b00000000010000010000000100010011;
ROM[3774] <= 32'b11111111110000010000000100010011;
ROM[3775] <= 32'b00000000000000010010001110000011;
ROM[3776] <= 32'b00000110011101101010101000100011;
ROM[3777] <= 32'b00000000000000000000001110010011;
ROM[3778] <= 32'b00000000011100010010000000100011;
ROM[3779] <= 32'b00000000010000010000000100010011;
ROM[3780] <= 32'b11111111110000010000000100010011;
ROM[3781] <= 32'b00000000000000010010001110000011;
ROM[3782] <= 32'b00000110011101101010110000100011;
ROM[3783] <= 32'b00000000000000000000001110010011;
ROM[3784] <= 32'b00000000011100010010000000100011;
ROM[3785] <= 32'b00000000010000010000000100010011;
ROM[3786] <= 32'b11111111110000010000000100010011;
ROM[3787] <= 32'b00000000000000010010001110000011;
ROM[3788] <= 32'b00000110011101101010111000100011;
ROM[3789] <= 32'b00000000000000000000001110010011;
ROM[3790] <= 32'b00000000011100010010000000100011;
ROM[3791] <= 32'b00000000010000010000000100010011;
ROM[3792] <= 32'b11111111110000010000000100010011;
ROM[3793] <= 32'b00000000000000010010001110000011;
ROM[3794] <= 32'b00001000011101101010000000100011;
ROM[3795] <= 32'b00000000000000000000001110010011;
ROM[3796] <= 32'b00000000011100010010000000100011;
ROM[3797] <= 32'b00000000010000010000000100010011;
ROM[3798] <= 32'b11111111110000010000000100010011;
ROM[3799] <= 32'b00000000000000010010001110000011;
ROM[3800] <= 32'b00001000011101101010001000100011;
ROM[3801] <= 32'b00000000000000000000001110010011;
ROM[3802] <= 32'b00000000011100010010000000100011;
ROM[3803] <= 32'b00000000010000010000000100010011;
ROM[3804] <= 32'b11111111110000010000000100010011;
ROM[3805] <= 32'b00000000000000010010001110000011;
ROM[3806] <= 32'b00001000011101101010010000100011;
ROM[3807] <= 32'b00000010010000000000001110010011;
ROM[3808] <= 32'b00000000011100010010000000100011;
ROM[3809] <= 32'b00000000010000010000000100010011;
ROM[3810] <= 32'b00000000000000000100001110110111;
ROM[3811] <= 32'b10111101010000111000001110010011;
ROM[3812] <= 32'b00000000111000111000001110110011;
ROM[3813] <= 32'b00000000011100010010000000100011;
ROM[3814] <= 32'b00000000010000010000000100010011;
ROM[3815] <= 32'b00000000001100010010000000100011;
ROM[3816] <= 32'b00000000010000010000000100010011;
ROM[3817] <= 32'b00000000010000010010000000100011;
ROM[3818] <= 32'b00000000010000010000000100010011;
ROM[3819] <= 32'b00000000010100010010000000100011;
ROM[3820] <= 32'b00000000010000010000000100010011;
ROM[3821] <= 32'b00000000011000010010000000100011;
ROM[3822] <= 32'b00000000010000010000000100010011;
ROM[3823] <= 32'b00000001010000000000001110010011;
ROM[3824] <= 32'b00000000010000111000001110010011;
ROM[3825] <= 32'b01000000011100010000001110110011;
ROM[3826] <= 32'b00000000011100000000001000110011;
ROM[3827] <= 32'b00000000001000000000000110110011;
ROM[3828] <= 32'b10000111000111111100000011101111;
ROM[3829] <= 32'b11111111110000010000000100010011;
ROM[3830] <= 32'b00000000000000010010001110000011;
ROM[3831] <= 32'b00001000011101101010011000100011;
ROM[3832] <= 32'b00000000000000000100001110110111;
ROM[3833] <= 32'b11000010110000111000001110010011;
ROM[3834] <= 32'b00000000111000111000001110110011;
ROM[3835] <= 32'b00000000011100010010000000100011;
ROM[3836] <= 32'b00000000010000010000000100010011;
ROM[3837] <= 32'b00000000001100010010000000100011;
ROM[3838] <= 32'b00000000010000010000000100010011;
ROM[3839] <= 32'b00000000010000010010000000100011;
ROM[3840] <= 32'b00000000010000010000000100010011;
ROM[3841] <= 32'b00000000010100010010000000100011;
ROM[3842] <= 32'b00000000010000010000000100010011;
ROM[3843] <= 32'b00000000011000010010000000100011;
ROM[3844] <= 32'b00000000010000010000000100010011;
ROM[3845] <= 32'b00000001010000000000001110010011;
ROM[3846] <= 32'b00000000000000111000001110010011;
ROM[3847] <= 32'b01000000011100010000001110110011;
ROM[3848] <= 32'b00000000011100000000001000110011;
ROM[3849] <= 32'b00000000001000000000000110110011;
ROM[3850] <= 32'b00001010110000000000000011101111;
ROM[3851] <= 32'b11111111110000010000000100010011;
ROM[3852] <= 32'b00000000000000010010001110000011;
ROM[3853] <= 32'b00000000011101100010000000100011;
ROM[3854] <= 32'b00000000000000000100001110110111;
ROM[3855] <= 32'b11001000010000111000001110010011;
ROM[3856] <= 32'b00000000111000111000001110110011;
ROM[3857] <= 32'b00000000011100010010000000100011;
ROM[3858] <= 32'b00000000010000010000000100010011;
ROM[3859] <= 32'b00000000001100010010000000100011;
ROM[3860] <= 32'b00000000010000010000000100010011;
ROM[3861] <= 32'b00000000010000010010000000100011;
ROM[3862] <= 32'b00000000010000010000000100010011;
ROM[3863] <= 32'b00000000010100010010000000100011;
ROM[3864] <= 32'b00000000010000010000000100010011;
ROM[3865] <= 32'b00000000011000010010000000100011;
ROM[3866] <= 32'b00000000010000010000000100010011;
ROM[3867] <= 32'b00000001010000000000001110010011;
ROM[3868] <= 32'b00000000000000111000001110010011;
ROM[3869] <= 32'b01000000011100010000001110110011;
ROM[3870] <= 32'b00000000011100000000001000110011;
ROM[3871] <= 32'b00000000001000000000000110110011;
ROM[3872] <= 32'b00101111010100000000000011101111;
ROM[3873] <= 32'b11111111110000010000000100010011;
ROM[3874] <= 32'b00000000000000010010001110000011;
ROM[3875] <= 32'b00000000011101100010000000100011;
ROM[3876] <= 32'b00000000000000000000001110010011;
ROM[3877] <= 32'b00000000011100010010000000100011;
ROM[3878] <= 32'b00000000010000010000000100010011;
ROM[3879] <= 32'b00000001010000000000001110010011;
ROM[3880] <= 32'b01000000011100011000001110110011;
ROM[3881] <= 32'b00000000000000111010000010000011;
ROM[3882] <= 32'b11111111110000010000000100010011;
ROM[3883] <= 32'b00000000000000010010001110000011;
ROM[3884] <= 32'b00000000011100100010000000100011;
ROM[3885] <= 32'b00000000010000100000000100010011;
ROM[3886] <= 32'b00000001010000000000001110010011;
ROM[3887] <= 32'b01000000011100011000001110110011;
ROM[3888] <= 32'b00000000010000111010000110000011;
ROM[3889] <= 32'b00000000100000111010001000000011;
ROM[3890] <= 32'b00000000110000111010001010000011;
ROM[3891] <= 32'b00000001000000111010001100000011;
ROM[3892] <= 32'b00000000000000001000000011100111;
ROM[3893] <= 32'b00000000000000010010000000100011;
ROM[3894] <= 32'b00000000010000010000000100010011;
ROM[3895] <= 32'b00000111111100000000001110010011;
ROM[3896] <= 32'b00000000011100010010000000100011;
ROM[3897] <= 32'b00000000010000010000000100010011;
ROM[3898] <= 32'b00000000000000000100001110110111;
ROM[3899] <= 32'b11010011010000111000001110010011;
ROM[3900] <= 32'b00000000111000111000001110110011;
ROM[3901] <= 32'b00000000011100010010000000100011;
ROM[3902] <= 32'b00000000010000010000000100010011;
ROM[3903] <= 32'b00000000001100010010000000100011;
ROM[3904] <= 32'b00000000010000010000000100010011;
ROM[3905] <= 32'b00000000010000010010000000100011;
ROM[3906] <= 32'b00000000010000010000000100010011;
ROM[3907] <= 32'b00000000010100010010000000100011;
ROM[3908] <= 32'b00000000010000010000000100010011;
ROM[3909] <= 32'b00000000011000010010000000100011;
ROM[3910] <= 32'b00000000010000010000000100010011;
ROM[3911] <= 32'b00000001010000000000001110010011;
ROM[3912] <= 32'b00000000010000111000001110010011;
ROM[3913] <= 32'b01000000011100010000001110110011;
ROM[3914] <= 32'b00000000011100000000001000110011;
ROM[3915] <= 32'b00000000001000000000000110110011;
ROM[3916] <= 32'b11110001000011111100000011101111;
ROM[3917] <= 32'b11111111110000010000000100010011;
ROM[3918] <= 32'b00000000000000010010001110000011;
ROM[3919] <= 32'b00001000011101101010100000100011;
ROM[3920] <= 32'b00000011000000000000001110010011;
ROM[3921] <= 32'b00000000011100010010000000100011;
ROM[3922] <= 32'b00000000010000010000000100010011;
ROM[3923] <= 32'b00000011111000000000001110010011;
ROM[3924] <= 32'b00000000011100010010000000100011;
ROM[3925] <= 32'b00000000010000010000000100010011;
ROM[3926] <= 32'b00000100001100000000001110010011;
ROM[3927] <= 32'b00000000011100010010000000100011;
ROM[3928] <= 32'b00000000010000010000000100010011;
ROM[3929] <= 32'b00000100010100000000001110010011;
ROM[3930] <= 32'b00000000011100010010000000100011;
ROM[3931] <= 32'b00000000010000010000000100010011;
ROM[3932] <= 32'b00000100100100000000001110010011;
ROM[3933] <= 32'b00000000011100010010000000100011;
ROM[3934] <= 32'b00000000010000010000000100010011;
ROM[3935] <= 32'b00000101000100000000001110010011;
ROM[3936] <= 32'b00000000011100010010000000100011;
ROM[3937] <= 32'b00000000010000010000000100010011;
ROM[3938] <= 32'b00000110000100000000001110010011;
ROM[3939] <= 32'b00000000011100010010000000100011;
ROM[3940] <= 32'b00000000010000010000000100010011;
ROM[3941] <= 32'b00000011111000000000001110010011;
ROM[3942] <= 32'b00000000011100010010000000100011;
ROM[3943] <= 32'b00000000010000010000000100010011;
ROM[3944] <= 32'b00000000000000000100001110110111;
ROM[3945] <= 32'b11011110110000111000001110010011;
ROM[3946] <= 32'b00000000111000111000001110110011;
ROM[3947] <= 32'b00000000011100010010000000100011;
ROM[3948] <= 32'b00000000010000010000000100010011;
ROM[3949] <= 32'b00000000001100010010000000100011;
ROM[3950] <= 32'b00000000010000010000000100010011;
ROM[3951] <= 32'b00000000010000010010000000100011;
ROM[3952] <= 32'b00000000010000010000000100010011;
ROM[3953] <= 32'b00000000010100010010000000100011;
ROM[3954] <= 32'b00000000010000010000000100010011;
ROM[3955] <= 32'b00000000011000010010000000100011;
ROM[3956] <= 32'b00000000010000010000000100010011;
ROM[3957] <= 32'b00000001010000000000001110010011;
ROM[3958] <= 32'b00000010000000111000001110010011;
ROM[3959] <= 32'b01000000011100010000001110110011;
ROM[3960] <= 32'b00000000011100000000001000110011;
ROM[3961] <= 32'b00000000001000000000000110110011;
ROM[3962] <= 32'b01001010010000000000000011101111;
ROM[3963] <= 32'b11111111110000010000000100010011;
ROM[3964] <= 32'b00000000000000010010001110000011;
ROM[3965] <= 32'b00000000011101100010000000100011;
ROM[3966] <= 32'b00000011000100000000001110010011;
ROM[3967] <= 32'b00000000011100010010000000100011;
ROM[3968] <= 32'b00000000010000010000000100010011;
ROM[3969] <= 32'b00000000100000000000001110010011;
ROM[3970] <= 32'b00000000011100010010000000100011;
ROM[3971] <= 32'b00000000010000010000000100010011;
ROM[3972] <= 32'b00000001100000000000001110010011;
ROM[3973] <= 32'b00000000011100010010000000100011;
ROM[3974] <= 32'b00000000010000010000000100010011;
ROM[3975] <= 32'b00000010100000000000001110010011;
ROM[3976] <= 32'b00000000011100010010000000100011;
ROM[3977] <= 32'b00000000010000010000000100010011;
ROM[3978] <= 32'b00000000100000000000001110010011;
ROM[3979] <= 32'b00000000011100010010000000100011;
ROM[3980] <= 32'b00000000010000010000000100010011;
ROM[3981] <= 32'b00000000100000000000001110010011;
ROM[3982] <= 32'b00000000011100010010000000100011;
ROM[3983] <= 32'b00000000010000010000000100010011;
ROM[3984] <= 32'b00000000100000000000001110010011;
ROM[3985] <= 32'b00000000011100010010000000100011;
ROM[3986] <= 32'b00000000010000010000000100010011;
ROM[3987] <= 32'b00000111111100000000001110010011;
ROM[3988] <= 32'b00000000011100010010000000100011;
ROM[3989] <= 32'b00000000010000010000000100010011;
ROM[3990] <= 32'b00000000000000000100001110110111;
ROM[3991] <= 32'b11101010010000111000001110010011;
ROM[3992] <= 32'b00000000111000111000001110110011;
ROM[3993] <= 32'b00000000011100010010000000100011;
ROM[3994] <= 32'b00000000010000010000000100010011;
ROM[3995] <= 32'b00000000001100010010000000100011;
ROM[3996] <= 32'b00000000010000010000000100010011;
ROM[3997] <= 32'b00000000010000010010000000100011;
ROM[3998] <= 32'b00000000010000010000000100010011;
ROM[3999] <= 32'b00000000010100010010000000100011;
ROM[4000] <= 32'b00000000010000010000000100010011;
ROM[4001] <= 32'b00000000011000010010000000100011;
ROM[4002] <= 32'b00000000010000010000000100010011;
ROM[4003] <= 32'b00000001010000000000001110010011;
ROM[4004] <= 32'b00000010000000111000001110010011;
ROM[4005] <= 32'b01000000011100010000001110110011;
ROM[4006] <= 32'b00000000011100000000001000110011;
ROM[4007] <= 32'b00000000001000000000000110110011;
ROM[4008] <= 32'b00111110110000000000000011101111;
ROM[4009] <= 32'b11111111110000010000000100010011;
ROM[4010] <= 32'b00000000000000010010001110000011;
ROM[4011] <= 32'b00000000011101100010000000100011;
ROM[4012] <= 32'b00000011001000000000001110010011;
ROM[4013] <= 32'b00000000011100010010000000100011;
ROM[4014] <= 32'b00000000010000010000000100010011;
ROM[4015] <= 32'b00000111111100000000001110010011;
ROM[4016] <= 32'b00000000011100010010000000100011;
ROM[4017] <= 32'b00000000010000010000000100010011;
ROM[4018] <= 32'b00000000000100000000001110010011;
ROM[4019] <= 32'b00000000011100010010000000100011;
ROM[4020] <= 32'b00000000010000010000000100010011;
ROM[4021] <= 32'b00000000000100000000001110010011;
ROM[4022] <= 32'b00000000011100010010000000100011;
ROM[4023] <= 32'b00000000010000010000000100010011;
ROM[4024] <= 32'b00000111111100000000001110010011;
ROM[4025] <= 32'b00000000011100010010000000100011;
ROM[4026] <= 32'b00000000010000010000000100010011;
ROM[4027] <= 32'b00000100000000000000001110010011;
ROM[4028] <= 32'b00000000011100010010000000100011;
ROM[4029] <= 32'b00000000010000010000000100010011;
ROM[4030] <= 32'b00000100000000000000001110010011;
ROM[4031] <= 32'b00000000011100010010000000100011;
ROM[4032] <= 32'b00000000010000010000000100010011;
ROM[4033] <= 32'b00000111111100000000001110010011;
ROM[4034] <= 32'b00000000011100010010000000100011;
ROM[4035] <= 32'b00000000010000010000000100010011;
ROM[4036] <= 32'b00000000000000000100001110110111;
ROM[4037] <= 32'b11110101110000111000001110010011;
ROM[4038] <= 32'b00000000111000111000001110110011;
ROM[4039] <= 32'b00000000011100010010000000100011;
ROM[4040] <= 32'b00000000010000010000000100010011;
ROM[4041] <= 32'b00000000001100010010000000100011;
ROM[4042] <= 32'b00000000010000010000000100010011;
ROM[4043] <= 32'b00000000010000010010000000100011;
ROM[4044] <= 32'b00000000010000010000000100010011;
ROM[4045] <= 32'b00000000010100010010000000100011;
ROM[4046] <= 32'b00000000010000010000000100010011;
ROM[4047] <= 32'b00000000011000010010000000100011;
ROM[4048] <= 32'b00000000010000010000000100010011;
ROM[4049] <= 32'b00000001010000000000001110010011;
ROM[4050] <= 32'b00000010000000111000001110010011;
ROM[4051] <= 32'b01000000011100010000001110110011;
ROM[4052] <= 32'b00000000011100000000001000110011;
ROM[4053] <= 32'b00000000001000000000000110110011;
ROM[4054] <= 32'b00110011010000000000000011101111;
ROM[4055] <= 32'b11111111110000010000000100010011;
ROM[4056] <= 32'b00000000000000010010001110000011;
ROM[4057] <= 32'b00000000011101100010000000100011;
ROM[4058] <= 32'b00000100000100000000001110010011;
ROM[4059] <= 32'b00000000011100010010000000100011;
ROM[4060] <= 32'b00000000010000010000000100010011;
ROM[4061] <= 32'b00000111111100000000001110010011;
ROM[4062] <= 32'b00000000011100010010000000100011;
ROM[4063] <= 32'b00000000010000010000000100010011;
ROM[4064] <= 32'b00000100000100000000001110010011;
ROM[4065] <= 32'b00000000011100010010000000100011;
ROM[4066] <= 32'b00000000010000010000000100010011;
ROM[4067] <= 32'b00000100000100000000001110010011;
ROM[4068] <= 32'b00000000011100010010000000100011;
ROM[4069] <= 32'b00000000010000010000000100010011;
ROM[4070] <= 32'b00000100000100000000001110010011;
ROM[4071] <= 32'b00000000011100010010000000100011;
ROM[4072] <= 32'b00000000010000010000000100010011;
ROM[4073] <= 32'b00000111111100000000001110010011;
ROM[4074] <= 32'b00000000011100010010000000100011;
ROM[4075] <= 32'b00000000010000010000000100010011;
ROM[4076] <= 32'b00000100000100000000001110010011;
ROM[4077] <= 32'b00000000011100010010000000100011;
ROM[4078] <= 32'b00000000010000010000000100010011;
ROM[4079] <= 32'b00000100000100000000001110010011;
ROM[4080] <= 32'b00000000011100010010000000100011;
ROM[4081] <= 32'b00000000010000010000000100010011;
ROM[4082] <= 32'b00000000000000000100001110110111;
ROM[4083] <= 32'b00000001010000111000001110010011;
ROM[4084] <= 32'b00000000111000111000001110110011;
ROM[4085] <= 32'b00000000011100010010000000100011;
ROM[4086] <= 32'b00000000010000010000000100010011;
ROM[4087] <= 32'b00000000001100010010000000100011;
ROM[4088] <= 32'b00000000010000010000000100010011;
ROM[4089] <= 32'b00000000010000010010000000100011;
ROM[4090] <= 32'b00000000010000010000000100010011;
ROM[4091] <= 32'b00000000010100010010000000100011;
ROM[4092] <= 32'b00000000010000010000000100010011;
ROM[4093] <= 32'b00000000011000010010000000100011;
ROM[4094] <= 32'b00000000010000010000000100010011;
ROM[4095] <= 32'b00000001010000000000001110010011;
ROM[4096] <= 32'b00000010000000111000001110010011;
ROM[4097] <= 32'b01000000011100010000001110110011;
ROM[4098] <= 32'b00000000011100000000001000110011;
ROM[4099] <= 32'b00000000001000000000000110110011;
ROM[4100] <= 32'b00100111110000000000000011101111;
ROM[4101] <= 32'b11111111110000010000000100010011;
ROM[4102] <= 32'b00000000000000010010001110000011;
ROM[4103] <= 32'b00000000011101100010000000100011;
ROM[4104] <= 32'b00000100001000000000001110010011;
ROM[4105] <= 32'b00000000011100010010000000100011;
ROM[4106] <= 32'b00000000010000010000000100010011;
ROM[4107] <= 32'b00000111111000000000001110010011;
ROM[4108] <= 32'b00000000011100010010000000100011;
ROM[4109] <= 32'b00000000010000010000000100010011;
ROM[4110] <= 32'b00000100000100000000001110010011;
ROM[4111] <= 32'b00000000011100010010000000100011;
ROM[4112] <= 32'b00000000010000010000000100010011;
ROM[4113] <= 32'b00000100000100000000001110010011;
ROM[4114] <= 32'b00000000011100010010000000100011;
ROM[4115] <= 32'b00000000010000010000000100010011;
ROM[4116] <= 32'b00000111111000000000001110010011;
ROM[4117] <= 32'b00000000011100010010000000100011;
ROM[4118] <= 32'b00000000010000010000000100010011;
ROM[4119] <= 32'b00000100000100000000001110010011;
ROM[4120] <= 32'b00000000011100010010000000100011;
ROM[4121] <= 32'b00000000010000010000000100010011;
ROM[4122] <= 32'b00000100000100000000001110010011;
ROM[4123] <= 32'b00000000011100010010000000100011;
ROM[4124] <= 32'b00000000010000010000000100010011;
ROM[4125] <= 32'b00000111111000000000001110010011;
ROM[4126] <= 32'b00000000011100010010000000100011;
ROM[4127] <= 32'b00000000010000010000000100010011;
ROM[4128] <= 32'b00000000000000000100001110110111;
ROM[4129] <= 32'b00001100110000111000001110010011;
ROM[4130] <= 32'b00000000111000111000001110110011;
ROM[4131] <= 32'b00000000011100010010000000100011;
ROM[4132] <= 32'b00000000010000010000000100010011;
ROM[4133] <= 32'b00000000001100010010000000100011;
ROM[4134] <= 32'b00000000010000010000000100010011;
ROM[4135] <= 32'b00000000010000010010000000100011;
ROM[4136] <= 32'b00000000010000010000000100010011;
ROM[4137] <= 32'b00000000010100010010000000100011;
ROM[4138] <= 32'b00000000010000010000000100010011;
ROM[4139] <= 32'b00000000011000010010000000100011;
ROM[4140] <= 32'b00000000010000010000000100010011;
ROM[4141] <= 32'b00000001010000000000001110010011;
ROM[4142] <= 32'b00000010000000111000001110010011;
ROM[4143] <= 32'b01000000011100010000001110110011;
ROM[4144] <= 32'b00000000011100000000001000110011;
ROM[4145] <= 32'b00000000001000000000000110110011;
ROM[4146] <= 32'b00011100010000000000000011101111;
ROM[4147] <= 32'b11111111110000010000000100010011;
ROM[4148] <= 32'b00000000000000010010001110000011;
ROM[4149] <= 32'b00000000011101100010000000100011;
ROM[4150] <= 32'b00000100001100000000001110010011;
ROM[4151] <= 32'b00000000011100010010000000100011;
ROM[4152] <= 32'b00000000010000010000000100010011;
ROM[4153] <= 32'b00000111111100000000001110010011;
ROM[4154] <= 32'b00000000011100010010000000100011;
ROM[4155] <= 32'b00000000010000010000000100010011;
ROM[4156] <= 32'b00000100000100000000001110010011;
ROM[4157] <= 32'b00000000011100010010000000100011;
ROM[4158] <= 32'b00000000010000010000000100010011;
ROM[4159] <= 32'b00000100000100000000001110010011;
ROM[4160] <= 32'b00000000011100010010000000100011;
ROM[4161] <= 32'b00000000010000010000000100010011;
ROM[4162] <= 32'b00000100000100000000001110010011;
ROM[4163] <= 32'b00000000011100010010000000100011;
ROM[4164] <= 32'b00000000010000010000000100010011;
ROM[4165] <= 32'b00000100000100000000001110010011;
ROM[4166] <= 32'b00000000011100010010000000100011;
ROM[4167] <= 32'b00000000010000010000000100010011;
ROM[4168] <= 32'b00000100000100000000001110010011;
ROM[4169] <= 32'b00000000011100010010000000100011;
ROM[4170] <= 32'b00000000010000010000000100010011;
ROM[4171] <= 32'b00000111111100000000001110010011;
ROM[4172] <= 32'b00000000011100010010000000100011;
ROM[4173] <= 32'b00000000010000010000000100010011;
ROM[4174] <= 32'b00000000000000000100001110110111;
ROM[4175] <= 32'b00011000010000111000001110010011;
ROM[4176] <= 32'b00000000111000111000001110110011;
ROM[4177] <= 32'b00000000011100010010000000100011;
ROM[4178] <= 32'b00000000010000010000000100010011;
ROM[4179] <= 32'b00000000001100010010000000100011;
ROM[4180] <= 32'b00000000010000010000000100010011;
ROM[4181] <= 32'b00000000010000010010000000100011;
ROM[4182] <= 32'b00000000010000010000000100010011;
ROM[4183] <= 32'b00000000010100010010000000100011;
ROM[4184] <= 32'b00000000010000010000000100010011;
ROM[4185] <= 32'b00000000011000010010000000100011;
ROM[4186] <= 32'b00000000010000010000000100010011;
ROM[4187] <= 32'b00000001010000000000001110010011;
ROM[4188] <= 32'b00000010000000111000001110010011;
ROM[4189] <= 32'b01000000011100010000001110110011;
ROM[4190] <= 32'b00000000011100000000001000110011;
ROM[4191] <= 32'b00000000001000000000000110110011;
ROM[4192] <= 32'b00010000110000000000000011101111;
ROM[4193] <= 32'b11111111110000010000000100010011;
ROM[4194] <= 32'b00000000000000010010001110000011;
ROM[4195] <= 32'b00000000011101100010000000100011;
ROM[4196] <= 32'b00000100010000000000001110010011;
ROM[4197] <= 32'b00000000011100010010000000100011;
ROM[4198] <= 32'b00000000010000010000000100010011;
ROM[4199] <= 32'b00000111110000000000001110010011;
ROM[4200] <= 32'b00000000011100010010000000100011;
ROM[4201] <= 32'b00000000010000010000000100010011;
ROM[4202] <= 32'b00000100011000000000001110010011;
ROM[4203] <= 32'b00000000011100010010000000100011;
ROM[4204] <= 32'b00000000010000010000000100010011;
ROM[4205] <= 32'b00000100001100000000001110010011;
ROM[4206] <= 32'b00000000011100010010000000100011;
ROM[4207] <= 32'b00000000010000010000000100010011;
ROM[4208] <= 32'b00000100001100000000001110010011;
ROM[4209] <= 32'b00000000011100010010000000100011;
ROM[4210] <= 32'b00000000010000010000000100010011;
ROM[4211] <= 32'b00000100001100000000001110010011;
ROM[4212] <= 32'b00000000011100010010000000100011;
ROM[4213] <= 32'b00000000010000010000000100010011;
ROM[4214] <= 32'b00000100011000000000001110010011;
ROM[4215] <= 32'b00000000011100010010000000100011;
ROM[4216] <= 32'b00000000010000010000000100010011;
ROM[4217] <= 32'b00000111110000000000001110010011;
ROM[4218] <= 32'b00000000011100010010000000100011;
ROM[4219] <= 32'b00000000010000010000000100010011;
ROM[4220] <= 32'b00000000000000000100001110110111;
ROM[4221] <= 32'b00100011110000111000001110010011;
ROM[4222] <= 32'b00000000111000111000001110110011;
ROM[4223] <= 32'b00000000011100010010000000100011;
ROM[4224] <= 32'b00000000010000010000000100010011;
ROM[4225] <= 32'b00000000001100010010000000100011;
ROM[4226] <= 32'b00000000010000010000000100010011;
ROM[4227] <= 32'b00000000010000010010000000100011;
ROM[4228] <= 32'b00000000010000010000000100010011;
ROM[4229] <= 32'b00000000010100010010000000100011;
ROM[4230] <= 32'b00000000010000010000000100010011;
ROM[4231] <= 32'b00000000011000010010000000100011;
ROM[4232] <= 32'b00000000010000010000000100010011;
ROM[4233] <= 32'b00000001010000000000001110010011;
ROM[4234] <= 32'b00000010000000111000001110010011;
ROM[4235] <= 32'b01000000011100010000001110110011;
ROM[4236] <= 32'b00000000011100000000001000110011;
ROM[4237] <= 32'b00000000001000000000000110110011;
ROM[4238] <= 32'b00000101010000000000000011101111;
ROM[4239] <= 32'b11111111110000010000000100010011;
ROM[4240] <= 32'b00000000000000010010001110000011;
ROM[4241] <= 32'b00000000011101100010000000100011;
ROM[4242] <= 32'b00000000000000000000001110010011;
ROM[4243] <= 32'b00000000011100010010000000100011;
ROM[4244] <= 32'b00000000010000010000000100010011;
ROM[4245] <= 32'b00000001010000000000001110010011;
ROM[4246] <= 32'b01000000011100011000001110110011;
ROM[4247] <= 32'b00000000000000111010000010000011;
ROM[4248] <= 32'b11111111110000010000000100010011;
ROM[4249] <= 32'b00000000000000010010001110000011;
ROM[4250] <= 32'b00000000011100100010000000100011;
ROM[4251] <= 32'b00000000010000100000000100010011;
ROM[4252] <= 32'b00000001010000000000001110010011;
ROM[4253] <= 32'b01000000011100011000001110110011;
ROM[4254] <= 32'b00000000010000111010000110000011;
ROM[4255] <= 32'b00000000100000111010001000000011;
ROM[4256] <= 32'b00000000110000111010001010000011;
ROM[4257] <= 32'b00000001000000111010001100000011;
ROM[4258] <= 32'b00000000000000001000000011100111;
ROM[4259] <= 32'b00000000000000010010000000100011;
ROM[4260] <= 32'b00000000010000010000000100010011;
ROM[4261] <= 32'b00000000000000010010000000100011;
ROM[4262] <= 32'b00000000010000010000000100010011;
ROM[4263] <= 32'b00000000011100000000001110010011;
ROM[4264] <= 32'b00000000011100010010000000100011;
ROM[4265] <= 32'b00000000010000010000000100010011;
ROM[4266] <= 32'b00000000000000000100001110110111;
ROM[4267] <= 32'b00101111010000111000001110010011;
ROM[4268] <= 32'b00000000111000111000001110110011;
ROM[4269] <= 32'b00000000011100010010000000100011;
ROM[4270] <= 32'b00000000010000010000000100010011;
ROM[4271] <= 32'b00000000001100010010000000100011;
ROM[4272] <= 32'b00000000010000010000000100010011;
ROM[4273] <= 32'b00000000010000010010000000100011;
ROM[4274] <= 32'b00000000010000010000000100010011;
ROM[4275] <= 32'b00000000010100010010000000100011;
ROM[4276] <= 32'b00000000010000010000000100010011;
ROM[4277] <= 32'b00000000011000010010000000100011;
ROM[4278] <= 32'b00000000010000010000000100010011;
ROM[4279] <= 32'b00000001010000000000001110010011;
ROM[4280] <= 32'b00000000010000111000001110010011;
ROM[4281] <= 32'b01000000011100010000001110110011;
ROM[4282] <= 32'b00000000011100000000001000110011;
ROM[4283] <= 32'b00000000001000000000000110110011;
ROM[4284] <= 32'b10010101000011111100000011101111;
ROM[4285] <= 32'b11111111110000010000000100010011;
ROM[4286] <= 32'b00000000000000010010001110000011;
ROM[4287] <= 32'b00000000011100011010000000100011;
ROM[4288] <= 32'b00000000000000100010001110000011;
ROM[4289] <= 32'b00000000011100010010000000100011;
ROM[4290] <= 32'b00000000010000010000000100010011;
ROM[4291] <= 32'b00000000000000100010001110000011;
ROM[4292] <= 32'b00000000011100010010000000100011;
ROM[4293] <= 32'b00000000010000010000000100010011;
ROM[4294] <= 32'b11111111110000010000000100010011;
ROM[4295] <= 32'b00000000000000010010001110000011;
ROM[4296] <= 32'b11111111110000010000000100010011;
ROM[4297] <= 32'b00000000000000010010010000000011;
ROM[4298] <= 32'b00000000011101000000001110110011;
ROM[4299] <= 32'b00000000011100010010000000100011;
ROM[4300] <= 32'b00000000010000010000000100010011;
ROM[4301] <= 32'b00000000000000100010001110000011;
ROM[4302] <= 32'b00000000011100010010000000100011;
ROM[4303] <= 32'b00000000010000010000000100010011;
ROM[4304] <= 32'b11111111110000010000000100010011;
ROM[4305] <= 32'b00000000000000010010001110000011;
ROM[4306] <= 32'b11111111110000010000000100010011;
ROM[4307] <= 32'b00000000000000010010010000000011;
ROM[4308] <= 32'b00000000011101000000001110110011;
ROM[4309] <= 32'b00000000011100010010000000100011;
ROM[4310] <= 32'b00000000010000010000000100010011;
ROM[4311] <= 32'b00000000000000100010001110000011;
ROM[4312] <= 32'b00000000011100010010000000100011;
ROM[4313] <= 32'b00000000010000010000000100010011;
ROM[4314] <= 32'b11111111110000010000000100010011;
ROM[4315] <= 32'b00000000000000010010001110000011;
ROM[4316] <= 32'b11111111110000010000000100010011;
ROM[4317] <= 32'b00000000000000010010010000000011;
ROM[4318] <= 32'b00000000011101000000001110110011;
ROM[4319] <= 32'b00000000011100010010000000100011;
ROM[4320] <= 32'b00000000010000010000000100010011;
ROM[4321] <= 32'b11111111110000010000000100010011;
ROM[4322] <= 32'b00000000000000010010001110000011;
ROM[4323] <= 32'b00000000011100011010001000100011;
ROM[4324] <= 32'b00000000010000011010001110000011;
ROM[4325] <= 32'b00000000011100010010000000100011;
ROM[4326] <= 32'b00000000010000010000000100010011;
ROM[4327] <= 32'b00001001000001101010001110000011;
ROM[4328] <= 32'b00000000011100010010000000100011;
ROM[4329] <= 32'b00000000010000010000000100010011;
ROM[4330] <= 32'b11111111110000010000000100010011;
ROM[4331] <= 32'b00000000000000010010001110000011;
ROM[4332] <= 32'b11111111110000010000000100010011;
ROM[4333] <= 32'b00000000000000010010010000000011;
ROM[4334] <= 32'b00000000011101000000001110110011;
ROM[4335] <= 32'b00000000011100010010000000100011;
ROM[4336] <= 32'b00000000010000010000000100010011;
ROM[4337] <= 32'b00000000000000011010001110000011;
ROM[4338] <= 32'b00000000011100010010000000100011;
ROM[4339] <= 32'b00000000010000010000000100010011;
ROM[4340] <= 32'b11111111110000010000000100010011;
ROM[4341] <= 32'b00000000000000010010001110000011;
ROM[4342] <= 32'b00000000011101100010000000100011;
ROM[4343] <= 32'b11111111110000010000000100010011;
ROM[4344] <= 32'b00000000000000010010001110000011;
ROM[4345] <= 32'b00000000000000111000001100010011;
ROM[4346] <= 32'b00000000000001100010001110000011;
ROM[4347] <= 32'b00000000011100010010000000100011;
ROM[4348] <= 32'b00000000010000010000000100010011;
ROM[4349] <= 32'b11111111110000010000000100010011;
ROM[4350] <= 32'b00000000000000010010001110000011;
ROM[4351] <= 32'b00000000110100110000010000110011;
ROM[4352] <= 32'b00000000011101000010000000100011;
ROM[4353] <= 32'b00000000000000000000001110010011;
ROM[4354] <= 32'b00000000011100010010000000100011;
ROM[4355] <= 32'b00000000010000010000000100010011;
ROM[4356] <= 32'b00000000000000011010001110000011;
ROM[4357] <= 32'b00000000011100010010000000100011;
ROM[4358] <= 32'b00000000010000010000000100010011;
ROM[4359] <= 32'b11111111110000010000000100010011;
ROM[4360] <= 32'b00000000000000010010001110000011;
ROM[4361] <= 32'b11111111110000010000000100010011;
ROM[4362] <= 32'b00000000000000010010010000000011;
ROM[4363] <= 32'b00000000011101000000001110110011;
ROM[4364] <= 32'b00000000011100010010000000100011;
ROM[4365] <= 32'b00000000010000010000000100010011;
ROM[4366] <= 32'b00000000010000100010001110000011;
ROM[4367] <= 32'b00000000011100010010000000100011;
ROM[4368] <= 32'b00000000010000010000000100010011;
ROM[4369] <= 32'b11111111110000010000000100010011;
ROM[4370] <= 32'b00000000000000010010001110000011;
ROM[4371] <= 32'b00000000011101100010000000100011;
ROM[4372] <= 32'b11111111110000010000000100010011;
ROM[4373] <= 32'b00000000000000010010001110000011;
ROM[4374] <= 32'b00000000000000111000001100010011;
ROM[4375] <= 32'b00000000000001100010001110000011;
ROM[4376] <= 32'b00000000011100010010000000100011;
ROM[4377] <= 32'b00000000010000010000000100010011;
ROM[4378] <= 32'b11111111110000010000000100010011;
ROM[4379] <= 32'b00000000000000010010001110000011;
ROM[4380] <= 32'b00000000110100110000010000110011;
ROM[4381] <= 32'b00000000011101000010000000100011;
ROM[4382] <= 32'b00000000010000000000001110010011;
ROM[4383] <= 32'b00000000011100010010000000100011;
ROM[4384] <= 32'b00000000010000010000000100010011;
ROM[4385] <= 32'b00000000000000011010001110000011;
ROM[4386] <= 32'b00000000011100010010000000100011;
ROM[4387] <= 32'b00000000010000010000000100010011;
ROM[4388] <= 32'b11111111110000010000000100010011;
ROM[4389] <= 32'b00000000000000010010001110000011;
ROM[4390] <= 32'b11111111110000010000000100010011;
ROM[4391] <= 32'b00000000000000010010010000000011;
ROM[4392] <= 32'b00000000011101000000001110110011;
ROM[4393] <= 32'b00000000011100010010000000100011;
ROM[4394] <= 32'b00000000010000010000000100010011;
ROM[4395] <= 32'b00000000100000100010001110000011;
ROM[4396] <= 32'b00000000011100010010000000100011;
ROM[4397] <= 32'b00000000010000010000000100010011;
ROM[4398] <= 32'b11111111110000010000000100010011;
ROM[4399] <= 32'b00000000000000010010001110000011;
ROM[4400] <= 32'b00000000011101100010000000100011;
ROM[4401] <= 32'b11111111110000010000000100010011;
ROM[4402] <= 32'b00000000000000010010001110000011;
ROM[4403] <= 32'b00000000000000111000001100010011;
ROM[4404] <= 32'b00000000000001100010001110000011;
ROM[4405] <= 32'b00000000011100010010000000100011;
ROM[4406] <= 32'b00000000010000010000000100010011;
ROM[4407] <= 32'b11111111110000010000000100010011;
ROM[4408] <= 32'b00000000000000010010001110000011;
ROM[4409] <= 32'b00000000110100110000010000110011;
ROM[4410] <= 32'b00000000011101000010000000100011;
ROM[4411] <= 32'b00000000100000000000001110010011;
ROM[4412] <= 32'b00000000011100010010000000100011;
ROM[4413] <= 32'b00000000010000010000000100010011;
ROM[4414] <= 32'b00000000000000011010001110000011;
ROM[4415] <= 32'b00000000011100010010000000100011;
ROM[4416] <= 32'b00000000010000010000000100010011;
ROM[4417] <= 32'b11111111110000010000000100010011;
ROM[4418] <= 32'b00000000000000010010001110000011;
ROM[4419] <= 32'b11111111110000010000000100010011;
ROM[4420] <= 32'b00000000000000010010010000000011;
ROM[4421] <= 32'b00000000011101000000001110110011;
ROM[4422] <= 32'b00000000011100010010000000100011;
ROM[4423] <= 32'b00000000010000010000000100010011;
ROM[4424] <= 32'b00000000110000100010001110000011;
ROM[4425] <= 32'b00000000011100010010000000100011;
ROM[4426] <= 32'b00000000010000010000000100010011;
ROM[4427] <= 32'b11111111110000010000000100010011;
ROM[4428] <= 32'b00000000000000010010001110000011;
ROM[4429] <= 32'b00000000011101100010000000100011;
ROM[4430] <= 32'b11111111110000010000000100010011;
ROM[4431] <= 32'b00000000000000010010001110000011;
ROM[4432] <= 32'b00000000000000111000001100010011;
ROM[4433] <= 32'b00000000000001100010001110000011;
ROM[4434] <= 32'b00000000011100010010000000100011;
ROM[4435] <= 32'b00000000010000010000000100010011;
ROM[4436] <= 32'b11111111110000010000000100010011;
ROM[4437] <= 32'b00000000000000010010001110000011;
ROM[4438] <= 32'b00000000110100110000010000110011;
ROM[4439] <= 32'b00000000011101000010000000100011;
ROM[4440] <= 32'b00000000110000000000001110010011;
ROM[4441] <= 32'b00000000011100010010000000100011;
ROM[4442] <= 32'b00000000010000010000000100010011;
ROM[4443] <= 32'b00000000000000011010001110000011;
ROM[4444] <= 32'b00000000011100010010000000100011;
ROM[4445] <= 32'b00000000010000010000000100010011;
ROM[4446] <= 32'b11111111110000010000000100010011;
ROM[4447] <= 32'b00000000000000010010001110000011;
ROM[4448] <= 32'b11111111110000010000000100010011;
ROM[4449] <= 32'b00000000000000010010010000000011;
ROM[4450] <= 32'b00000000011101000000001110110011;
ROM[4451] <= 32'b00000000011100010010000000100011;
ROM[4452] <= 32'b00000000010000010000000100010011;
ROM[4453] <= 32'b00000001000000100010001110000011;
ROM[4454] <= 32'b00000000011100010010000000100011;
ROM[4455] <= 32'b00000000010000010000000100010011;
ROM[4456] <= 32'b11111111110000010000000100010011;
ROM[4457] <= 32'b00000000000000010010001110000011;
ROM[4458] <= 32'b00000000011101100010000000100011;
ROM[4459] <= 32'b11111111110000010000000100010011;
ROM[4460] <= 32'b00000000000000010010001110000011;
ROM[4461] <= 32'b00000000000000111000001100010011;
ROM[4462] <= 32'b00000000000001100010001110000011;
ROM[4463] <= 32'b00000000011100010010000000100011;
ROM[4464] <= 32'b00000000010000010000000100010011;
ROM[4465] <= 32'b11111111110000010000000100010011;
ROM[4466] <= 32'b00000000000000010010001110000011;
ROM[4467] <= 32'b00000000110100110000010000110011;
ROM[4468] <= 32'b00000000011101000010000000100011;
ROM[4469] <= 32'b00000001000000000000001110010011;
ROM[4470] <= 32'b00000000011100010010000000100011;
ROM[4471] <= 32'b00000000010000010000000100010011;
ROM[4472] <= 32'b00000000000000011010001110000011;
ROM[4473] <= 32'b00000000011100010010000000100011;
ROM[4474] <= 32'b00000000010000010000000100010011;
ROM[4475] <= 32'b11111111110000010000000100010011;
ROM[4476] <= 32'b00000000000000010010001110000011;
ROM[4477] <= 32'b11111111110000010000000100010011;
ROM[4478] <= 32'b00000000000000010010010000000011;
ROM[4479] <= 32'b00000000011101000000001110110011;
ROM[4480] <= 32'b00000000011100010010000000100011;
ROM[4481] <= 32'b00000000010000010000000100010011;
ROM[4482] <= 32'b00000001010000100010001110000011;
ROM[4483] <= 32'b00000000011100010010000000100011;
ROM[4484] <= 32'b00000000010000010000000100010011;
ROM[4485] <= 32'b11111111110000010000000100010011;
ROM[4486] <= 32'b00000000000000010010001110000011;
ROM[4487] <= 32'b00000000011101100010000000100011;
ROM[4488] <= 32'b11111111110000010000000100010011;
ROM[4489] <= 32'b00000000000000010010001110000011;
ROM[4490] <= 32'b00000000000000111000001100010011;
ROM[4491] <= 32'b00000000000001100010001110000011;
ROM[4492] <= 32'b00000000011100010010000000100011;
ROM[4493] <= 32'b00000000010000010000000100010011;
ROM[4494] <= 32'b11111111110000010000000100010011;
ROM[4495] <= 32'b00000000000000010010001110000011;
ROM[4496] <= 32'b00000000110100110000010000110011;
ROM[4497] <= 32'b00000000011101000010000000100011;
ROM[4498] <= 32'b00000001010000000000001110010011;
ROM[4499] <= 32'b00000000011100010010000000100011;
ROM[4500] <= 32'b00000000010000010000000100010011;
ROM[4501] <= 32'b00000000000000011010001110000011;
ROM[4502] <= 32'b00000000011100010010000000100011;
ROM[4503] <= 32'b00000000010000010000000100010011;
ROM[4504] <= 32'b11111111110000010000000100010011;
ROM[4505] <= 32'b00000000000000010010001110000011;
ROM[4506] <= 32'b11111111110000010000000100010011;
ROM[4507] <= 32'b00000000000000010010010000000011;
ROM[4508] <= 32'b00000000011101000000001110110011;
ROM[4509] <= 32'b00000000011100010010000000100011;
ROM[4510] <= 32'b00000000010000010000000100010011;
ROM[4511] <= 32'b00000001100000100010001110000011;
ROM[4512] <= 32'b00000000011100010010000000100011;
ROM[4513] <= 32'b00000000010000010000000100010011;
ROM[4514] <= 32'b11111111110000010000000100010011;
ROM[4515] <= 32'b00000000000000010010001110000011;
ROM[4516] <= 32'b00000000011101100010000000100011;
ROM[4517] <= 32'b11111111110000010000000100010011;
ROM[4518] <= 32'b00000000000000010010001110000011;
ROM[4519] <= 32'b00000000000000111000001100010011;
ROM[4520] <= 32'b00000000000001100010001110000011;
ROM[4521] <= 32'b00000000011100010010000000100011;
ROM[4522] <= 32'b00000000010000010000000100010011;
ROM[4523] <= 32'b11111111110000010000000100010011;
ROM[4524] <= 32'b00000000000000010010001110000011;
ROM[4525] <= 32'b00000000110100110000010000110011;
ROM[4526] <= 32'b00000000011101000010000000100011;
ROM[4527] <= 32'b00000001100000000000001110010011;
ROM[4528] <= 32'b00000000011100010010000000100011;
ROM[4529] <= 32'b00000000010000010000000100010011;
ROM[4530] <= 32'b00000000000000011010001110000011;
ROM[4531] <= 32'b00000000011100010010000000100011;
ROM[4532] <= 32'b00000000010000010000000100010011;
ROM[4533] <= 32'b11111111110000010000000100010011;
ROM[4534] <= 32'b00000000000000010010001110000011;
ROM[4535] <= 32'b11111111110000010000000100010011;
ROM[4536] <= 32'b00000000000000010010010000000011;
ROM[4537] <= 32'b00000000011101000000001110110011;
ROM[4538] <= 32'b00000000011100010010000000100011;
ROM[4539] <= 32'b00000000010000010000000100010011;
ROM[4540] <= 32'b00000001110000100010001110000011;
ROM[4541] <= 32'b00000000011100010010000000100011;
ROM[4542] <= 32'b00000000010000010000000100010011;
ROM[4543] <= 32'b11111111110000010000000100010011;
ROM[4544] <= 32'b00000000000000010010001110000011;
ROM[4545] <= 32'b00000000011101100010000000100011;
ROM[4546] <= 32'b11111111110000010000000100010011;
ROM[4547] <= 32'b00000000000000010010001110000011;
ROM[4548] <= 32'b00000000000000111000001100010011;
ROM[4549] <= 32'b00000000000001100010001110000011;
ROM[4550] <= 32'b00000000011100010010000000100011;
ROM[4551] <= 32'b00000000010000010000000100010011;
ROM[4552] <= 32'b11111111110000010000000100010011;
ROM[4553] <= 32'b00000000000000010010001110000011;
ROM[4554] <= 32'b00000000110100110000010000110011;
ROM[4555] <= 32'b00000000011101000010000000100011;
ROM[4556] <= 32'b00000000000000000000001110010011;
ROM[4557] <= 32'b00000000011100010010000000100011;
ROM[4558] <= 32'b00000000010000010000000100010011;
ROM[4559] <= 32'b00000001010000000000001110010011;
ROM[4560] <= 32'b01000000011100011000001110110011;
ROM[4561] <= 32'b00000000000000111010000010000011;
ROM[4562] <= 32'b11111111110000010000000100010011;
ROM[4563] <= 32'b00000000000000010010001110000011;
ROM[4564] <= 32'b00000000011100100010000000100011;
ROM[4565] <= 32'b00000000010000100000000100010011;
ROM[4566] <= 32'b00000001010000000000001110010011;
ROM[4567] <= 32'b01000000011100011000001110110011;
ROM[4568] <= 32'b00000000010000111010000110000011;
ROM[4569] <= 32'b00000000100000111010001000000011;
ROM[4570] <= 32'b00000000110000111010001010000011;
ROM[4571] <= 32'b00000001000000111010001100000011;
ROM[4572] <= 32'b00000000000000001000000011100111;
ROM[4573] <= 32'b00000000000000010010000000100011;
ROM[4574] <= 32'b00000000010000010000000100010011;
ROM[4575] <= 32'b00000000000000010010000000100011;
ROM[4576] <= 32'b00000000010000010000000100010011;
ROM[4577] <= 32'b00000000000000010010000000100011;
ROM[4578] <= 32'b00000000010000010000000100010011;
ROM[4579] <= 32'b00000000000000010010000000100011;
ROM[4580] <= 32'b00000000010000010000000100010011;
ROM[4581] <= 32'b00000000000000010010000000100011;
ROM[4582] <= 32'b00000000010000010000000100010011;
ROM[4583] <= 32'b00000000000000010010000000100011;
ROM[4584] <= 32'b00000000010000010000000100010011;
ROM[4585] <= 32'b00000000000000000000001110010011;
ROM[4586] <= 32'b00000000011100010010000000100011;
ROM[4587] <= 32'b00000000010000010000000100010011;
ROM[4588] <= 32'b11111111110000010000000100010011;
ROM[4589] <= 32'b00000000000000010010001110000011;
ROM[4590] <= 32'b00000000011100011010000000100011;
ROM[4591] <= 32'b00000000000000000000001110010011;
ROM[4592] <= 32'b00000000011100010010000000100011;
ROM[4593] <= 32'b00000000010000010000000100010011;
ROM[4594] <= 32'b11111111110000010000000100010011;
ROM[4595] <= 32'b00000000000000010010001110000011;
ROM[4596] <= 32'b00000000011100011010001000100011;
ROM[4597] <= 32'b00000000000000000000001110010011;
ROM[4598] <= 32'b00000000011100010010000000100011;
ROM[4599] <= 32'b00000000010000010000000100010011;
ROM[4600] <= 32'b11111111110000010000000100010011;
ROM[4601] <= 32'b00000000000000010010001110000011;
ROM[4602] <= 32'b00000000011100011010010000100011;
ROM[4603] <= 32'b00000000000000000000001110010011;
ROM[4604] <= 32'b00000000011100010010000000100011;
ROM[4605] <= 32'b00000000010000010000000100010011;
ROM[4606] <= 32'b11111111110000010000000100010011;
ROM[4607] <= 32'b00000000000000010010001110000011;
ROM[4608] <= 32'b00000000011100011010011000100011;
ROM[4609] <= 32'b00000000010000011010001110000011;
ROM[4610] <= 32'b00000000011100010010000000100011;
ROM[4611] <= 32'b00000000010000010000000100010011;
ROM[4612] <= 32'b00010011011000000000001110010011;
ROM[4613] <= 32'b00000000011100010010000000100011;
ROM[4614] <= 32'b00000000010000010000000100010011;
ROM[4615] <= 32'b11111111110000010000000100010011;
ROM[4616] <= 32'b00000000000000010010001110000011;
ROM[4617] <= 32'b11111111110000010000000100010011;
ROM[4618] <= 32'b00000000000000010010010000000011;
ROM[4619] <= 32'b00000000011101000010001110110011;
ROM[4620] <= 32'b00000000011100010010000000100011;
ROM[4621] <= 32'b00000000010000010000000100010011;
ROM[4622] <= 32'b11111111110000010000000100010011;
ROM[4623] <= 32'b00000000000000010010001110000011;
ROM[4624] <= 32'b01000000011100000000001110110011;
ROM[4625] <= 32'b00000000000100111000001110010011;
ROM[4626] <= 32'b00000000011100010010000000100011;
ROM[4627] <= 32'b00000000010000010000000100010011;
ROM[4628] <= 32'b11111111110000010000000100010011;
ROM[4629] <= 32'b00000000000000010010001110000011;
ROM[4630] <= 32'b00000000000000111000101001100011;
ROM[4631] <= 32'b00000000000000001000001110110111;
ROM[4632] <= 32'b11001110010000111000001110010011;
ROM[4633] <= 32'b00000000111000111000001110110011;
ROM[4634] <= 32'b00000000000000111000000011100111;
ROM[4635] <= 32'b00000000010000011010001110000011;
ROM[4636] <= 32'b00000000011100010010000000100011;
ROM[4637] <= 32'b00000000010000010000000100010011;
ROM[4638] <= 32'b00000010000000000000001110010011;
ROM[4639] <= 32'b00000000011100010010000000100011;
ROM[4640] <= 32'b00000000010000010000000100010011;
ROM[4641] <= 32'b00000000000000000101001110110111;
ROM[4642] <= 32'b10001101000000111000001110010011;
ROM[4643] <= 32'b00000000111000111000001110110011;
ROM[4644] <= 32'b00000000011100010010000000100011;
ROM[4645] <= 32'b00000000010000010000000100010011;
ROM[4646] <= 32'b00000000001100010010000000100011;
ROM[4647] <= 32'b00000000010000010000000100010011;
ROM[4648] <= 32'b00000000010000010010000000100011;
ROM[4649] <= 32'b00000000010000010000000100010011;
ROM[4650] <= 32'b00000000010100010010000000100011;
ROM[4651] <= 32'b00000000010000010000000100010011;
ROM[4652] <= 32'b00000000011000010010000000100011;
ROM[4653] <= 32'b00000000010000010000000100010011;
ROM[4654] <= 32'b00000001010000000000001110010011;
ROM[4655] <= 32'b00000000100000111000001110010011;
ROM[4656] <= 32'b01000000011100010000001110110011;
ROM[4657] <= 32'b00000000011100000000001000110011;
ROM[4658] <= 32'b00000000001000000000000110110011;
ROM[4659] <= 32'b10000100010011111110000011101111;
ROM[4660] <= 32'b11111111110000010000000100010011;
ROM[4661] <= 32'b00000000000000010010001110000011;
ROM[4662] <= 32'b00000000011100011010100000100011;
ROM[4663] <= 32'b00000001000000011010001110000011;
ROM[4664] <= 32'b00000000011100010010000000100011;
ROM[4665] <= 32'b00000000010000010000000100010011;
ROM[4666] <= 32'b00000000001100000000001110010011;
ROM[4667] <= 32'b00000000011100010010000000100011;
ROM[4668] <= 32'b00000000010000010000000100010011;
ROM[4669] <= 32'b00000000000000000101001110110111;
ROM[4670] <= 32'b10010100000000111000001110010011;
ROM[4671] <= 32'b00000000111000111000001110110011;
ROM[4672] <= 32'b00000000011100010010000000100011;
ROM[4673] <= 32'b00000000010000010000000100010011;
ROM[4674] <= 32'b00000000001100010010000000100011;
ROM[4675] <= 32'b00000000010000010000000100010011;
ROM[4676] <= 32'b00000000010000010010000000100011;
ROM[4677] <= 32'b00000000010000010000000100010011;
ROM[4678] <= 32'b00000000010100010010000000100011;
ROM[4679] <= 32'b00000000010000010000000100010011;
ROM[4680] <= 32'b00000000011000010010000000100011;
ROM[4681] <= 32'b00000000010000010000000100010011;
ROM[4682] <= 32'b00000001010000000000001110010011;
ROM[4683] <= 32'b00000000100000111000001110010011;
ROM[4684] <= 32'b01000000011100010000001110110011;
ROM[4685] <= 32'b00000000011100000000001000110011;
ROM[4686] <= 32'b00000000001000000000000110110011;
ROM[4687] <= 32'b11111101010111111101000011101111;
ROM[4688] <= 32'b11111111110000010000000100010011;
ROM[4689] <= 32'b00000000000000010010001110000011;
ROM[4690] <= 32'b00000000011100011010101000100011;
ROM[4691] <= 32'b00000001010000011010001110000011;
ROM[4692] <= 32'b00000000011100010010000000100011;
ROM[4693] <= 32'b00000000010000010000000100010011;
ROM[4694] <= 32'b00000000000100000000001110010011;
ROM[4695] <= 32'b00000000011100010010000000100011;
ROM[4696] <= 32'b00000000010000010000000100010011;
ROM[4697] <= 32'b11111111110000010000000100010011;
ROM[4698] <= 32'b00000000000000010010001110000011;
ROM[4699] <= 32'b11111111110000010000000100010011;
ROM[4700] <= 32'b00000000000000010010010000000011;
ROM[4701] <= 32'b00000000011101000010010010110011;
ROM[4702] <= 32'b00000000100000111010010100110011;
ROM[4703] <= 32'b00000000101001001000001110110011;
ROM[4704] <= 32'b00000000000100111000001110010011;
ROM[4705] <= 32'b00000000000100111111001110010011;
ROM[4706] <= 32'b00000000011100010010000000100011;
ROM[4707] <= 32'b00000000010000010000000100010011;
ROM[4708] <= 32'b11111111110000010000000100010011;
ROM[4709] <= 32'b00000000000000010010001110000011;
ROM[4710] <= 32'b00000000000000111000101001100011;
ROM[4711] <= 32'b00000000000000000111001110110111;
ROM[4712] <= 32'b10001110100000111000001110010011;
ROM[4713] <= 32'b00000000111000111000001110110011;
ROM[4714] <= 32'b00000000000000111000000011100111;
ROM[4715] <= 32'b01110101100100000001000011101111;
ROM[4716] <= 32'b00000000110000011010001110000011;
ROM[4717] <= 32'b00000000011100010010000000100011;
ROM[4718] <= 32'b00000000010000010000000100010011;
ROM[4719] <= 32'b00000000000000000000001110010011;
ROM[4720] <= 32'b00000000011100010010000000100011;
ROM[4721] <= 32'b00000000010000010000000100010011;
ROM[4722] <= 32'b11111111110000010000000100010011;
ROM[4723] <= 32'b00000000000000010010001110000011;
ROM[4724] <= 32'b11111111110000010000000100010011;
ROM[4725] <= 32'b00000000000000010010010000000011;
ROM[4726] <= 32'b00000000011101000010010010110011;
ROM[4727] <= 32'b00000000100000111010010100110011;
ROM[4728] <= 32'b00000000101001001000001110110011;
ROM[4729] <= 32'b00000000000100111000001110010011;
ROM[4730] <= 32'b00000000000100111111001110010011;
ROM[4731] <= 32'b00000000011100010010000000100011;
ROM[4732] <= 32'b00000000010000010000000100010011;
ROM[4733] <= 32'b11111111110000010000000100010011;
ROM[4734] <= 32'b00000000000000010010001110000011;
ROM[4735] <= 32'b00000000000000111000101001100011;
ROM[4736] <= 32'b00000000000000000111001110110111;
ROM[4737] <= 32'b11000011000000111000001110010011;
ROM[4738] <= 32'b00000000111000111000001110110011;
ROM[4739] <= 32'b00000000000000111000000011100111;
ROM[4740] <= 32'b00101110100000000010000011101111;
ROM[4741] <= 32'b00000000100000011010001110000011;
ROM[4742] <= 32'b00000000011100010010000000100011;
ROM[4743] <= 32'b00000000010000010000000100010011;
ROM[4744] <= 32'b00001000110001101010001110000011;
ROM[4745] <= 32'b00000000011100010010000000100011;
ROM[4746] <= 32'b00000000010000010000000100010011;
ROM[4747] <= 32'b11111111110000010000000100010011;
ROM[4748] <= 32'b00000000000000010010001110000011;
ROM[4749] <= 32'b11111111110000010000000100010011;
ROM[4750] <= 32'b00000000000000010010010000000011;
ROM[4751] <= 32'b00000000011101000000001110110011;
ROM[4752] <= 32'b00000000011100010010000000100011;
ROM[4753] <= 32'b00000000010000010000000100010011;
ROM[4754] <= 32'b00000000010000011010001110000011;
ROM[4755] <= 32'b00000000011100010010000000100011;
ROM[4756] <= 32'b00000000010000010000000100010011;
ROM[4757] <= 32'b11111111110000010000000100010011;
ROM[4758] <= 32'b00000000000000010010001110000011;
ROM[4759] <= 32'b00000000011101100010000000100011;
ROM[4760] <= 32'b11111111110000010000000100010011;
ROM[4761] <= 32'b00000000000000010010001110000011;
ROM[4762] <= 32'b00000000000000111000001100010011;
ROM[4763] <= 32'b00000000000001100010001110000011;
ROM[4764] <= 32'b00000000011100010010000000100011;
ROM[4765] <= 32'b00000000010000010000000100010011;
ROM[4766] <= 32'b11111111110000010000000100010011;
ROM[4767] <= 32'b00000000000000010010001110000011;
ROM[4768] <= 32'b00000000110100110000010000110011;
ROM[4769] <= 32'b00000000011101000010000000100011;
ROM[4770] <= 32'b00000000100000011010001110000011;
ROM[4771] <= 32'b00000000011100010010000000100011;
ROM[4772] <= 32'b00000000010000010000000100010011;
ROM[4773] <= 32'b00000000010000000000001110010011;
ROM[4774] <= 32'b00000000011100010010000000100011;
ROM[4775] <= 32'b00000000010000010000000100010011;
ROM[4776] <= 32'b11111111110000010000000100010011;
ROM[4777] <= 32'b00000000000000010010001110000011;
ROM[4778] <= 32'b11111111110000010000000100010011;
ROM[4779] <= 32'b00000000000000010010010000000011;
ROM[4780] <= 32'b00000000011101000000001110110011;
ROM[4781] <= 32'b00000000011100010010000000100011;
ROM[4782] <= 32'b00000000010000010000000100010011;
ROM[4783] <= 32'b11111111110000010000000100010011;
ROM[4784] <= 32'b00000000000000010010001110000011;
ROM[4785] <= 32'b00000000011100011010010000100011;
ROM[4786] <= 32'b00100011000000000010000011101111;
ROM[4787] <= 32'b00000000110000011010001110000011;
ROM[4788] <= 32'b00000000011100010010000000100011;
ROM[4789] <= 32'b00000000010000010000000100010011;
ROM[4790] <= 32'b00000000000100000000001110010011;
ROM[4791] <= 32'b00000000011100010010000000100011;
ROM[4792] <= 32'b00000000010000010000000100010011;
ROM[4793] <= 32'b11111111110000010000000100010011;
ROM[4794] <= 32'b00000000000000010010001110000011;
ROM[4795] <= 32'b11111111110000010000000100010011;
ROM[4796] <= 32'b00000000000000010010010000000011;
ROM[4797] <= 32'b00000000011101000000001110110011;
ROM[4798] <= 32'b00000000011100010010000000100011;
ROM[4799] <= 32'b00000000010000010000000100010011;
ROM[4800] <= 32'b11111111110000010000000100010011;
ROM[4801] <= 32'b00000000000000010010001110000011;
ROM[4802] <= 32'b00000000011100011010011000100011;
ROM[4803] <= 32'b00000000110000011010001110000011;
ROM[4804] <= 32'b00000000011100010010000000100011;
ROM[4805] <= 32'b00000000010000010000000100010011;
ROM[4806] <= 32'b00000000001100000000001110010011;
ROM[4807] <= 32'b00000000011100010010000000100011;
ROM[4808] <= 32'b00000000010000010000000100010011;
ROM[4809] <= 32'b00000000000000000101001110110111;
ROM[4810] <= 32'b10110111000000111000001110010011;
ROM[4811] <= 32'b00000000111000111000001110110011;
ROM[4812] <= 32'b00000000011100010010000000100011;
ROM[4813] <= 32'b00000000010000010000000100010011;
ROM[4814] <= 32'b00000000001100010010000000100011;
ROM[4815] <= 32'b00000000010000010000000100010011;
ROM[4816] <= 32'b00000000010000010010000000100011;
ROM[4817] <= 32'b00000000010000010000000100010011;
ROM[4818] <= 32'b00000000010100010010000000100011;
ROM[4819] <= 32'b00000000010000010000000100010011;
ROM[4820] <= 32'b00000000011000010010000000100011;
ROM[4821] <= 32'b00000000010000010000000100010011;
ROM[4822] <= 32'b00000001010000000000001110010011;
ROM[4823] <= 32'b00000000100000111000001110010011;
ROM[4824] <= 32'b01000000011100010000001110110011;
ROM[4825] <= 32'b00000000011100000000001000110011;
ROM[4826] <= 32'b00000000001000000000000110110011;
ROM[4827] <= 32'b11011010010111111101000011101111;
ROM[4828] <= 32'b11111111110000010000000100010011;
ROM[4829] <= 32'b00000000000000010010001110000011;
ROM[4830] <= 32'b00000000011100011010011000100011;
ROM[4831] <= 32'b01011000100100000001000011101111;
ROM[4832] <= 32'b00000000010000011010001110000011;
ROM[4833] <= 32'b00000000011100010010000000100011;
ROM[4834] <= 32'b00000000010000010000000100010011;
ROM[4835] <= 32'b00000000000100000000001110010011;
ROM[4836] <= 32'b00000000011100010010000000100011;
ROM[4837] <= 32'b00000000010000010000000100010011;
ROM[4838] <= 32'b11111111110000010000000100010011;
ROM[4839] <= 32'b00000000000000010010001110000011;
ROM[4840] <= 32'b11111111110000010000000100010011;
ROM[4841] <= 32'b00000000000000010010010000000011;
ROM[4842] <= 32'b00000000011101000000001110110011;
ROM[4843] <= 32'b00000000011100010010000000100011;
ROM[4844] <= 32'b00000000010000010000000100010011;
ROM[4845] <= 32'b11111111110000010000000100010011;
ROM[4846] <= 32'b00000000000000010010001110000011;
ROM[4847] <= 32'b00000000011100011010001000100011;
ROM[4848] <= 32'b00001100100000000011000011101111;
ROM[4849] <= 32'b00000000000000000000001110010011;
ROM[4850] <= 32'b00000000011100010010000000100011;
ROM[4851] <= 32'b00000000010000010000000100010011;
ROM[4852] <= 32'b00000001010000000000001110010011;
ROM[4853] <= 32'b01000000011100011000001110110011;
ROM[4854] <= 32'b00000000000000111010000010000011;
ROM[4855] <= 32'b11111111110000010000000100010011;
ROM[4856] <= 32'b00000000000000010010001110000011;
ROM[4857] <= 32'b00000000011100100010000000100011;
ROM[4858] <= 32'b00000000010000100000000100010011;
ROM[4859] <= 32'b00000001010000000000001110010011;
ROM[4860] <= 32'b01000000011100011000001110110011;
ROM[4861] <= 32'b00000000010000111010000110000011;
ROM[4862] <= 32'b00000000100000111010001000000011;
ROM[4863] <= 32'b00000000110000111010001010000011;
ROM[4864] <= 32'b00000001000000111010001100000011;
ROM[4865] <= 32'b00000000000000001000000011100111;
ROM[4866] <= 32'b00000000000000100010001110000011;
ROM[4867] <= 32'b00000000011100010010000000100011;
ROM[4868] <= 32'b00000000010000010000000100010011;
ROM[4869] <= 32'b00000010000000000000001110010011;
ROM[4870] <= 32'b00000000011100010010000000100011;
ROM[4871] <= 32'b00000000010000010000000100010011;
ROM[4872] <= 32'b11111111110000010000000100010011;
ROM[4873] <= 32'b00000000000000010010001110000011;
ROM[4874] <= 32'b11111111110000010000000100010011;
ROM[4875] <= 32'b00000000000000010010010000000011;
ROM[4876] <= 32'b00000000011101000010001110110011;
ROM[4877] <= 32'b00000000011100010010000000100011;
ROM[4878] <= 32'b00000000010000010000000100010011;
ROM[4879] <= 32'b00000000000000100010001110000011;
ROM[4880] <= 32'b00000000011100010010000000100011;
ROM[4881] <= 32'b00000000010000010000000100010011;
ROM[4882] <= 32'b00000111111000000000001110010011;
ROM[4883] <= 32'b00000000011100010010000000100011;
ROM[4884] <= 32'b00000000010000010000000100010011;
ROM[4885] <= 32'b11111111110000010000000100010011;
ROM[4886] <= 32'b00000000000000010010001110000011;
ROM[4887] <= 32'b11111111110000010000000100010011;
ROM[4888] <= 32'b00000000000000010010010000000011;
ROM[4889] <= 32'b00000000100000111010001110110011;
ROM[4890] <= 32'b00000000011100010010000000100011;
ROM[4891] <= 32'b00000000010000010000000100010011;
ROM[4892] <= 32'b11111111110000010000000100010011;
ROM[4893] <= 32'b00000000000000010010001110000011;
ROM[4894] <= 32'b11111111110000010000000100010011;
ROM[4895] <= 32'b00000000000000010010010000000011;
ROM[4896] <= 32'b00000000011101000110001110110011;
ROM[4897] <= 32'b00000000011100010010000000100011;
ROM[4898] <= 32'b00000000010000010000000100010011;
ROM[4899] <= 32'b11111111110000010000000100010011;
ROM[4900] <= 32'b00000000000000010010001110000011;
ROM[4901] <= 32'b00000000000000111000101001100011;
ROM[4902] <= 32'b00000000000000000111001110110111;
ROM[4903] <= 32'b11011011000000111000001110010011;
ROM[4904] <= 32'b00000000111000111000001110110011;
ROM[4905] <= 32'b00000000000000111000000011100111;
ROM[4906] <= 32'b00010101010000000010000011101111;
ROM[4907] <= 32'b00000000000000000000001110010011;
ROM[4908] <= 32'b00000000011100010010000000100011;
ROM[4909] <= 32'b00000000010000010000000100010011;
ROM[4910] <= 32'b11111111110000010000000100010011;
ROM[4911] <= 32'b00000000000000010010001110000011;
ROM[4912] <= 32'b00000000011100100010000000100011;
ROM[4913] <= 32'b00010011100000000010000011101111;
ROM[4914] <= 32'b00000000000000100010001110000011;
ROM[4915] <= 32'b00000000011100010010000000100011;
ROM[4916] <= 32'b00000000010000010000000100010011;
ROM[4917] <= 32'b00000000000000100010001110000011;
ROM[4918] <= 32'b00000000011100010010000000100011;
ROM[4919] <= 32'b00000000010000010000000100010011;
ROM[4920] <= 32'b11111111110000010000000100010011;
ROM[4921] <= 32'b00000000000000010010001110000011;
ROM[4922] <= 32'b11111111110000010000000100010011;
ROM[4923] <= 32'b00000000000000010010010000000011;
ROM[4924] <= 32'b00000000011101000000001110110011;
ROM[4925] <= 32'b00000000011100010010000000100011;
ROM[4926] <= 32'b00000000010000010000000100010011;
ROM[4927] <= 32'b00000000000000100010001110000011;
ROM[4928] <= 32'b00000000011100010010000000100011;
ROM[4929] <= 32'b00000000010000010000000100010011;
ROM[4930] <= 32'b11111111110000010000000100010011;
ROM[4931] <= 32'b00000000000000010010001110000011;
ROM[4932] <= 32'b11111111110000010000000100010011;
ROM[4933] <= 32'b00000000000000010010010000000011;
ROM[4934] <= 32'b00000000011101000000001110110011;
ROM[4935] <= 32'b00000000011100010010000000100011;
ROM[4936] <= 32'b00000000010000010000000100010011;
ROM[4937] <= 32'b00000000000000100010001110000011;
ROM[4938] <= 32'b00000000011100010010000000100011;
ROM[4939] <= 32'b00000000010000010000000100010011;
ROM[4940] <= 32'b11111111110000010000000100010011;
ROM[4941] <= 32'b00000000000000010010001110000011;
ROM[4942] <= 32'b11111111110000010000000100010011;
ROM[4943] <= 32'b00000000000000010010010000000011;
ROM[4944] <= 32'b00000000011101000000001110110011;
ROM[4945] <= 32'b00000000011100010010000000100011;
ROM[4946] <= 32'b00000000010000010000000100010011;
ROM[4947] <= 32'b11111111110000010000000100010011;
ROM[4948] <= 32'b00000000000000010010001110000011;
ROM[4949] <= 32'b00000000011100100010000000100011;
ROM[4950] <= 32'b00000000000000100010001110000011;
ROM[4951] <= 32'b00000000011100010010000000100011;
ROM[4952] <= 32'b00000000010000010000000100010011;
ROM[4953] <= 32'b00001001000001101010001110000011;
ROM[4954] <= 32'b00000000011100010010000000100011;
ROM[4955] <= 32'b00000000010000010000000100010011;
ROM[4956] <= 32'b11111111110000010000000100010011;
ROM[4957] <= 32'b00000000000000010010001110000011;
ROM[4958] <= 32'b11111111110000010000000100010011;
ROM[4959] <= 32'b00000000000000010010010000000011;
ROM[4960] <= 32'b00000000011101000000001110110011;
ROM[4961] <= 32'b00000000011100010010000000100011;
ROM[4962] <= 32'b00000000010000010000000100010011;
ROM[4963] <= 32'b11111111110000010000000100010011;
ROM[4964] <= 32'b00000000000000010010001110000011;
ROM[4965] <= 32'b00000000000000111000001100010011;
ROM[4966] <= 32'b00000000110100110000010000110011;
ROM[4967] <= 32'b00000000000001000010001110000011;
ROM[4968] <= 32'b00000000011100010010000000100011;
ROM[4969] <= 32'b00000000010000010000000100010011;
ROM[4970] <= 32'b00000001010000000000001110010011;
ROM[4971] <= 32'b01000000011100011000001110110011;
ROM[4972] <= 32'b00000000000000111010000010000011;
ROM[4973] <= 32'b11111111110000010000000100010011;
ROM[4974] <= 32'b00000000000000010010001110000011;
ROM[4975] <= 32'b00000000011100100010000000100011;
ROM[4976] <= 32'b00000000010000100000000100010011;
ROM[4977] <= 32'b00000001010000000000001110010011;
ROM[4978] <= 32'b01000000011100011000001110110011;
ROM[4979] <= 32'b00000000010000111010000110000011;
ROM[4980] <= 32'b00000000100000111010001000000011;
ROM[4981] <= 32'b00000000110000111010001010000011;
ROM[4982] <= 32'b00000001000000111010001100000011;
ROM[4983] <= 32'b00000000000000001000000011100111;
ROM[4984] <= 32'b00000000010000100010001110000011;
ROM[4985] <= 32'b00000000011100010010000000100011;
ROM[4986] <= 32'b00000000010000010000000100010011;
ROM[4987] <= 32'b11111111110000010000000100010011;
ROM[4988] <= 32'b00000000000000010010001110000011;
ROM[4989] <= 32'b00000110011101101010110000100011;
ROM[4990] <= 32'b00000000000000100010001110000011;
ROM[4991] <= 32'b00000000011100010010000000100011;
ROM[4992] <= 32'b00000000010000010000000100010011;
ROM[4993] <= 32'b11111111110000010000000100010011;
ROM[4994] <= 32'b00000000000000010010001110000011;
ROM[4995] <= 32'b00000110011101101010111000100011;
ROM[4996] <= 32'b00000000000000000000001110010011;
ROM[4997] <= 32'b00000000011100010010000000100011;
ROM[4998] <= 32'b00000000010000010000000100010011;
ROM[4999] <= 32'b00000001010000000000001110010011;
ROM[5000] <= 32'b01000000011100011000001110110011;
ROM[5001] <= 32'b00000000000000111010000010000011;
ROM[5002] <= 32'b11111111110000010000000100010011;
ROM[5003] <= 32'b00000000000000010010001110000011;
ROM[5004] <= 32'b00000000011100100010000000100011;
ROM[5005] <= 32'b00000000010000100000000100010011;
ROM[5006] <= 32'b00000001010000000000001110010011;
ROM[5007] <= 32'b01000000011100011000001110110011;
ROM[5008] <= 32'b00000000010000111010000110000011;
ROM[5009] <= 32'b00000000100000111010001000000011;
ROM[5010] <= 32'b00000000110000111010001010000011;
ROM[5011] <= 32'b00000001000000111010001100000011;
ROM[5012] <= 32'b00000000000000001000000011100111;
ROM[5013] <= 32'b00000000000000010010000000100011;
ROM[5014] <= 32'b00000000010000010000000100010011;
ROM[5015] <= 32'b00000000000100000000001110010011;
ROM[5016] <= 32'b00000000011100010010000000100011;
ROM[5017] <= 32'b00000000010000010000000100010011;
ROM[5018] <= 32'b11111111110000010000000100010011;
ROM[5019] <= 32'b00000000000000010010001110000011;
ROM[5020] <= 32'b00000000011100011010000000100011;
ROM[5021] <= 32'b00000000010000100010001110000011;
ROM[5022] <= 32'b00000000011100010010000000100011;
ROM[5023] <= 32'b00000000010000010000000100010011;
ROM[5024] <= 32'b00000000000000000000001110010011;
ROM[5025] <= 32'b00000000011100010010000000100011;
ROM[5026] <= 32'b00000000010000010000000100010011;
ROM[5027] <= 32'b11111111110000010000000100010011;
ROM[5028] <= 32'b00000000000000010010001110000011;
ROM[5029] <= 32'b11111111110000010000000100010011;
ROM[5030] <= 32'b00000000000000010010010000000011;
ROM[5031] <= 32'b00000000100000111010001110110011;
ROM[5032] <= 32'b00000000011100010010000000100011;
ROM[5033] <= 32'b00000000010000010000000100010011;
ROM[5034] <= 32'b11111111110000010000000100010011;
ROM[5035] <= 32'b00000000000000010010001110000011;
ROM[5036] <= 32'b01000000011100000000001110110011;
ROM[5037] <= 32'b00000000000100111000001110010011;
ROM[5038] <= 32'b00000000011100010010000000100011;
ROM[5039] <= 32'b00000000010000010000000100010011;
ROM[5040] <= 32'b11111111110000010000000100010011;
ROM[5041] <= 32'b00000000000000010010001110000011;
ROM[5042] <= 32'b00000000000000111000101001100011;
ROM[5043] <= 32'b00000000000000001000001110110111;
ROM[5044] <= 32'b11101100000000111000001110010011;
ROM[5045] <= 32'b00000000111000111000001110110011;
ROM[5046] <= 32'b00000000000000111000000011100111;
ROM[5047] <= 32'b00000000000000011010001110000011;
ROM[5048] <= 32'b00000000011100010010000000100011;
ROM[5049] <= 32'b00000000010000010000000100010011;
ROM[5050] <= 32'b00000000000000100010001110000011;
ROM[5051] <= 32'b00000000011100010010000000100011;
ROM[5052] <= 32'b00000000010000010000000100010011;
ROM[5053] <= 32'b00000000000000000101001110110111;
ROM[5054] <= 32'b11110100000000111000001110010011;
ROM[5055] <= 32'b00000000111000111000001110110011;
ROM[5056] <= 32'b00000000011100010010000000100011;
ROM[5057] <= 32'b00000000010000010000000100010011;
ROM[5058] <= 32'b00000000001100010010000000100011;
ROM[5059] <= 32'b00000000010000010000000100010011;
ROM[5060] <= 32'b00000000010000010010000000100011;
ROM[5061] <= 32'b00000000010000010000000100010011;
ROM[5062] <= 32'b00000000010100010010000000100011;
ROM[5063] <= 32'b00000000010000010000000100010011;
ROM[5064] <= 32'b00000000011000010010000000100011;
ROM[5065] <= 32'b00000000010000010000000100010011;
ROM[5066] <= 32'b00000001010000000000001110010011;
ROM[5067] <= 32'b00000000100000111000001110010011;
ROM[5068] <= 32'b01000000011100010000001110110011;
ROM[5069] <= 32'b00000000011100000000001000110011;
ROM[5070] <= 32'b00000000001000000000000110110011;
ROM[5071] <= 32'b10000000110011111101000011101111;
ROM[5072] <= 32'b11111111110000010000000100010011;
ROM[5073] <= 32'b00000000000000010010001110000011;
ROM[5074] <= 32'b00000000011100011010000000100011;
ROM[5075] <= 32'b00000000010000100010001110000011;
ROM[5076] <= 32'b00000000011100010010000000100011;
ROM[5077] <= 32'b00000000010000010000000100010011;
ROM[5078] <= 32'b00000000000100000000001110010011;
ROM[5079] <= 32'b00000000011100010010000000100011;
ROM[5080] <= 32'b00000000010000010000000100010011;
ROM[5081] <= 32'b11111111110000010000000100010011;
ROM[5082] <= 32'b00000000000000010010001110000011;
ROM[5083] <= 32'b11111111110000010000000100010011;
ROM[5084] <= 32'b00000000000000010010010000000011;
ROM[5085] <= 32'b01000000011101000000001110110011;
ROM[5086] <= 32'b00000000011100010010000000100011;
ROM[5087] <= 32'b00000000010000010000000100010011;
ROM[5088] <= 32'b11111111110000010000000100010011;
ROM[5089] <= 32'b00000000000000010010001110000011;
ROM[5090] <= 32'b00000000011100100010001000100011;
ROM[5091] <= 32'b01011100010100000010000011101111;
ROM[5092] <= 32'b00000000000000011010001110000011;
ROM[5093] <= 32'b00000000011100010010000000100011;
ROM[5094] <= 32'b00000000010000010000000100010011;
ROM[5095] <= 32'b00000001010000000000001110010011;
ROM[5096] <= 32'b01000000011100011000001110110011;
ROM[5097] <= 32'b00000000000000111010000010000011;
ROM[5098] <= 32'b11111111110000010000000100010011;
ROM[5099] <= 32'b00000000000000010010001110000011;
ROM[5100] <= 32'b00000000011100100010000000100011;
ROM[5101] <= 32'b00000000010000100000000100010011;
ROM[5102] <= 32'b00000001010000000000001110010011;
ROM[5103] <= 32'b01000000011100011000001110110011;
ROM[5104] <= 32'b00000000010000111010000110000011;
ROM[5105] <= 32'b00000000100000111010001000000011;
ROM[5106] <= 32'b00000000110000111010001010000011;
ROM[5107] <= 32'b00000001000000111010001100000011;
ROM[5108] <= 32'b00000000000000001000000011100111;
ROM[5109] <= 32'b00000000000000010010000000100011;
ROM[5110] <= 32'b00000000010000010000000100010011;
ROM[5111] <= 32'b00000000000000010010000000100011;
ROM[5112] <= 32'b00000000010000010000000100010011;
ROM[5113] <= 32'b00000000000000010010000000100011;
ROM[5114] <= 32'b00000000010000010000000100010011;
ROM[5115] <= 32'b00000000000000010010000000100011;
ROM[5116] <= 32'b00000000010000010000000100010011;
ROM[5117] <= 32'b00000000000000010010000000100011;
ROM[5118] <= 32'b00000000010000010000000100010011;
ROM[5119] <= 32'b00000000000000010010000000100011;
ROM[5120] <= 32'b00000000010000010000000100010011;
ROM[5121] <= 32'b00000000000000010010000000100011;
ROM[5122] <= 32'b00000000010000010000000100010011;
ROM[5123] <= 32'b00000000000000010010000000100011;
ROM[5124] <= 32'b00000000010000010000000100010011;
ROM[5125] <= 32'b00000000000000010010000000100011;
ROM[5126] <= 32'b00000000010000010000000100010011;
ROM[5127] <= 32'b00000000000000010010000000100011;
ROM[5128] <= 32'b00000000010000010000000100010011;
ROM[5129] <= 32'b00000000000000010010000000100011;
ROM[5130] <= 32'b00000000010000010000000100010011;
ROM[5131] <= 32'b00000000000000010010000000100011;
ROM[5132] <= 32'b00000000010000010000000100010011;
ROM[5133] <= 32'b00000000000000010010000000100011;
ROM[5134] <= 32'b00000000010000010000000100010011;
ROM[5135] <= 32'b00000000000000010010000000100011;
ROM[5136] <= 32'b00000000010000010000000100010011;
ROM[5137] <= 32'b00000000000000010010000000100011;
ROM[5138] <= 32'b00000000010000010000000100010011;
ROM[5139] <= 32'b00000000000000010010000000100011;
ROM[5140] <= 32'b00000000010000010000000100010011;
ROM[5141] <= 32'b00000000000000010010000000100011;
ROM[5142] <= 32'b00000000010000010000000100010011;
ROM[5143] <= 32'b00001000000001101010001110000011;
ROM[5144] <= 32'b00000000011100010010000000100011;
ROM[5145] <= 32'b00000000010000010000000100010011;
ROM[5146] <= 32'b00001000000001101010001110000011;
ROM[5147] <= 32'b00000000011100010010000000100011;
ROM[5148] <= 32'b00000000010000010000000100010011;
ROM[5149] <= 32'b11111111110000010000000100010011;
ROM[5150] <= 32'b00000000000000010010001110000011;
ROM[5151] <= 32'b11111111110000010000000100010011;
ROM[5152] <= 32'b00000000000000010010010000000011;
ROM[5153] <= 32'b00000000011101000000001110110011;
ROM[5154] <= 32'b00000000011100010010000000100011;
ROM[5155] <= 32'b00000000010000010000000100010011;
ROM[5156] <= 32'b00001000000001101010001110000011;
ROM[5157] <= 32'b00000000011100010010000000100011;
ROM[5158] <= 32'b00000000010000010000000100010011;
ROM[5159] <= 32'b11111111110000010000000100010011;
ROM[5160] <= 32'b00000000000000010010001110000011;
ROM[5161] <= 32'b11111111110000010000000100010011;
ROM[5162] <= 32'b00000000000000010010010000000011;
ROM[5163] <= 32'b00000000011101000000001110110011;
ROM[5164] <= 32'b00000000011100010010000000100011;
ROM[5165] <= 32'b00000000010000010000000100010011;
ROM[5166] <= 32'b00001000000001101010001110000011;
ROM[5167] <= 32'b00000000011100010010000000100011;
ROM[5168] <= 32'b00000000010000010000000100010011;
ROM[5169] <= 32'b11111111110000010000000100010011;
ROM[5170] <= 32'b00000000000000010010001110000011;
ROM[5171] <= 32'b11111111110000010000000100010011;
ROM[5172] <= 32'b00000000000000010010010000000011;
ROM[5173] <= 32'b00000000011101000000001110110011;
ROM[5174] <= 32'b00000000011100010010000000100011;
ROM[5175] <= 32'b00000000010000010000000100010011;
ROM[5176] <= 32'b11111111110000010000000100010011;
ROM[5177] <= 32'b00000000000000010010001110000011;
ROM[5178] <= 32'b00001000011101101010001000100011;
ROM[5179] <= 32'b00001000010001101010001110000011;
ROM[5180] <= 32'b00000000011100010010000000100011;
ROM[5181] <= 32'b00000000010000010000000100010011;
ROM[5182] <= 32'b00001000110001101010001110000011;
ROM[5183] <= 32'b00000000011100010010000000100011;
ROM[5184] <= 32'b00000000010000010000000100010011;
ROM[5185] <= 32'b11111111110000010000000100010011;
ROM[5186] <= 32'b00000000000000010010001110000011;
ROM[5187] <= 32'b11111111110000010000000100010011;
ROM[5188] <= 32'b00000000000000010010010000000011;
ROM[5189] <= 32'b00000000011101000000001110110011;
ROM[5190] <= 32'b00000000011100010010000000100011;
ROM[5191] <= 32'b00000000010000010000000100010011;
ROM[5192] <= 32'b11111111110000010000000100010011;
ROM[5193] <= 32'b00000000000000010010001110000011;
ROM[5194] <= 32'b00000000000000111000001100010011;
ROM[5195] <= 32'b00000000110100110000010000110011;
ROM[5196] <= 32'b00000000000001000010001110000011;
ROM[5197] <= 32'b00000000011100010010000000100011;
ROM[5198] <= 32'b00000000010000010000000100010011;
ROM[5199] <= 32'b11111111110000010000000100010011;
ROM[5200] <= 32'b00000000000000010010001110000011;
ROM[5201] <= 32'b00000000011100011010001000100011;
ROM[5202] <= 32'b00001000100001101010001110000011;
ROM[5203] <= 32'b00000000011100010010000000100011;
ROM[5204] <= 32'b00000000010000010000000100010011;
ROM[5205] <= 32'b00000110010000000000001110010011;
ROM[5206] <= 32'b00000000011100010010000000100011;
ROM[5207] <= 32'b00000000010000010000000100010011;
ROM[5208] <= 32'b00000000000000000101001110110111;
ROM[5209] <= 32'b00011010110000111000001110010011;
ROM[5210] <= 32'b00000000111000111000001110110011;
ROM[5211] <= 32'b00000000011100010010000000100011;
ROM[5212] <= 32'b00000000010000010000000100010011;
ROM[5213] <= 32'b00000000001100010010000000100011;
ROM[5214] <= 32'b00000000010000010000000100010011;
ROM[5215] <= 32'b00000000010000010010000000100011;
ROM[5216] <= 32'b00000000010000010000000100010011;
ROM[5217] <= 32'b00000000010100010010000000100011;
ROM[5218] <= 32'b00000000010000010000000100010011;
ROM[5219] <= 32'b00000000011000010010000000100011;
ROM[5220] <= 32'b00000000010000010000000100010011;
ROM[5221] <= 32'b00000001010000000000001110010011;
ROM[5222] <= 32'b00000000100000111000001110010011;
ROM[5223] <= 32'b01000000011100010000001110110011;
ROM[5224] <= 32'b00000000011100000000001000110011;
ROM[5225] <= 32'b00000000001000000000000110110011;
ROM[5226] <= 32'b11011010000111111100000011101111;
ROM[5227] <= 32'b00000000010000011010001110000011;
ROM[5228] <= 32'b00000000011100010010000000100011;
ROM[5229] <= 32'b00000000010000010000000100010011;
ROM[5230] <= 32'b00000010000000000000001110010011;
ROM[5231] <= 32'b00000000011100010010000000100011;
ROM[5232] <= 32'b00000000010000010000000100010011;
ROM[5233] <= 32'b00000000000000000101001110110111;
ROM[5234] <= 32'b00100001000000111000001110010011;
ROM[5235] <= 32'b00000000111000111000001110110011;
ROM[5236] <= 32'b00000000011100010010000000100011;
ROM[5237] <= 32'b00000000010000010000000100010011;
ROM[5238] <= 32'b00000000001100010010000000100011;
ROM[5239] <= 32'b00000000010000010000000100010011;
ROM[5240] <= 32'b00000000010000010010000000100011;
ROM[5241] <= 32'b00000000010000010000000100010011;
ROM[5242] <= 32'b00000000010100010010000000100011;
ROM[5243] <= 32'b00000000010000010000000100010011;
ROM[5244] <= 32'b00000000011000010010000000100011;
ROM[5245] <= 32'b00000000010000010000000100010011;
ROM[5246] <= 32'b00000001010000000000001110010011;
ROM[5247] <= 32'b00000000100000111000001110010011;
ROM[5248] <= 32'b01000000011100010000001110110011;
ROM[5249] <= 32'b00000000011100000000001000110011;
ROM[5250] <= 32'b00000000001000000000000110110011;
ROM[5251] <= 32'b10001100000011111101000011101111;
ROM[5252] <= 32'b11111111110000010000000100010011;
ROM[5253] <= 32'b00000000000000010010001110000011;
ROM[5254] <= 32'b11111111110000010000000100010011;
ROM[5255] <= 32'b00000000000000010010010000000011;
ROM[5256] <= 32'b00000000011101000000001110110011;
ROM[5257] <= 32'b00000000011100010010000000100011;
ROM[5258] <= 32'b00000000010000010000000100010011;
ROM[5259] <= 32'b11111111110000010000000100010011;
ROM[5260] <= 32'b00000000000000010010001110000011;
ROM[5261] <= 32'b00000000011100011010010000100011;
ROM[5262] <= 32'b00000000010000011010001110000011;
ROM[5263] <= 32'b00000000011100010010000000100011;
ROM[5264] <= 32'b00000000010000010000000100010011;
ROM[5265] <= 32'b00000010000000000000001110010011;
ROM[5266] <= 32'b00000000011100010010000000100011;
ROM[5267] <= 32'b00000000010000010000000100010011;
ROM[5268] <= 32'b00000000000000000101001110110111;
ROM[5269] <= 32'b00101001110000111000001110010011;
ROM[5270] <= 32'b00000000111000111000001110110011;
ROM[5271] <= 32'b00000000011100010010000000100011;
ROM[5272] <= 32'b00000000010000010000000100010011;
ROM[5273] <= 32'b00000000001100010010000000100011;
ROM[5274] <= 32'b00000000010000010000000100010011;
ROM[5275] <= 32'b00000000010000010010000000100011;
ROM[5276] <= 32'b00000000010000010000000100010011;
ROM[5277] <= 32'b00000000010100010010000000100011;
ROM[5278] <= 32'b00000000010000010000000100010011;
ROM[5279] <= 32'b00000000011000010010000000100011;
ROM[5280] <= 32'b00000000010000010000000100010011;
ROM[5281] <= 32'b00000001010000000000001110010011;
ROM[5282] <= 32'b00000000100000111000001110010011;
ROM[5283] <= 32'b01000000011100010000001110110011;
ROM[5284] <= 32'b00000000011100000000001000110011;
ROM[5285] <= 32'b00000000001000000000000110110011;
ROM[5286] <= 32'b11100111100011111101000011101111;
ROM[5287] <= 32'b11111111110000010000000100010011;
ROM[5288] <= 32'b00000000000000010010001110000011;
ROM[5289] <= 32'b00000000011100011010000000100011;
ROM[5290] <= 32'b00000000000000000000001110010011;
ROM[5291] <= 32'b00000000011100010010000000100011;
ROM[5292] <= 32'b00000000010000010000000100010011;
ROM[5293] <= 32'b11111111110000010000000100010011;
ROM[5294] <= 32'b00000000000000010010001110000011;
ROM[5295] <= 32'b00000000011100011010011000100011;
ROM[5296] <= 32'b00000000000000100010001110000011;
ROM[5297] <= 32'b00000000011100010010000000100011;
ROM[5298] <= 32'b00000000010000010000000100010011;
ROM[5299] <= 32'b00000000000000000101001110110111;
ROM[5300] <= 32'b00110001100000111000001110010011;
ROM[5301] <= 32'b00000000111000111000001110110011;
ROM[5302] <= 32'b00000000011100010010000000100011;
ROM[5303] <= 32'b00000000010000010000000100010011;
ROM[5304] <= 32'b00000000001100010010000000100011;
ROM[5305] <= 32'b00000000010000010000000100010011;
ROM[5306] <= 32'b00000000010000010010000000100011;
ROM[5307] <= 32'b00000000010000010000000100010011;
ROM[5308] <= 32'b00000000010100010010000000100011;
ROM[5309] <= 32'b00000000010000010000000100010011;
ROM[5310] <= 32'b00000000011000010010000000100011;
ROM[5311] <= 32'b00000000010000010000000100010011;
ROM[5312] <= 32'b00000001010000000000001110010011;
ROM[5313] <= 32'b00000000010000111000001110010011;
ROM[5314] <= 32'b01000000011100010000001110110011;
ROM[5315] <= 32'b00000000011100000000001000110011;
ROM[5316] <= 32'b00000000001000000000000110110011;
ROM[5317] <= 32'b10001111010111111111000011101111;
ROM[5318] <= 32'b11111111110000010000000100010011;
ROM[5319] <= 32'b00000000000000010010001110000011;
ROM[5320] <= 32'b00000000011100011010100000100011;
ROM[5321] <= 32'b00000000110000011010001110000011;
ROM[5322] <= 32'b00000000011100010010000000100011;
ROM[5323] <= 32'b00000000010000010000000100010011;
ROM[5324] <= 32'b00000000011100000000001110010011;
ROM[5325] <= 32'b00000000011100010010000000100011;
ROM[5326] <= 32'b00000000010000010000000100010011;
ROM[5327] <= 32'b11111111110000010000000100010011;
ROM[5328] <= 32'b00000000000000010010001110000011;
ROM[5329] <= 32'b11111111110000010000000100010011;
ROM[5330] <= 32'b00000000000000010010010000000011;
ROM[5331] <= 32'b00000000011101000010001110110011;
ROM[5332] <= 32'b00000000011100010010000000100011;
ROM[5333] <= 32'b00000000010000010000000100010011;
ROM[5334] <= 32'b11111111110000010000000100010011;
ROM[5335] <= 32'b00000000000000010010001110000011;
ROM[5336] <= 32'b01000000011100000000001110110011;
ROM[5337] <= 32'b00000000000100111000001110010011;
ROM[5338] <= 32'b00000000011100010010000000100011;
ROM[5339] <= 32'b00000000010000010000000100010011;
ROM[5340] <= 32'b11111111110000010000000100010011;
ROM[5341] <= 32'b00000000000000010010001110000011;
ROM[5342] <= 32'b00000000000000111000101001100011;
ROM[5343] <= 32'b00000000000000001000001110110111;
ROM[5344] <= 32'b11100111110000111000001110010011;
ROM[5345] <= 32'b00000000111000111000001110110011;
ROM[5346] <= 32'b00000000000000111000000011100111;
ROM[5347] <= 32'b00000000000000000000001110010011;
ROM[5348] <= 32'b00000000011100010010000000100011;
ROM[5349] <= 32'b00000000010000010000000100010011;
ROM[5350] <= 32'b11111111110000010000000100010011;
ROM[5351] <= 32'b00000000000000010010001110000011;
ROM[5352] <= 32'b00000000011100011010101000100011;
ROM[5353] <= 32'b00000001010000011010001110000011;
ROM[5354] <= 32'b00000000011100010010000000100011;
ROM[5355] <= 32'b00000000010000010000000100010011;
ROM[5356] <= 32'b00000000011100000000001110010011;
ROM[5357] <= 32'b00000000011100010010000000100011;
ROM[5358] <= 32'b00000000010000010000000100010011;
ROM[5359] <= 32'b11111111110000010000000100010011;
ROM[5360] <= 32'b00000000000000010010001110000011;
ROM[5361] <= 32'b11111111110000010000000100010011;
ROM[5362] <= 32'b00000000000000010010010000000011;
ROM[5363] <= 32'b00000000011101000010001110110011;
ROM[5364] <= 32'b00000000011100010010000000100011;
ROM[5365] <= 32'b00000000010000010000000100010011;
ROM[5366] <= 32'b11111111110000010000000100010011;
ROM[5367] <= 32'b00000000000000010010001110000011;
ROM[5368] <= 32'b01000000011100000000001110110011;
ROM[5369] <= 32'b00000000000100111000001110010011;
ROM[5370] <= 32'b00000000011100010010000000100011;
ROM[5371] <= 32'b00000000010000010000000100010011;
ROM[5372] <= 32'b11111111110000010000000100010011;
ROM[5373] <= 32'b00000000000000010010001110000011;
ROM[5374] <= 32'b00000000000000111000101001100011;
ROM[5375] <= 32'b00000000000000000110001110110111;
ROM[5376] <= 32'b10100110110000111000001110010011;
ROM[5377] <= 32'b00000000111000111000001110110011;
ROM[5378] <= 32'b00000000000000111000000011100111;
ROM[5379] <= 32'b00000001010000011010001110000011;
ROM[5380] <= 32'b00000000011100010010000000100011;
ROM[5381] <= 32'b00000000010000010000000100010011;
ROM[5382] <= 32'b00000001010000011010001110000011;
ROM[5383] <= 32'b00000000011100010010000000100011;
ROM[5384] <= 32'b00000000010000010000000100010011;
ROM[5385] <= 32'b11111111110000010000000100010011;
ROM[5386] <= 32'b00000000000000010010001110000011;
ROM[5387] <= 32'b11111111110000010000000100010011;
ROM[5388] <= 32'b00000000000000010010010000000011;
ROM[5389] <= 32'b00000000011101000000001110110011;
ROM[5390] <= 32'b00000000011100010010000000100011;
ROM[5391] <= 32'b00000000010000010000000100010011;
ROM[5392] <= 32'b00000001010000011010001110000011;
ROM[5393] <= 32'b00000000011100010010000000100011;
ROM[5394] <= 32'b00000000010000010000000100010011;
ROM[5395] <= 32'b11111111110000010000000100010011;
ROM[5396] <= 32'b00000000000000010010001110000011;
ROM[5397] <= 32'b11111111110000010000000100010011;
ROM[5398] <= 32'b00000000000000010010010000000011;
ROM[5399] <= 32'b00000000011101000000001110110011;
ROM[5400] <= 32'b00000000011100010010000000100011;
ROM[5401] <= 32'b00000000010000010000000100010011;
ROM[5402] <= 32'b00000001010000011010001110000011;
ROM[5403] <= 32'b00000000011100010010000000100011;
ROM[5404] <= 32'b00000000010000010000000100010011;
ROM[5405] <= 32'b11111111110000010000000100010011;
ROM[5406] <= 32'b00000000000000010010001110000011;
ROM[5407] <= 32'b11111111110000010000000100010011;
ROM[5408] <= 32'b00000000000000010010010000000011;
ROM[5409] <= 32'b00000000011101000000001110110011;
ROM[5410] <= 32'b00000000011100010010000000100011;
ROM[5411] <= 32'b00000000010000010000000100010011;
ROM[5412] <= 32'b11111111110000010000000100010011;
ROM[5413] <= 32'b00000000000000010010001110000011;
ROM[5414] <= 32'b00000010011100011010111000100011;
ROM[5415] <= 32'b00000011110000011010001110000011;
ROM[5416] <= 32'b00000000011100010010000000100011;
ROM[5417] <= 32'b00000000010000010000000100010011;
ROM[5418] <= 32'b00000001000000011010001110000011;
ROM[5419] <= 32'b00000000011100010010000000100011;
ROM[5420] <= 32'b00000000010000010000000100010011;
ROM[5421] <= 32'b11111111110000010000000100010011;
ROM[5422] <= 32'b00000000000000010010001110000011;
ROM[5423] <= 32'b11111111110000010000000100010011;
ROM[5424] <= 32'b00000000000000010010010000000011;
ROM[5425] <= 32'b00000000011101000000001110110011;
ROM[5426] <= 32'b00000000011100010010000000100011;
ROM[5427] <= 32'b00000000010000010000000100010011;
ROM[5428] <= 32'b11111111110000010000000100010011;
ROM[5429] <= 32'b00000000000000010010001110000011;
ROM[5430] <= 32'b00000000000000111000001100010011;
ROM[5431] <= 32'b00000000110100110000010000110011;
ROM[5432] <= 32'b00000000000001000010001110000011;
ROM[5433] <= 32'b00000000011100010010000000100011;
ROM[5434] <= 32'b00000000010000010000000100010011;
ROM[5435] <= 32'b11111111110000010000000100010011;
ROM[5436] <= 32'b00000000000000010010001110000011;
ROM[5437] <= 32'b00000000011100011010110000100011;
ROM[5438] <= 32'b00000000100000011010001110000011;
ROM[5439] <= 32'b00000000011100010010000000100011;
ROM[5440] <= 32'b00000000010000010000000100010011;
ROM[5441] <= 32'b00000000100000011010001110000011;
ROM[5442] <= 32'b00000000011100010010000000100011;
ROM[5443] <= 32'b00000000010000010000000100010011;
ROM[5444] <= 32'b11111111110000010000000100010011;
ROM[5445] <= 32'b00000000000000010010001110000011;
ROM[5446] <= 32'b11111111110000010000000100010011;
ROM[5447] <= 32'b00000000000000010010010000000011;
ROM[5448] <= 32'b00000000011101000000001110110011;
ROM[5449] <= 32'b00000000011100010010000000100011;
ROM[5450] <= 32'b00000000010000010000000100010011;
ROM[5451] <= 32'b00000000100000011010001110000011;
ROM[5452] <= 32'b00000000011100010010000000100011;
ROM[5453] <= 32'b00000000010000010000000100010011;
ROM[5454] <= 32'b11111111110000010000000100010011;
ROM[5455] <= 32'b00000000000000010010001110000011;
ROM[5456] <= 32'b11111111110000010000000100010011;
ROM[5457] <= 32'b00000000000000010010010000000011;
ROM[5458] <= 32'b00000000011101000000001110110011;
ROM[5459] <= 32'b00000000011100010010000000100011;
ROM[5460] <= 32'b00000000010000010000000100010011;
ROM[5461] <= 32'b00000000100000011010001110000011;
ROM[5462] <= 32'b00000000011100010010000000100011;
ROM[5463] <= 32'b00000000010000010000000100010011;
ROM[5464] <= 32'b11111111110000010000000100010011;
ROM[5465] <= 32'b00000000000000010010001110000011;
ROM[5466] <= 32'b11111111110000010000000100010011;
ROM[5467] <= 32'b00000000000000010010010000000011;
ROM[5468] <= 32'b00000000011101000000001110110011;
ROM[5469] <= 32'b00000000011100010010000000100011;
ROM[5470] <= 32'b00000000010000010000000100010011;
ROM[5471] <= 32'b11111111110000010000000100010011;
ROM[5472] <= 32'b00000000000000010010001110000011;
ROM[5473] <= 32'b00000100011100011010000000100011;
ROM[5474] <= 32'b00000100000000011010001110000011;
ROM[5475] <= 32'b00000000011100010010000000100011;
ROM[5476] <= 32'b00000000010000010000000100010011;
ROM[5477] <= 32'b00000111010001101010001110000011;
ROM[5478] <= 32'b00000000011100010010000000100011;
ROM[5479] <= 32'b00000000010000010000000100010011;
ROM[5480] <= 32'b11111111110000010000000100010011;
ROM[5481] <= 32'b00000000000000010010001110000011;
ROM[5482] <= 32'b11111111110000010000000100010011;
ROM[5483] <= 32'b00000000000000010010010000000011;
ROM[5484] <= 32'b00000000011101000000001110110011;
ROM[5485] <= 32'b00000000011100010010000000100011;
ROM[5486] <= 32'b00000000010000010000000100010011;
ROM[5487] <= 32'b11111111110000010000000100010011;
ROM[5488] <= 32'b00000000000000010010001110000011;
ROM[5489] <= 32'b00000000000000111000001100010011;
ROM[5490] <= 32'b00000000110100110000010000110011;
ROM[5491] <= 32'b00000000000001000010001110000011;
ROM[5492] <= 32'b00000000011100010010000000100011;
ROM[5493] <= 32'b00000000010000010000000100010011;
ROM[5494] <= 32'b11111111110000010000000100010011;
ROM[5495] <= 32'b00000000000000010010001110000011;
ROM[5496] <= 32'b00000010011100011010000000100011;
ROM[5497] <= 32'b00000001111100000000001110010011;
ROM[5498] <= 32'b00000000011100010010000000100011;
ROM[5499] <= 32'b00000000010000010000000100010011;
ROM[5500] <= 32'b00000000000000011010001110000011;
ROM[5501] <= 32'b00000000011100010010000000100011;
ROM[5502] <= 32'b00000000010000010000000100010011;
ROM[5503] <= 32'b11111111110000010000000100010011;
ROM[5504] <= 32'b00000000000000010010001110000011;
ROM[5505] <= 32'b11111111110000010000000100010011;
ROM[5506] <= 32'b00000000000000010010010000000011;
ROM[5507] <= 32'b01000000011101000000001110110011;
ROM[5508] <= 32'b00000000011100010010000000100011;
ROM[5509] <= 32'b00000000010000010000000100010011;
ROM[5510] <= 32'b11111111110000010000000100010011;
ROM[5511] <= 32'b00000000000000010010001110000011;
ROM[5512] <= 32'b00000000011100011010111000100011;
ROM[5513] <= 32'b00000000001000000000001110010011;
ROM[5514] <= 32'b00000000011100010010000000100011;
ROM[5515] <= 32'b00000000010000010000000100010011;
ROM[5516] <= 32'b00000001110000011010001110000011;
ROM[5517] <= 32'b00000000011100010010000000100011;
ROM[5518] <= 32'b00000000010000010000000100010011;
ROM[5519] <= 32'b00000000000000000101001110110111;
ROM[5520] <= 32'b01101000100000111000001110010011;
ROM[5521] <= 32'b00000000111000111000001110110011;
ROM[5522] <= 32'b00000000011100010010000000100011;
ROM[5523] <= 32'b00000000010000010000000100010011;
ROM[5524] <= 32'b00000000001100010010000000100011;
ROM[5525] <= 32'b00000000010000010000000100010011;
ROM[5526] <= 32'b00000000010000010010000000100011;
ROM[5527] <= 32'b00000000010000010000000100010011;
ROM[5528] <= 32'b00000000010100010010000000100011;
ROM[5529] <= 32'b00000000010000010000000100010011;
ROM[5530] <= 32'b00000000011000010010000000100011;
ROM[5531] <= 32'b00000000010000010000000100010011;
ROM[5532] <= 32'b00000001010000000000001110010011;
ROM[5533] <= 32'b00000000100000111000001110010011;
ROM[5534] <= 32'b01000000011100010000001110110011;
ROM[5535] <= 32'b00000000011100000000001000110011;
ROM[5536] <= 32'b00000000001000000000000110110011;
ROM[5537] <= 32'b11111101000011111111000011101111;
ROM[5538] <= 32'b11111111110000010000000100010011;
ROM[5539] <= 32'b00000000000000010010001110000011;
ROM[5540] <= 32'b00000010011100011010001000100011;
ROM[5541] <= 32'b00000010000000011010001110000011;
ROM[5542] <= 32'b00000000011100010010000000100011;
ROM[5543] <= 32'b00000000010000010000000100010011;
ROM[5544] <= 32'b00000010010000011010001110000011;
ROM[5545] <= 32'b00000000011100010010000000100011;
ROM[5546] <= 32'b00000000010000010000000100010011;
ROM[5547] <= 32'b00000000000000000101001110110111;
ROM[5548] <= 32'b01101111100000111000001110010011;
ROM[5549] <= 32'b00000000111000111000001110110011;
ROM[5550] <= 32'b00000000011100010010000000100011;
ROM[5551] <= 32'b00000000010000010000000100010011;
ROM[5552] <= 32'b00000000001100010010000000100011;
ROM[5553] <= 32'b00000000010000010000000100010011;
ROM[5554] <= 32'b00000000010000010010000000100011;
ROM[5555] <= 32'b00000000010000010000000100010011;
ROM[5556] <= 32'b00000000010100010010000000100011;
ROM[5557] <= 32'b00000000010000010000000100010011;
ROM[5558] <= 32'b00000000011000010010000000100011;
ROM[5559] <= 32'b00000000010000010000000100010011;
ROM[5560] <= 32'b00000001010000000000001110010011;
ROM[5561] <= 32'b00000000100000111000001110010011;
ROM[5562] <= 32'b01000000011100010000001110110011;
ROM[5563] <= 32'b00000000011100000000001000110011;
ROM[5564] <= 32'b00000000001000000000000110110011;
ROM[5565] <= 32'b10111101100111111100000011101111;
ROM[5566] <= 32'b11111111110000010000000100010011;
ROM[5567] <= 32'b00000000000000010010001110000011;
ROM[5568] <= 32'b00000010011100011010010000100011;
ROM[5569] <= 32'b00000010100000011010001110000011;
ROM[5570] <= 32'b00000000011100010010000000100011;
ROM[5571] <= 32'b00000000010000010000000100010011;
ROM[5572] <= 32'b00000000000100000000001110010011;
ROM[5573] <= 32'b00000000011100010010000000100011;
ROM[5574] <= 32'b00000000010000010000000100010011;
ROM[5575] <= 32'b11111111110000010000000100010011;
ROM[5576] <= 32'b00000000000000010010001110000011;
ROM[5577] <= 32'b11111111110000010000000100010011;
ROM[5578] <= 32'b00000000000000010010010000000011;
ROM[5579] <= 32'b00000000011101000111001110110011;
ROM[5580] <= 32'b00000000011100010010000000100011;
ROM[5581] <= 32'b00000000010000010000000100010011;
ROM[5582] <= 32'b11111111110000010000000100010011;
ROM[5583] <= 32'b00000000000000010010001110000011;
ROM[5584] <= 32'b00000010011100011010011000100011;
ROM[5585] <= 32'b00000010110000011010001110000011;
ROM[5586] <= 32'b00000000011100010010000000100011;
ROM[5587] <= 32'b00000000010000010000000100010011;
ROM[5588] <= 32'b00000000000100000000001110010011;
ROM[5589] <= 32'b00000000011100010010000000100011;
ROM[5590] <= 32'b00000000010000010000000100010011;
ROM[5591] <= 32'b11111111110000010000000100010011;
ROM[5592] <= 32'b00000000000000010010001110000011;
ROM[5593] <= 32'b11111111110000010000000100010011;
ROM[5594] <= 32'b00000000000000010010010000000011;
ROM[5595] <= 32'b00000000011101000010010010110011;
ROM[5596] <= 32'b00000000100000111010010100110011;
ROM[5597] <= 32'b00000000101001001000001110110011;
ROM[5598] <= 32'b00000000000100111000001110010011;
ROM[5599] <= 32'b00000000000100111111001110010011;
ROM[5600] <= 32'b00000000011100010010000000100011;
ROM[5601] <= 32'b00000000010000010000000100010011;
ROM[5602] <= 32'b11111111110000010000000100010011;
ROM[5603] <= 32'b00000000000000010010001110000011;
ROM[5604] <= 32'b00000000000000111000101001100011;
ROM[5605] <= 32'b00000000000000000111001110110111;
ROM[5606] <= 32'b11111000100000111000001110010011;
ROM[5607] <= 32'b00000000111000111000001110110011;
ROM[5608] <= 32'b00000000000000111000000011100111;
ROM[5609] <= 32'b00000011000100000001000011101111;
ROM[5610] <= 32'b00000010000000011010001110000011;
ROM[5611] <= 32'b00000000011100010010000000100011;
ROM[5612] <= 32'b00000000010000010000000100010011;
ROM[5613] <= 32'b00000010010000011010001110000011;
ROM[5614] <= 32'b00000000011100010010000000100011;
ROM[5615] <= 32'b00000000010000010000000100010011;
ROM[5616] <= 32'b11111111110000010000000100010011;
ROM[5617] <= 32'b00000000000000010010001110000011;
ROM[5618] <= 32'b11111111110000010000000100010011;
ROM[5619] <= 32'b00000000000000010010010000000011;
ROM[5620] <= 32'b01000000011101000000001110110011;
ROM[5621] <= 32'b00000000011100010010000000100011;
ROM[5622] <= 32'b00000000010000010000000100010011;
ROM[5623] <= 32'b11111111110000010000000100010011;
ROM[5624] <= 32'b00000000000000010010001110000011;
ROM[5625] <= 32'b00000010011100011010000000100011;
ROM[5626] <= 32'b00000001110100000001000011101111;
ROM[5627] <= 32'b00000000011000000000001110010011;
ROM[5628] <= 32'b00000000011100010010000000100011;
ROM[5629] <= 32'b00000000010000010000000100010011;
ROM[5630] <= 32'b00000000110000011010001110000011;
ROM[5631] <= 32'b00000000011100010010000000100011;
ROM[5632] <= 32'b00000000010000010000000100010011;
ROM[5633] <= 32'b11111111110000010000000100010011;
ROM[5634] <= 32'b00000000000000010010001110000011;
ROM[5635] <= 32'b11111111110000010000000100010011;
ROM[5636] <= 32'b00000000000000010010010000000011;
ROM[5637] <= 32'b01000000011101000000001110110011;
ROM[5638] <= 32'b00000000011100010010000000100011;
ROM[5639] <= 32'b00000000010000010000000100010011;
ROM[5640] <= 32'b11111111110000010000000100010011;
ROM[5641] <= 32'b00000000000000010010001110000011;
ROM[5642] <= 32'b00000010011100011010100000100011;
ROM[5643] <= 32'b00000000001000000000001110010011;
ROM[5644] <= 32'b00000000011100010010000000100011;
ROM[5645] <= 32'b00000000010000010000000100010011;
ROM[5646] <= 32'b00000011000000011010001110000011;
ROM[5647] <= 32'b00000000011100010010000000100011;
ROM[5648] <= 32'b00000000010000010000000100010011;
ROM[5649] <= 32'b00000000000000000110001110110111;
ROM[5650] <= 32'b10001001000000111000001110010011;
ROM[5651] <= 32'b00000000111000111000001110110011;
ROM[5652] <= 32'b00000000011100010010000000100011;
ROM[5653] <= 32'b00000000010000010000000100010011;
ROM[5654] <= 32'b00000000001100010010000000100011;
ROM[5655] <= 32'b00000000010000010000000100010011;
ROM[5656] <= 32'b00000000010000010010000000100011;
ROM[5657] <= 32'b00000000010000010000000100010011;
ROM[5658] <= 32'b00000000010100010010000000100011;
ROM[5659] <= 32'b00000000010000010000000100010011;
ROM[5660] <= 32'b00000000011000010010000000100011;
ROM[5661] <= 32'b00000000010000010000000100010011;
ROM[5662] <= 32'b00000001010000000000001110010011;
ROM[5663] <= 32'b00000000100000111000001110010011;
ROM[5664] <= 32'b01000000011100010000001110110011;
ROM[5665] <= 32'b00000000011100000000001000110011;
ROM[5666] <= 32'b00000000001000000000000110110011;
ROM[5667] <= 32'b11011100100011111111000011101111;
ROM[5668] <= 32'b11111111110000010000000100010011;
ROM[5669] <= 32'b00000000000000010010001110000011;
ROM[5670] <= 32'b00000010011100011010101000100011;
ROM[5671] <= 32'b00000001100000011010001110000011;
ROM[5672] <= 32'b00000000011100010010000000100011;
ROM[5673] <= 32'b00000000010000010000000100010011;
ROM[5674] <= 32'b00000011010000011010001110000011;
ROM[5675] <= 32'b00000000011100010010000000100011;
ROM[5676] <= 32'b00000000010000010000000100010011;
ROM[5677] <= 32'b00000000000000000110001110110111;
ROM[5678] <= 32'b10010000000000111000001110010011;
ROM[5679] <= 32'b00000000111000111000001110110011;
ROM[5680] <= 32'b00000000011100010010000000100011;
ROM[5681] <= 32'b00000000010000010000000100010011;
ROM[5682] <= 32'b00000000001100010010000000100011;
ROM[5683] <= 32'b00000000010000010000000100010011;
ROM[5684] <= 32'b00000000010000010010000000100011;
ROM[5685] <= 32'b00000000010000010000000100010011;
ROM[5686] <= 32'b00000000010100010010000000100011;
ROM[5687] <= 32'b00000000010000010000000100010011;
ROM[5688] <= 32'b00000000011000010010000000100011;
ROM[5689] <= 32'b00000000010000010000000100010011;
ROM[5690] <= 32'b00000001010000000000001110010011;
ROM[5691] <= 32'b00000000100000111000001110010011;
ROM[5692] <= 32'b01000000011100010000001110110011;
ROM[5693] <= 32'b00000000011100000000001000110011;
ROM[5694] <= 32'b00000000001000000000000110110011;
ROM[5695] <= 32'b10011101000111111100000011101111;
ROM[5696] <= 32'b11111111110000010000000100010011;
ROM[5697] <= 32'b00000000000000010010001110000011;
ROM[5698] <= 32'b00000010011100011010110000100011;
ROM[5699] <= 32'b00000011100000011010001110000011;
ROM[5700] <= 32'b00000000011100010010000000100011;
ROM[5701] <= 32'b00000000010000010000000100010011;
ROM[5702] <= 32'b00000000000100000000001110010011;
ROM[5703] <= 32'b00000000011100010010000000100011;
ROM[5704] <= 32'b00000000010000010000000100010011;
ROM[5705] <= 32'b11111111110000010000000100010011;
ROM[5706] <= 32'b00000000000000010010001110000011;
ROM[5707] <= 32'b11111111110000010000000100010011;
ROM[5708] <= 32'b00000000000000010010010000000011;
ROM[5709] <= 32'b00000000011101000111001110110011;
ROM[5710] <= 32'b00000000011100010010000000100011;
ROM[5711] <= 32'b00000000010000010000000100010011;
ROM[5712] <= 32'b11111111110000010000000100010011;
ROM[5713] <= 32'b00000000000000010010001110000011;
ROM[5714] <= 32'b00000010011100011010011000100011;
ROM[5715] <= 32'b00000010110000011010001110000011;
ROM[5716] <= 32'b00000000011100010010000000100011;
ROM[5717] <= 32'b00000000010000010000000100010011;
ROM[5718] <= 32'b00000000000100000000001110010011;
ROM[5719] <= 32'b00000000011100010010000000100011;
ROM[5720] <= 32'b00000000010000010000000100010011;
ROM[5721] <= 32'b11111111110000010000000100010011;
ROM[5722] <= 32'b00000000000000010010001110000011;
ROM[5723] <= 32'b11111111110000010000000100010011;
ROM[5724] <= 32'b00000000000000010010010000000011;
ROM[5725] <= 32'b00000000011101000010010010110011;
ROM[5726] <= 32'b00000000100000111010010100110011;
ROM[5727] <= 32'b00000000101001001000001110110011;
ROM[5728] <= 32'b00000000000100111000001110010011;
ROM[5729] <= 32'b00000000000100111111001110010011;
ROM[5730] <= 32'b00000000011100010010000000100011;
ROM[5731] <= 32'b00000000010000010000000100010011;
ROM[5732] <= 32'b11111111110000010000000100010011;
ROM[5733] <= 32'b00000000000000010010001110000011;
ROM[5734] <= 32'b00000000000000111000101001100011;
ROM[5735] <= 32'b00000000000000000111001110110111;
ROM[5736] <= 32'b00101100100000111000001110010011;
ROM[5737] <= 32'b00000000111000111000001110110011;
ROM[5738] <= 32'b00000000000000111000000011100111;
ROM[5739] <= 32'b00010111100100000001000011101111;
ROM[5740] <= 32'b00000010000000011010001110000011;
ROM[5741] <= 32'b00000000011100010010000000100011;
ROM[5742] <= 32'b00000000010000010000000100010011;
ROM[5743] <= 32'b00000010010000011010001110000011;
ROM[5744] <= 32'b00000000011100010010000000100011;
ROM[5745] <= 32'b00000000010000010000000100010011;
ROM[5746] <= 32'b11111111110000010000000100010011;
ROM[5747] <= 32'b00000000000000010010001110000011;
ROM[5748] <= 32'b11111111110000010000000100010011;
ROM[5749] <= 32'b00000000000000010010010000000011;
ROM[5750] <= 32'b00000000011101000000001110110011;
ROM[5751] <= 32'b00000000011100010010000000100011;
ROM[5752] <= 32'b00000000010000010000000100010011;
ROM[5753] <= 32'b11111111110000010000000100010011;
ROM[5754] <= 32'b00000000000000010010001110000011;
ROM[5755] <= 32'b00000010011100011010000000100011;
ROM[5756] <= 32'b00010111100100000001000011101111;
ROM[5757] <= 32'b00000100000000011010001110000011;
ROM[5758] <= 32'b00000000011100010010000000100011;
ROM[5759] <= 32'b00000000010000010000000100010011;
ROM[5760] <= 32'b00000111010001101010001110000011;
ROM[5761] <= 32'b00000000011100010010000000100011;
ROM[5762] <= 32'b00000000010000010000000100010011;
ROM[5763] <= 32'b11111111110000010000000100010011;
ROM[5764] <= 32'b00000000000000010010001110000011;
ROM[5765] <= 32'b11111111110000010000000100010011;
ROM[5766] <= 32'b00000000000000010010010000000011;
ROM[5767] <= 32'b00000000011101000000001110110011;
ROM[5768] <= 32'b00000000011100010010000000100011;
ROM[5769] <= 32'b00000000010000010000000100010011;
ROM[5770] <= 32'b00000010000000011010001110000011;
ROM[5771] <= 32'b00000000011100010010000000100011;
ROM[5772] <= 32'b00000000010000010000000100010011;
ROM[5773] <= 32'b11111111110000010000000100010011;
ROM[5774] <= 32'b00000000000000010010001110000011;
ROM[5775] <= 32'b00000000011101100010000000100011;
ROM[5776] <= 32'b11111111110000010000000100010011;
ROM[5777] <= 32'b00000000000000010010001110000011;
ROM[5778] <= 32'b00000000000000111000001100010011;
ROM[5779] <= 32'b00000000000001100010001110000011;
ROM[5780] <= 32'b00000000011100010010000000100011;
ROM[5781] <= 32'b00000000010000010000000100010011;
ROM[5782] <= 32'b11111111110000010000000100010011;
ROM[5783] <= 32'b00000000000000010010001110000011;
ROM[5784] <= 32'b00000000110100110000010000110011;
ROM[5785] <= 32'b00000000011101000010000000100011;
ROM[5786] <= 32'b10010011110111111111000011101111;
ROM[5787] <= 32'b00000000000000011010001110000011;
ROM[5788] <= 32'b00000000011100010010000000100011;
ROM[5789] <= 32'b00000000010000010000000100010011;
ROM[5790] <= 32'b00000000000100000000001110010011;
ROM[5791] <= 32'b00000000011100010010000000100011;
ROM[5792] <= 32'b00000000010000010000000100010011;
ROM[5793] <= 32'b11111111110000010000000100010011;
ROM[5794] <= 32'b00000000000000010010001110000011;
ROM[5795] <= 32'b11111111110000010000000100010011;
ROM[5796] <= 32'b00000000000000010010010000000011;
ROM[5797] <= 32'b00000000011101000000001110110011;
ROM[5798] <= 32'b00000000011100010010000000100011;
ROM[5799] <= 32'b00000000010000010000000100010011;
ROM[5800] <= 32'b11111111110000010000000100010011;
ROM[5801] <= 32'b00000000000000010010001110000011;
ROM[5802] <= 32'b00000000011100011010000000100011;
ROM[5803] <= 32'b00000000110000011010001110000011;
ROM[5804] <= 32'b00000000011100010010000000100011;
ROM[5805] <= 32'b00000000010000010000000100010011;
ROM[5806] <= 32'b00000000000100000000001110010011;
ROM[5807] <= 32'b00000000011100010010000000100011;
ROM[5808] <= 32'b00000000010000010000000100010011;
ROM[5809] <= 32'b11111111110000010000000100010011;
ROM[5810] <= 32'b00000000000000010010001110000011;
ROM[5811] <= 32'b11111111110000010000000100010011;
ROM[5812] <= 32'b00000000000000010010010000000011;
ROM[5813] <= 32'b00000000011101000000001110110011;
ROM[5814] <= 32'b00000000011100010010000000100011;
ROM[5815] <= 32'b00000000010000010000000100010011;
ROM[5816] <= 32'b11111111110000010000000100010011;
ROM[5817] <= 32'b00000000000000010010001110000011;
ROM[5818] <= 32'b00000000011100011010011000100011;
ROM[5819] <= 32'b00000000000000011010001110000011;
ROM[5820] <= 32'b00000000011100010010000000100011;
ROM[5821] <= 32'b00000000010000010000000100010011;
ROM[5822] <= 32'b00000010000000000000001110010011;
ROM[5823] <= 32'b00000000011100010010000000100011;
ROM[5824] <= 32'b00000000010000010000000100010011;
ROM[5825] <= 32'b11111111110000010000000100010011;
ROM[5826] <= 32'b00000000000000010010001110000011;
ROM[5827] <= 32'b11111111110000010000000100010011;
ROM[5828] <= 32'b00000000000000010010010000000011;
ROM[5829] <= 32'b00000000011101000010010010110011;
ROM[5830] <= 32'b00000000100000111010010100110011;
ROM[5831] <= 32'b00000000101001001000001110110011;
ROM[5832] <= 32'b00000000000100111000001110010011;
ROM[5833] <= 32'b00000000000100111111001110010011;
ROM[5834] <= 32'b00000000011100010010000000100011;
ROM[5835] <= 32'b00000000010000010000000100010011;
ROM[5836] <= 32'b11111111110000010000000100010011;
ROM[5837] <= 32'b00000000000000010010001110000011;
ROM[5838] <= 32'b00000000000000111000101001100011;
ROM[5839] <= 32'b00000000000000000111001110110111;
ROM[5840] <= 32'b01011011010000111000001110010011;
ROM[5841] <= 32'b00000000111000111000001110110011;
ROM[5842] <= 32'b00000000000000111000000011100111;
ROM[5843] <= 32'b00110000010100000001000011101111;
ROM[5844] <= 32'b00000000000000000000001110010011;
ROM[5845] <= 32'b00000000011100010010000000100011;
ROM[5846] <= 32'b00000000010000010000000100010011;
ROM[5847] <= 32'b11111111110000010000000100010011;
ROM[5848] <= 32'b00000000000000010010001110000011;
ROM[5849] <= 32'b00000000011100011010000000100011;
ROM[5850] <= 32'b00000000100000011010001110000011;
ROM[5851] <= 32'b00000000011100010010000000100011;
ROM[5852] <= 32'b00000000010000010000000100010011;
ROM[5853] <= 32'b00000000000100000000001110010011;
ROM[5854] <= 32'b00000000011100010010000000100011;
ROM[5855] <= 32'b00000000010000010000000100010011;
ROM[5856] <= 32'b11111111110000010000000100010011;
ROM[5857] <= 32'b00000000000000010010001110000011;
ROM[5858] <= 32'b11111111110000010000000100010011;
ROM[5859] <= 32'b00000000000000010010010000000011;
ROM[5860] <= 32'b00000000011101000000001110110011;
ROM[5861] <= 32'b00000000011100010010000000100011;
ROM[5862] <= 32'b00000000010000010000000100010011;
ROM[5863] <= 32'b11111111110000010000000100010011;
ROM[5864] <= 32'b00000000000000010010001110000011;
ROM[5865] <= 32'b00000000011100011010010000100011;
ROM[5866] <= 32'b00101010100100000001000011101111;
ROM[5867] <= 32'b00100010010000000010000011101111;
ROM[5868] <= 32'b00001000000001101010001110000011;
ROM[5869] <= 32'b00000000011100010010000000100011;
ROM[5870] <= 32'b00000000010000010000000100010011;
ROM[5871] <= 32'b00000010001100000000001110010011;
ROM[5872] <= 32'b00000000011100010010000000100011;
ROM[5873] <= 32'b00000000010000010000000100010011;
ROM[5874] <= 32'b11111111110000010000000100010011;
ROM[5875] <= 32'b00000000000000010010001110000011;
ROM[5876] <= 32'b11111111110000010000000100010011;
ROM[5877] <= 32'b00000000000000010010010000000011;
ROM[5878] <= 32'b00000000011101000010010010110011;
ROM[5879] <= 32'b00000000100000111010010100110011;
ROM[5880] <= 32'b00000000101001001000001110110011;
ROM[5881] <= 32'b00000000000100111000001110010011;
ROM[5882] <= 32'b00000000000100111111001110010011;
ROM[5883] <= 32'b00000000011100010010000000100011;
ROM[5884] <= 32'b00000000010000010000000100010011;
ROM[5885] <= 32'b11111111110000010000000100010011;
ROM[5886] <= 32'b00000000000000010010001110000011;
ROM[5887] <= 32'b00000000000000111000101001100011;
ROM[5888] <= 32'b00000000000000000111001110110111;
ROM[5889] <= 32'b01110111010000111000001110010011;
ROM[5890] <= 32'b00000000111000111000001110110011;
ROM[5891] <= 32'b00000000000000111000000011100111;
ROM[5892] <= 32'b01000010000100000001000011101111;
ROM[5893] <= 32'b00000000000000000000001110010011;
ROM[5894] <= 32'b00000000011100010010000000100011;
ROM[5895] <= 32'b00000000010000010000000100010011;
ROM[5896] <= 32'b11111111110000010000000100010011;
ROM[5897] <= 32'b00000000000000010010001110000011;
ROM[5898] <= 32'b00001000011101101010000000100011;
ROM[5899] <= 32'b00001000100001101010001110000011;
ROM[5900] <= 32'b00000000011100010010000000100011;
ROM[5901] <= 32'b00000000010000010000000100010011;
ROM[5902] <= 32'b00000000000100000000001110010011;
ROM[5903] <= 32'b00000000011100010010000000100011;
ROM[5904] <= 32'b00000000010000010000000100010011;
ROM[5905] <= 32'b11111111110000010000000100010011;
ROM[5906] <= 32'b00000000000000010010001110000011;
ROM[5907] <= 32'b11111111110000010000000100010011;
ROM[5908] <= 32'b00000000000000010010010000000011;
ROM[5909] <= 32'b00000000011101000000001110110011;
ROM[5910] <= 32'b00000000011100010010000000100011;
ROM[5911] <= 32'b00000000010000010000000100010011;
ROM[5912] <= 32'b11111111110000010000000100010011;
ROM[5913] <= 32'b00000000000000010010001110000011;
ROM[5914] <= 32'b00001000011101101010010000100011;
ROM[5915] <= 32'b01011101100100000001000011101111;
ROM[5916] <= 32'b00001000000001101010001110000011;
ROM[5917] <= 32'b00000000011100010010000000100011;
ROM[5918] <= 32'b00000000010000010000000100010011;
ROM[5919] <= 32'b00000000000100000000001110010011;
ROM[5920] <= 32'b00000000011100010010000000100011;
ROM[5921] <= 32'b00000000010000010000000100010011;
ROM[5922] <= 32'b11111111110000010000000100010011;
ROM[5923] <= 32'b00000000000000010010001110000011;
ROM[5924] <= 32'b11111111110000010000000100010011;
ROM[5925] <= 32'b00000000000000010010010000000011;
ROM[5926] <= 32'b00000000011101000000001110110011;
ROM[5927] <= 32'b00000000011100010010000000100011;
ROM[5928] <= 32'b00000000010000010000000100010011;
ROM[5929] <= 32'b11111111110000010000000100010011;
ROM[5930] <= 32'b00000000000000010010001110000011;
ROM[5931] <= 32'b00001000011101101010000000100011;
ROM[5932] <= 32'b00000000000000000000001110010011;
ROM[5933] <= 32'b00000000011100010010000000100011;
ROM[5934] <= 32'b00000000010000010000000100010011;
ROM[5935] <= 32'b00000001010000000000001110010011;
ROM[5936] <= 32'b01000000011100011000001110110011;
ROM[5937] <= 32'b00000000000000111010000010000011;
ROM[5938] <= 32'b11111111110000010000000100010011;
ROM[5939] <= 32'b00000000000000010010001110000011;
ROM[5940] <= 32'b00000000011100100010000000100011;
ROM[5941] <= 32'b00000000010000100000000100010011;
ROM[5942] <= 32'b00000001010000000000001110010011;
ROM[5943] <= 32'b01000000011100011000001110110011;
ROM[5944] <= 32'b00000000010000111010000110000011;
ROM[5945] <= 32'b00000000100000111010001000000011;
ROM[5946] <= 32'b00000000110000111010001010000011;
ROM[5947] <= 32'b00000001000000111010001100000011;
ROM[5948] <= 32'b00000000000000001000000011100111;
ROM[5949] <= 32'b00000000000000000000001110010011;
ROM[5950] <= 32'b00000000011100010010000000100011;
ROM[5951] <= 32'b00000000010000010000000100010011;
ROM[5952] <= 32'b11111111110000010000000100010011;
ROM[5953] <= 32'b00000000000000010010001110000011;
ROM[5954] <= 32'b00001000011101101010000000100011;
ROM[5955] <= 32'b00001000100001101010001110000011;
ROM[5956] <= 32'b00000000011100010010000000100011;
ROM[5957] <= 32'b00000000010000010000000100010011;
ROM[5958] <= 32'b00000000000100000000001110010011;
ROM[5959] <= 32'b00000000011100010010000000100011;
ROM[5960] <= 32'b00000000010000010000000100010011;
ROM[5961] <= 32'b11111111110000010000000100010011;
ROM[5962] <= 32'b00000000000000010010001110000011;
ROM[5963] <= 32'b11111111110000010000000100010011;
ROM[5964] <= 32'b00000000000000010010010000000011;
ROM[5965] <= 32'b00000000011101000000001110110011;
ROM[5966] <= 32'b00000000011100010010000000100011;
ROM[5967] <= 32'b00000000010000010000000100010011;
ROM[5968] <= 32'b11111111110000010000000100010011;
ROM[5969] <= 32'b00000000000000010010001110000011;
ROM[5970] <= 32'b00001000011101101010010000100011;
ROM[5971] <= 32'b00000000000000000000001110010011;
ROM[5972] <= 32'b00000000011100010010000000100011;
ROM[5973] <= 32'b00000000010000010000000100010011;
ROM[5974] <= 32'b00000001010000000000001110010011;
ROM[5975] <= 32'b01000000011100011000001110110011;
ROM[5976] <= 32'b00000000000000111010000010000011;
ROM[5977] <= 32'b11111111110000010000000100010011;
ROM[5978] <= 32'b00000000000000010010001110000011;
ROM[5979] <= 32'b00000000011100100010000000100011;
ROM[5980] <= 32'b00000000010000100000000100010011;
ROM[5981] <= 32'b00000001010000000000001110010011;
ROM[5982] <= 32'b01000000011100011000001110110011;
ROM[5983] <= 32'b00000000010000111010000110000011;
ROM[5984] <= 32'b00000000100000111010001000000011;
ROM[5985] <= 32'b00000000110000111010001010000011;
ROM[5986] <= 32'b00000001000000111010001100000011;
ROM[5987] <= 32'b00000000000000001000000011100111;
ROM[5988] <= 32'b00000000000000010010000000100011;
ROM[5989] <= 32'b00000000010000010000000100010011;
ROM[5990] <= 32'b00000000000000010010000000100011;
ROM[5991] <= 32'b00000000010000010000000100010011;
ROM[5992] <= 32'b00000000000000010010000000100011;
ROM[5993] <= 32'b00000000010000010000000100010011;
ROM[5994] <= 32'b00000000000000010010000000100011;
ROM[5995] <= 32'b00000000010000010000000100010011;
ROM[5996] <= 32'b00000000000000010010000000100011;
ROM[5997] <= 32'b00000000010000010000000100010011;
ROM[5998] <= 32'b00000000000000010010000000100011;
ROM[5999] <= 32'b00000000010000010000000100010011;
ROM[6000] <= 32'b00000000000000010010000000100011;
ROM[6001] <= 32'b00000000010000010000000100010011;
ROM[6002] <= 32'b00000000000000010010000000100011;
ROM[6003] <= 32'b00000000010000010000000100010011;
ROM[6004] <= 32'b00000000000000010010000000100011;
ROM[6005] <= 32'b00000000010000010000000100010011;
ROM[6006] <= 32'b00000000000000010010000000100011;
ROM[6007] <= 32'b00000000010000010000000100010011;
ROM[6008] <= 32'b00000000000000010010000000100011;
ROM[6009] <= 32'b00000000010000010000000100010011;
ROM[6010] <= 32'b00000000000000010010000000100011;
ROM[6011] <= 32'b00000000010000010000000100010011;
ROM[6012] <= 32'b00000000000000010010000000100011;
ROM[6013] <= 32'b00000000010000010000000100010011;
ROM[6014] <= 32'b00001000000001101010001110000011;
ROM[6015] <= 32'b00000000011100010010000000100011;
ROM[6016] <= 32'b00000000010000010000000100010011;
ROM[6017] <= 32'b00001000000001101010001110000011;
ROM[6018] <= 32'b00000000011100010010000000100011;
ROM[6019] <= 32'b00000000010000010000000100010011;
ROM[6020] <= 32'b11111111110000010000000100010011;
ROM[6021] <= 32'b00000000000000010010001110000011;
ROM[6022] <= 32'b11111111110000010000000100010011;
ROM[6023] <= 32'b00000000000000010010010000000011;
ROM[6024] <= 32'b00000000011101000000001110110011;
ROM[6025] <= 32'b00000000011100010010000000100011;
ROM[6026] <= 32'b00000000010000010000000100010011;
ROM[6027] <= 32'b00001000000001101010001110000011;
ROM[6028] <= 32'b00000000011100010010000000100011;
ROM[6029] <= 32'b00000000010000010000000100010011;
ROM[6030] <= 32'b11111111110000010000000100010011;
ROM[6031] <= 32'b00000000000000010010001110000011;
ROM[6032] <= 32'b11111111110000010000000100010011;
ROM[6033] <= 32'b00000000000000010010010000000011;
ROM[6034] <= 32'b00000000011101000000001110110011;
ROM[6035] <= 32'b00000000011100010010000000100011;
ROM[6036] <= 32'b00000000010000010000000100010011;
ROM[6037] <= 32'b00001000000001101010001110000011;
ROM[6038] <= 32'b00000000011100010010000000100011;
ROM[6039] <= 32'b00000000010000010000000100010011;
ROM[6040] <= 32'b11111111110000010000000100010011;
ROM[6041] <= 32'b00000000000000010010001110000011;
ROM[6042] <= 32'b11111111110000010000000100010011;
ROM[6043] <= 32'b00000000000000010010010000000011;
ROM[6044] <= 32'b00000000011101000000001110110011;
ROM[6045] <= 32'b00000000011100010010000000100011;
ROM[6046] <= 32'b00000000010000010000000100010011;
ROM[6047] <= 32'b11111111110000010000000100010011;
ROM[6048] <= 32'b00000000000000010010001110000011;
ROM[6049] <= 32'b00001000011101101010001000100011;
ROM[6050] <= 32'b00001000010001101010001110000011;
ROM[6051] <= 32'b00000000011100010010000000100011;
ROM[6052] <= 32'b00000000010000010000000100010011;
ROM[6053] <= 32'b00001000110001101010001110000011;
ROM[6054] <= 32'b00000000011100010010000000100011;
ROM[6055] <= 32'b00000000010000010000000100010011;
ROM[6056] <= 32'b11111111110000010000000100010011;
ROM[6057] <= 32'b00000000000000010010001110000011;
ROM[6058] <= 32'b11111111110000010000000100010011;
ROM[6059] <= 32'b00000000000000010010010000000011;
ROM[6060] <= 32'b00000000011101000000001110110011;
ROM[6061] <= 32'b00000000011100010010000000100011;
ROM[6062] <= 32'b00000000010000010000000100010011;
ROM[6063] <= 32'b11111111110000010000000100010011;
ROM[6064] <= 32'b00000000000000010010001110000011;
ROM[6065] <= 32'b00000000000000111000001100010011;
ROM[6066] <= 32'b00000000110100110000010000110011;
ROM[6067] <= 32'b00000000000001000010001110000011;
ROM[6068] <= 32'b00000000011100010010000000100011;
ROM[6069] <= 32'b00000000010000010000000100010011;
ROM[6070] <= 32'b11111111110000010000000100010011;
ROM[6071] <= 32'b00000000000000010010001110000011;
ROM[6072] <= 32'b00000000011100011010001000100011;
ROM[6073] <= 32'b00001000100001101010001110000011;
ROM[6074] <= 32'b00000000011100010010000000100011;
ROM[6075] <= 32'b00000000010000010000000100010011;
ROM[6076] <= 32'b00000110010000000000001110010011;
ROM[6077] <= 32'b00000000011100010010000000100011;
ROM[6078] <= 32'b00000000010000010000000100010011;
ROM[6079] <= 32'b00000000000000000110001110110111;
ROM[6080] <= 32'b11110100100000111000001110010011;
ROM[6081] <= 32'b00000000111000111000001110110011;
ROM[6082] <= 32'b00000000011100010010000000100011;
ROM[6083] <= 32'b00000000010000010000000100010011;
ROM[6084] <= 32'b00000000001100010010000000100011;
ROM[6085] <= 32'b00000000010000010000000100010011;
ROM[6086] <= 32'b00000000010000010010000000100011;
ROM[6087] <= 32'b00000000010000010000000100010011;
ROM[6088] <= 32'b00000000010100010010000000100011;
ROM[6089] <= 32'b00000000010000010000000100010011;
ROM[6090] <= 32'b00000000011000010010000000100011;
ROM[6091] <= 32'b00000000010000010000000100010011;
ROM[6092] <= 32'b00000001010000000000001110010011;
ROM[6093] <= 32'b00000000100000111000001110010011;
ROM[6094] <= 32'b01000000011100010000001110110011;
ROM[6095] <= 32'b00000000011100000000001000110011;
ROM[6096] <= 32'b00000000001000000000000110110011;
ROM[6097] <= 32'b10000000010011111100000011101111;
ROM[6098] <= 32'b00000000010000011010001110000011;
ROM[6099] <= 32'b00000000011100010010000000100011;
ROM[6100] <= 32'b00000000010000010000000100010011;
ROM[6101] <= 32'b00000010000000000000001110010011;
ROM[6102] <= 32'b00000000011100010010000000100011;
ROM[6103] <= 32'b00000000010000010000000100010011;
ROM[6104] <= 32'b00000000000000000110001110110111;
ROM[6105] <= 32'b11111010110000111000001110010011;
ROM[6106] <= 32'b00000000111000111000001110110011;
ROM[6107] <= 32'b00000000011100010010000000100011;
ROM[6108] <= 32'b00000000010000010000000100010011;
ROM[6109] <= 32'b00000000001100010010000000100011;
ROM[6110] <= 32'b00000000010000010000000100010011;
ROM[6111] <= 32'b00000000010000010010000000100011;
ROM[6112] <= 32'b00000000010000010000000100010011;
ROM[6113] <= 32'b00000000010100010010000000100011;
ROM[6114] <= 32'b00000000010000010000000100010011;
ROM[6115] <= 32'b00000000011000010010000000100011;
ROM[6116] <= 32'b00000000010000010000000100010011;
ROM[6117] <= 32'b00000001010000000000001110010011;
ROM[6118] <= 32'b00000000100000111000001110010011;
ROM[6119] <= 32'b01000000011100010000001110110011;
ROM[6120] <= 32'b00000000011100000000001000110011;
ROM[6121] <= 32'b00000000001000000000000110110011;
ROM[6122] <= 32'b10110010010011111100000011101111;
ROM[6123] <= 32'b11111111110000010000000100010011;
ROM[6124] <= 32'b00000000000000010010001110000011;
ROM[6125] <= 32'b11111111110000010000000100010011;
ROM[6126] <= 32'b00000000000000010010010000000011;
ROM[6127] <= 32'b00000000011101000000001110110011;
ROM[6128] <= 32'b00000000011100010010000000100011;
ROM[6129] <= 32'b00000000010000010000000100010011;
ROM[6130] <= 32'b11111111110000010000000100010011;
ROM[6131] <= 32'b00000000000000010010001110000011;
ROM[6132] <= 32'b00000000011100011010010000100011;
ROM[6133] <= 32'b00000000010000011010001110000011;
ROM[6134] <= 32'b00000000011100010010000000100011;
ROM[6135] <= 32'b00000000010000010000000100010011;
ROM[6136] <= 32'b00000010000000000000001110010011;
ROM[6137] <= 32'b00000000011100010010000000100011;
ROM[6138] <= 32'b00000000010000010000000100010011;
ROM[6139] <= 32'b00000000000000000110001110110111;
ROM[6140] <= 32'b00000011100000111000001110010011;
ROM[6141] <= 32'b00000000111000111000001110110011;
ROM[6142] <= 32'b00000000011100010010000000100011;
ROM[6143] <= 32'b00000000010000010000000100010011;
ROM[6144] <= 32'b00000000001100010010000000100011;
ROM[6145] <= 32'b00000000010000010000000100010011;
ROM[6146] <= 32'b00000000010000010010000000100011;
ROM[6147] <= 32'b00000000010000010000000100010011;
ROM[6148] <= 32'b00000000010100010010000000100011;
ROM[6149] <= 32'b00000000010000010000000100010011;
ROM[6150] <= 32'b00000000011000010010000000100011;
ROM[6151] <= 32'b00000000010000010000000100010011;
ROM[6152] <= 32'b00000001010000000000001110010011;
ROM[6153] <= 32'b00000000100000111000001110010011;
ROM[6154] <= 32'b01000000011100010000001110110011;
ROM[6155] <= 32'b00000000011100000000001000110011;
ROM[6156] <= 32'b00000000001000000000000110110011;
ROM[6157] <= 32'b10001101110111111100000011101111;
ROM[6158] <= 32'b11111111110000010000000100010011;
ROM[6159] <= 32'b00000000000000010010001110000011;
ROM[6160] <= 32'b00000000011100011010000000100011;
ROM[6161] <= 32'b00000000000000000000001110010011;
ROM[6162] <= 32'b00000000011100010010000000100011;
ROM[6163] <= 32'b00000000010000010000000100010011;
ROM[6164] <= 32'b11111111110000010000000100010011;
ROM[6165] <= 32'b00000000000000010010001110000011;
ROM[6166] <= 32'b00000000011100011010011000100011;
ROM[6167] <= 32'b00001000000001101010001110000011;
ROM[6168] <= 32'b00000000011100010010000000100011;
ROM[6169] <= 32'b00000000010000010000000100010011;
ROM[6170] <= 32'b00000000000000000000001110010011;
ROM[6171] <= 32'b00000000011100010010000000100011;
ROM[6172] <= 32'b00000000010000010000000100010011;
ROM[6173] <= 32'b11111111110000010000000100010011;
ROM[6174] <= 32'b00000000000000010010001110000011;
ROM[6175] <= 32'b11111111110000010000000100010011;
ROM[6176] <= 32'b00000000000000010010010000000011;
ROM[6177] <= 32'b00000000011101000010010010110011;
ROM[6178] <= 32'b00000000100000111010010100110011;
ROM[6179] <= 32'b00000000101001001000001110110011;
ROM[6180] <= 32'b00000000000100111000001110010011;
ROM[6181] <= 32'b00000000000100111111001110010011;
ROM[6182] <= 32'b00000000011100010010000000100011;
ROM[6183] <= 32'b00000000010000010000000100010011;
ROM[6184] <= 32'b11111111110000010000000100010011;
ROM[6185] <= 32'b00000000000000010010001110000011;
ROM[6186] <= 32'b00000000000000111000101001100011;
ROM[6187] <= 32'b00000000000000000110001110110111;
ROM[6188] <= 32'b00001100000000111000001110010011;
ROM[6189] <= 32'b00000000111000111000001110110011;
ROM[6190] <= 32'b00000000000000111000000011100111;
ROM[6191] <= 32'b00001011100000000000000011101111;
ROM[6192] <= 32'b00001000100001101010001110000011;
ROM[6193] <= 32'b00000000011100010010000000100011;
ROM[6194] <= 32'b00000000010000010000000100010011;
ROM[6195] <= 32'b00000000000000000000001110010011;
ROM[6196] <= 32'b00000000011100010010000000100011;
ROM[6197] <= 32'b00000000010000010000000100010011;
ROM[6198] <= 32'b11111111110000010000000100010011;
ROM[6199] <= 32'b00000000000000010010001110000011;
ROM[6200] <= 32'b11111111110000010000000100010011;
ROM[6201] <= 32'b00000000000000010010010000000011;
ROM[6202] <= 32'b00000000100000111010001110110011;
ROM[6203] <= 32'b00000000011100010010000000100011;
ROM[6204] <= 32'b00000000010000010000000100010011;
ROM[6205] <= 32'b11111111110000010000000100010011;
ROM[6206] <= 32'b00000000000000010010001110000011;
ROM[6207] <= 32'b00000000000000111000101001100011;
ROM[6208] <= 32'b00000000000000000110001110110111;
ROM[6209] <= 32'b00010001010000111000001110010011;
ROM[6210] <= 32'b00000000111000111000001110110011;
ROM[6211] <= 32'b00000000000000111000000011100111;
ROM[6212] <= 32'b00000110000000000000000011101111;
ROM[6213] <= 32'b00001000100001101010001110000011;
ROM[6214] <= 32'b00000000011100010010000000100011;
ROM[6215] <= 32'b00000000010000010000000100010011;
ROM[6216] <= 32'b00000000000100000000001110010011;
ROM[6217] <= 32'b00000000011100010010000000100011;
ROM[6218] <= 32'b00000000010000010000000100010011;
ROM[6219] <= 32'b11111111110000010000000100010011;
ROM[6220] <= 32'b00000000000000010010001110000011;
ROM[6221] <= 32'b11111111110000010000000100010011;
ROM[6222] <= 32'b00000000000000010010010000000011;
ROM[6223] <= 32'b01000000011101000000001110110011;
ROM[6224] <= 32'b00000000011100010010000000100011;
ROM[6225] <= 32'b00000000010000010000000100010011;
ROM[6226] <= 32'b11111111110000010000000100010011;
ROM[6227] <= 32'b00000000000000010010001110000011;
ROM[6228] <= 32'b00001000011101101010010000100011;
ROM[6229] <= 32'b00000010001100000000001110010011;
ROM[6230] <= 32'b00000000011100010010000000100011;
ROM[6231] <= 32'b00000000010000010000000100010011;
ROM[6232] <= 32'b11111111110000010000000100010011;
ROM[6233] <= 32'b00000000000000010010001110000011;
ROM[6234] <= 32'b00001000011101101010000000100011;
ROM[6235] <= 32'b00000000010000000000000011101111;
ROM[6236] <= 32'b00000100010000000000000011101111;
ROM[6237] <= 32'b00001000000001101010001110000011;
ROM[6238] <= 32'b00000000011100010010000000100011;
ROM[6239] <= 32'b00000000010000010000000100010011;
ROM[6240] <= 32'b00000000000100000000001110010011;
ROM[6241] <= 32'b00000000011100010010000000100011;
ROM[6242] <= 32'b00000000010000010000000100010011;
ROM[6243] <= 32'b11111111110000010000000100010011;
ROM[6244] <= 32'b00000000000000010010001110000011;
ROM[6245] <= 32'b11111111110000010000000100010011;
ROM[6246] <= 32'b00000000000000010010010000000011;
ROM[6247] <= 32'b01000000011101000000001110110011;
ROM[6248] <= 32'b00000000011100010010000000100011;
ROM[6249] <= 32'b00000000010000010000000100010011;
ROM[6250] <= 32'b11111111110000010000000100010011;
ROM[6251] <= 32'b00000000000000010010001110000011;
ROM[6252] <= 32'b00001000011101101010000000100011;
ROM[6253] <= 32'b00000000110000011010001110000011;
ROM[6254] <= 32'b00000000011100010010000000100011;
ROM[6255] <= 32'b00000000010000010000000100010011;
ROM[6256] <= 32'b00000000011100000000001110010011;
ROM[6257] <= 32'b00000000011100010010000000100011;
ROM[6258] <= 32'b00000000010000010000000100010011;
ROM[6259] <= 32'b11111111110000010000000100010011;
ROM[6260] <= 32'b00000000000000010010001110000011;
ROM[6261] <= 32'b11111111110000010000000100010011;
ROM[6262] <= 32'b00000000000000010010010000000011;
ROM[6263] <= 32'b00000000011101000010001110110011;
ROM[6264] <= 32'b00000000011100010010000000100011;
ROM[6265] <= 32'b00000000010000010000000100010011;
ROM[6266] <= 32'b11111111110000010000000100010011;
ROM[6267] <= 32'b00000000000000010010001110000011;
ROM[6268] <= 32'b01000000011100000000001110110011;
ROM[6269] <= 32'b00000000000100111000001110010011;
ROM[6270] <= 32'b00000000011100010010000000100011;
ROM[6271] <= 32'b00000000010000010000000100010011;
ROM[6272] <= 32'b11111111110000010000000100010011;
ROM[6273] <= 32'b00000000000000010010001110000011;
ROM[6274] <= 32'b00000000000000111000101001100011;
ROM[6275] <= 32'b00000000000000000110001110110111;
ROM[6276] <= 32'b01111101110000111000001110010011;
ROM[6277] <= 32'b00000000111000111000001110110011;
ROM[6278] <= 32'b00000000000000111000000011100111;
ROM[6279] <= 32'b00000000000000000000001110010011;
ROM[6280] <= 32'b00000000011100010010000000100011;
ROM[6281] <= 32'b00000000010000010000000100010011;
ROM[6282] <= 32'b11111111110000010000000100010011;
ROM[6283] <= 32'b00000000000000010010001110000011;
ROM[6284] <= 32'b00000000011100011010100000100011;
ROM[6285] <= 32'b00000001000000011010001110000011;
ROM[6286] <= 32'b00000000011100010010000000100011;
ROM[6287] <= 32'b00000000010000010000000100010011;
ROM[6288] <= 32'b00000000011100000000001110010011;
ROM[6289] <= 32'b00000000011100010010000000100011;
ROM[6290] <= 32'b00000000010000010000000100010011;
ROM[6291] <= 32'b11111111110000010000000100010011;
ROM[6292] <= 32'b00000000000000010010001110000011;
ROM[6293] <= 32'b11111111110000010000000100010011;
ROM[6294] <= 32'b00000000000000010010010000000011;
ROM[6295] <= 32'b00000000011101000010001110110011;
ROM[6296] <= 32'b00000000011100010010000000100011;
ROM[6297] <= 32'b00000000010000010000000100010011;
ROM[6298] <= 32'b11111111110000010000000100010011;
ROM[6299] <= 32'b00000000000000010010001110000011;
ROM[6300] <= 32'b01000000011100000000001110110011;
ROM[6301] <= 32'b00000000000100111000001110010011;
ROM[6302] <= 32'b00000000011100010010000000100011;
ROM[6303] <= 32'b00000000010000010000000100010011;
ROM[6304] <= 32'b11111111110000010000000100010011;
ROM[6305] <= 32'b00000000000000010010001110000011;
ROM[6306] <= 32'b00000000000000111000101001100011;
ROM[6307] <= 32'b00000000000000000110001110110111;
ROM[6308] <= 32'b01101001100000111000001110010011;
ROM[6309] <= 32'b00000000111000111000001110110011;
ROM[6310] <= 32'b00000000000000111000000011100111;
ROM[6311] <= 32'b00000001000000011010001110000011;
ROM[6312] <= 32'b00000000011100010010000000100011;
ROM[6313] <= 32'b00000000010000010000000100010011;
ROM[6314] <= 32'b00000001000000011010001110000011;
ROM[6315] <= 32'b00000000011100010010000000100011;
ROM[6316] <= 32'b00000000010000010000000100010011;
ROM[6317] <= 32'b11111111110000010000000100010011;
ROM[6318] <= 32'b00000000000000010010001110000011;
ROM[6319] <= 32'b11111111110000010000000100010011;
ROM[6320] <= 32'b00000000000000010010010000000011;
ROM[6321] <= 32'b00000000011101000000001110110011;
ROM[6322] <= 32'b00000000011100010010000000100011;
ROM[6323] <= 32'b00000000010000010000000100010011;
ROM[6324] <= 32'b00000001000000011010001110000011;
ROM[6325] <= 32'b00000000011100010010000000100011;
ROM[6326] <= 32'b00000000010000010000000100010011;
ROM[6327] <= 32'b11111111110000010000000100010011;
ROM[6328] <= 32'b00000000000000010010001110000011;
ROM[6329] <= 32'b11111111110000010000000100010011;
ROM[6330] <= 32'b00000000000000010010010000000011;
ROM[6331] <= 32'b00000000011101000000001110110011;
ROM[6332] <= 32'b00000000011100010010000000100011;
ROM[6333] <= 32'b00000000010000010000000100010011;
ROM[6334] <= 32'b00000001000000011010001110000011;
ROM[6335] <= 32'b00000000011100010010000000100011;
ROM[6336] <= 32'b00000000010000010000000100010011;
ROM[6337] <= 32'b11111111110000010000000100010011;
ROM[6338] <= 32'b00000000000000010010001110000011;
ROM[6339] <= 32'b11111111110000010000000100010011;
ROM[6340] <= 32'b00000000000000010010010000000011;
ROM[6341] <= 32'b00000000011101000000001110110011;
ROM[6342] <= 32'b00000000011100010010000000100011;
ROM[6343] <= 32'b00000000010000010000000100010011;
ROM[6344] <= 32'b11111111110000010000000100010011;
ROM[6345] <= 32'b00000000000000010010001110000011;
ROM[6346] <= 32'b00000010011100011010100000100011;
ROM[6347] <= 32'b00000000100000011010001110000011;
ROM[6348] <= 32'b00000000011100010010000000100011;
ROM[6349] <= 32'b00000000010000010000000100010011;
ROM[6350] <= 32'b00000000100000011010001110000011;
ROM[6351] <= 32'b00000000011100010010000000100011;
ROM[6352] <= 32'b00000000010000010000000100010011;
ROM[6353] <= 32'b11111111110000010000000100010011;
ROM[6354] <= 32'b00000000000000010010001110000011;
ROM[6355] <= 32'b11111111110000010000000100010011;
ROM[6356] <= 32'b00000000000000010010010000000011;
ROM[6357] <= 32'b00000000011101000000001110110011;
ROM[6358] <= 32'b00000000011100010010000000100011;
ROM[6359] <= 32'b00000000010000010000000100010011;
ROM[6360] <= 32'b00000000100000011010001110000011;
ROM[6361] <= 32'b00000000011100010010000000100011;
ROM[6362] <= 32'b00000000010000010000000100010011;
ROM[6363] <= 32'b11111111110000010000000100010011;
ROM[6364] <= 32'b00000000000000010010001110000011;
ROM[6365] <= 32'b11111111110000010000000100010011;
ROM[6366] <= 32'b00000000000000010010010000000011;
ROM[6367] <= 32'b00000000011101000000001110110011;
ROM[6368] <= 32'b00000000011100010010000000100011;
ROM[6369] <= 32'b00000000010000010000000100010011;
ROM[6370] <= 32'b00000000100000011010001110000011;
ROM[6371] <= 32'b00000000011100010010000000100011;
ROM[6372] <= 32'b00000000010000010000000100010011;
ROM[6373] <= 32'b11111111110000010000000100010011;
ROM[6374] <= 32'b00000000000000010010001110000011;
ROM[6375] <= 32'b11111111110000010000000100010011;
ROM[6376] <= 32'b00000000000000010010010000000011;
ROM[6377] <= 32'b00000000011101000000001110110011;
ROM[6378] <= 32'b00000000011100010010000000100011;
ROM[6379] <= 32'b00000000010000010000000100010011;
ROM[6380] <= 32'b11111111110000010000000100010011;
ROM[6381] <= 32'b00000000000000010010001110000011;
ROM[6382] <= 32'b00000010011100011010011000100011;
ROM[6383] <= 32'b00000010110000011010001110000011;
ROM[6384] <= 32'b00000000011100010010000000100011;
ROM[6385] <= 32'b00000000010000010000000100010011;
ROM[6386] <= 32'b00000111010001101010001110000011;
ROM[6387] <= 32'b00000000011100010010000000100011;
ROM[6388] <= 32'b00000000010000010000000100010011;
ROM[6389] <= 32'b11111111110000010000000100010011;
ROM[6390] <= 32'b00000000000000010010001110000011;
ROM[6391] <= 32'b11111111110000010000000100010011;
ROM[6392] <= 32'b00000000000000010010010000000011;
ROM[6393] <= 32'b00000000011101000000001110110011;
ROM[6394] <= 32'b00000000011100010010000000100011;
ROM[6395] <= 32'b00000000010000010000000100010011;
ROM[6396] <= 32'b11111111110000010000000100010011;
ROM[6397] <= 32'b00000000000000010010001110000011;
ROM[6398] <= 32'b00000000000000111000001100010011;
ROM[6399] <= 32'b00000000110100110000010000110011;
ROM[6400] <= 32'b00000000000001000010001110000011;
ROM[6401] <= 32'b00000000011100010010000000100011;
ROM[6402] <= 32'b00000000010000010000000100010011;
ROM[6403] <= 32'b11111111110000010000000100010011;
ROM[6404] <= 32'b00000000000000010010001110000011;
ROM[6405] <= 32'b00000000011100011010111000100011;
ROM[6406] <= 32'b00000001111100000000001110010011;
ROM[6407] <= 32'b00000000011100010010000000100011;
ROM[6408] <= 32'b00000000010000010000000100010011;
ROM[6409] <= 32'b00000000000000011010001110000011;
ROM[6410] <= 32'b00000000011100010010000000100011;
ROM[6411] <= 32'b00000000010000010000000100010011;
ROM[6412] <= 32'b11111111110000010000000100010011;
ROM[6413] <= 32'b00000000000000010010001110000011;
ROM[6414] <= 32'b11111111110000010000000100010011;
ROM[6415] <= 32'b00000000000000010010010000000011;
ROM[6416] <= 32'b01000000011101000000001110110011;
ROM[6417] <= 32'b00000000011100010010000000100011;
ROM[6418] <= 32'b00000000010000010000000100010011;
ROM[6419] <= 32'b11111111110000010000000100010011;
ROM[6420] <= 32'b00000000000000010010001110000011;
ROM[6421] <= 32'b00000000011100011010110000100011;
ROM[6422] <= 32'b00000000001000000000001110010011;
ROM[6423] <= 32'b00000000011100010010000000100011;
ROM[6424] <= 32'b00000000010000010000000100010011;
ROM[6425] <= 32'b00000001100000011010001110000011;
ROM[6426] <= 32'b00000000011100010010000000100011;
ROM[6427] <= 32'b00000000010000010000000100010011;
ROM[6428] <= 32'b00000000000000000110001110110111;
ROM[6429] <= 32'b01001011110000111000001110010011;
ROM[6430] <= 32'b00000000111000111000001110110011;
ROM[6431] <= 32'b00000000011100010010000000100011;
ROM[6432] <= 32'b00000000010000010000000100010011;
ROM[6433] <= 32'b00000000001100010010000000100011;
ROM[6434] <= 32'b00000000010000010000000100010011;
ROM[6435] <= 32'b00000000010000010010000000100011;
ROM[6436] <= 32'b00000000010000010000000100010011;
ROM[6437] <= 32'b00000000010100010010000000100011;
ROM[6438] <= 32'b00000000010000010000000100010011;
ROM[6439] <= 32'b00000000011000010010000000100011;
ROM[6440] <= 32'b00000000010000010000000100010011;
ROM[6441] <= 32'b00000001010000000000001110010011;
ROM[6442] <= 32'b00000000100000111000001110010011;
ROM[6443] <= 32'b01000000011100010000001110110011;
ROM[6444] <= 32'b00000000011100000000001000110011;
ROM[6445] <= 32'b00000000001000000000000110110011;
ROM[6446] <= 32'b10011001110111111110000011101111;
ROM[6447] <= 32'b11111111110000010000000100010011;
ROM[6448] <= 32'b00000000000000010010001110000011;
ROM[6449] <= 32'b00000010011100011010000000100011;
ROM[6450] <= 32'b00000001110000011010001110000011;
ROM[6451] <= 32'b00000000011100010010000000100011;
ROM[6452] <= 32'b00000000010000010000000100010011;
ROM[6453] <= 32'b00000010000000011010001110000011;
ROM[6454] <= 32'b00000000011100010010000000100011;
ROM[6455] <= 32'b00000000010000010000000100010011;
ROM[6456] <= 32'b00000000000000000110001110110111;
ROM[6457] <= 32'b01010010110000111000001110010011;
ROM[6458] <= 32'b00000000111000111000001110110011;
ROM[6459] <= 32'b00000000011100010010000000100011;
ROM[6460] <= 32'b00000000010000010000000100010011;
ROM[6461] <= 32'b00000000001100010010000000100011;
ROM[6462] <= 32'b00000000010000010000000100010011;
ROM[6463] <= 32'b00000000010000010010000000100011;
ROM[6464] <= 32'b00000000010000010000000100010011;
ROM[6465] <= 32'b00000000010100010010000000100011;
ROM[6466] <= 32'b00000000010000010000000100010011;
ROM[6467] <= 32'b00000000011000010010000000100011;
ROM[6468] <= 32'b00000000010000010000000100010011;
ROM[6469] <= 32'b00000001010000000000001110010011;
ROM[6470] <= 32'b00000000100000111000001110010011;
ROM[6471] <= 32'b01000000011100010000001110110011;
ROM[6472] <= 32'b00000000011100000000001000110011;
ROM[6473] <= 32'b00000000001000000000000110110011;
ROM[6474] <= 32'b11011010010111111011000011101111;
ROM[6475] <= 32'b11111111110000010000000100010011;
ROM[6476] <= 32'b00000000000000010010001110000011;
ROM[6477] <= 32'b00000010011100011010001000100011;
ROM[6478] <= 32'b00000010010000011010001110000011;
ROM[6479] <= 32'b00000000011100010010000000100011;
ROM[6480] <= 32'b00000000010000010000000100010011;
ROM[6481] <= 32'b00000000000100000000001110010011;
ROM[6482] <= 32'b00000000011100010010000000100011;
ROM[6483] <= 32'b00000000010000010000000100010011;
ROM[6484] <= 32'b11111111110000010000000100010011;
ROM[6485] <= 32'b00000000000000010010001110000011;
ROM[6486] <= 32'b11111111110000010000000100010011;
ROM[6487] <= 32'b00000000000000010010010000000011;
ROM[6488] <= 32'b00000000011101000111001110110011;
ROM[6489] <= 32'b00000000011100010010000000100011;
ROM[6490] <= 32'b00000000010000010000000100010011;
ROM[6491] <= 32'b11111111110000010000000100010011;
ROM[6492] <= 32'b00000000000000010010001110000011;
ROM[6493] <= 32'b00000010011100011010010000100011;
ROM[6494] <= 32'b00000010100000011010001110000011;
ROM[6495] <= 32'b00000000011100010010000000100011;
ROM[6496] <= 32'b00000000010000010000000100010011;
ROM[6497] <= 32'b00000000000100000000001110010011;
ROM[6498] <= 32'b00000000011100010010000000100011;
ROM[6499] <= 32'b00000000010000010000000100010011;
ROM[6500] <= 32'b11111111110000010000000100010011;
ROM[6501] <= 32'b00000000000000010010001110000011;
ROM[6502] <= 32'b11111111110000010000000100010011;
ROM[6503] <= 32'b00000000000000010010010000000011;
ROM[6504] <= 32'b00000000011101000010010010110011;
ROM[6505] <= 32'b00000000100000111010010100110011;
ROM[6506] <= 32'b00000000101001001000001110110011;
ROM[6507] <= 32'b00000000000100111000001110010011;
ROM[6508] <= 32'b00000000000100111111001110010011;
ROM[6509] <= 32'b00000000011100010010000000100011;
ROM[6510] <= 32'b00000000010000010000000100010011;
ROM[6511] <= 32'b11111111110000010000000100010011;
ROM[6512] <= 32'b00000000000000010010001110000011;
ROM[6513] <= 32'b00000000000000111000101001100011;
ROM[6514] <= 32'b00000000000000000110001110110111;
ROM[6515] <= 32'b01011101110000111000001110010011;
ROM[6516] <= 32'b00000000111000111000001110110011;
ROM[6517] <= 32'b00000000000000111000000011100111;
ROM[6518] <= 32'b00000100100000000000000011101111;
ROM[6519] <= 32'b00000001110000011010001110000011;
ROM[6520] <= 32'b00000000011100010010000000100011;
ROM[6521] <= 32'b00000000010000010000000100010011;
ROM[6522] <= 32'b00000010000000011010001110000011;
ROM[6523] <= 32'b00000000011100010010000000100011;
ROM[6524] <= 32'b00000000010000010000000100010011;
ROM[6525] <= 32'b11111111110000010000000100010011;
ROM[6526] <= 32'b00000000000000010010001110000011;
ROM[6527] <= 32'b11111111110000010000000100010011;
ROM[6528] <= 32'b00000000000000010010010000000011;
ROM[6529] <= 32'b01000000011101000000001110110011;
ROM[6530] <= 32'b00000000011100010010000000100011;
ROM[6531] <= 32'b00000000010000010000000100010011;
ROM[6532] <= 32'b11111111110000010000000100010011;
ROM[6533] <= 32'b00000000000000010010001110000011;
ROM[6534] <= 32'b00000000011100011010111000100011;
ROM[6535] <= 32'b00000000010000000000000011101111;
ROM[6536] <= 32'b00000010110000011010001110000011;
ROM[6537] <= 32'b00000000011100010010000000100011;
ROM[6538] <= 32'b00000000010000010000000100010011;
ROM[6539] <= 32'b00000111010001101010001110000011;
ROM[6540] <= 32'b00000000011100010010000000100011;
ROM[6541] <= 32'b00000000010000010000000100010011;
ROM[6542] <= 32'b11111111110000010000000100010011;
ROM[6543] <= 32'b00000000000000010010001110000011;
ROM[6544] <= 32'b11111111110000010000000100010011;
ROM[6545] <= 32'b00000000000000010010010000000011;
ROM[6546] <= 32'b00000000011101000000001110110011;
ROM[6547] <= 32'b00000000011100010010000000100011;
ROM[6548] <= 32'b00000000010000010000000100010011;
ROM[6549] <= 32'b00000001110000011010001110000011;
ROM[6550] <= 32'b00000000011100010010000000100011;
ROM[6551] <= 32'b00000000010000010000000100010011;
ROM[6552] <= 32'b11111111110000010000000100010011;
ROM[6553] <= 32'b00000000000000010010001110000011;
ROM[6554] <= 32'b00000000011101100010000000100011;
ROM[6555] <= 32'b11111111110000010000000100010011;
ROM[6556] <= 32'b00000000000000010010001110000011;
ROM[6557] <= 32'b00000000000000111000001100010011;
ROM[6558] <= 32'b00000000000001100010001110000011;
ROM[6559] <= 32'b00000000011100010010000000100011;
ROM[6560] <= 32'b00000000010000010000000100010011;
ROM[6561] <= 32'b11111111110000010000000100010011;
ROM[6562] <= 32'b00000000000000010010001110000011;
ROM[6563] <= 32'b00000000110100110000010000110011;
ROM[6564] <= 32'b00000000011101000010000000100011;
ROM[6565] <= 32'b10111010000111111111000011101111;
ROM[6566] <= 32'b00000000000000011010001110000011;
ROM[6567] <= 32'b00000000011100010010000000100011;
ROM[6568] <= 32'b00000000010000010000000100010011;
ROM[6569] <= 32'b00000000000100000000001110010011;
ROM[6570] <= 32'b00000000011100010010000000100011;
ROM[6571] <= 32'b00000000010000010000000100010011;
ROM[6572] <= 32'b11111111110000010000000100010011;
ROM[6573] <= 32'b00000000000000010010001110000011;
ROM[6574] <= 32'b11111111110000010000000100010011;
ROM[6575] <= 32'b00000000000000010010010000000011;
ROM[6576] <= 32'b00000000011101000000001110110011;
ROM[6577] <= 32'b00000000011100010010000000100011;
ROM[6578] <= 32'b00000000010000010000000100010011;
ROM[6579] <= 32'b11111111110000010000000100010011;
ROM[6580] <= 32'b00000000000000010010001110000011;
ROM[6581] <= 32'b00000000011100011010000000100011;
ROM[6582] <= 32'b00000000110000011010001110000011;
ROM[6583] <= 32'b00000000011100010010000000100011;
ROM[6584] <= 32'b00000000010000010000000100010011;
ROM[6585] <= 32'b00000000000100000000001110010011;
ROM[6586] <= 32'b00000000011100010010000000100011;
ROM[6587] <= 32'b00000000010000010000000100010011;
ROM[6588] <= 32'b11111111110000010000000100010011;
ROM[6589] <= 32'b00000000000000010010001110000011;
ROM[6590] <= 32'b11111111110000010000000100010011;
ROM[6591] <= 32'b00000000000000010010010000000011;
ROM[6592] <= 32'b00000000011101000000001110110011;
ROM[6593] <= 32'b00000000011100010010000000100011;
ROM[6594] <= 32'b00000000010000010000000100010011;
ROM[6595] <= 32'b11111111110000010000000100010011;
ROM[6596] <= 32'b00000000000000010010001110000011;
ROM[6597] <= 32'b00000000011100011010011000100011;
ROM[6598] <= 32'b00000000000000011010001110000011;
ROM[6599] <= 32'b00000000011100010010000000100011;
ROM[6600] <= 32'b00000000010000010000000100010011;
ROM[6601] <= 32'b00000010000000000000001110010011;
ROM[6602] <= 32'b00000000011100010010000000100011;
ROM[6603] <= 32'b00000000010000010000000100010011;
ROM[6604] <= 32'b11111111110000010000000100010011;
ROM[6605] <= 32'b00000000000000010010001110000011;
ROM[6606] <= 32'b11111111110000010000000100010011;
ROM[6607] <= 32'b00000000000000010010010000000011;
ROM[6608] <= 32'b00000000011101000010010010110011;
ROM[6609] <= 32'b00000000100000111010010100110011;
ROM[6610] <= 32'b00000000101001001000001110110011;
ROM[6611] <= 32'b00000000000100111000001110010011;
ROM[6612] <= 32'b00000000000100111111001110010011;
ROM[6613] <= 32'b00000000011100010010000000100011;
ROM[6614] <= 32'b00000000010000010000000100010011;
ROM[6615] <= 32'b11111111110000010000000100010011;
ROM[6616] <= 32'b00000000000000010010001110000011;
ROM[6617] <= 32'b00000000000000111000101001100011;
ROM[6618] <= 32'b00000000000000000110001110110111;
ROM[6619] <= 32'b01110111110000111000001110010011;
ROM[6620] <= 32'b00000000111000111000001110110011;
ROM[6621] <= 32'b00000000000000111000000011100111;
ROM[6622] <= 32'b00000110000000000000000011101111;
ROM[6623] <= 32'b00000000000000000000001110010011;
ROM[6624] <= 32'b00000000011100010010000000100011;
ROM[6625] <= 32'b00000000010000010000000100010011;
ROM[6626] <= 32'b11111111110000010000000100010011;
ROM[6627] <= 32'b00000000000000010010001110000011;
ROM[6628] <= 32'b00000000011100011010000000100011;
ROM[6629] <= 32'b00000000100000011010001110000011;
ROM[6630] <= 32'b00000000011100010010000000100011;
ROM[6631] <= 32'b00000000010000010000000100010011;
ROM[6632] <= 32'b00000000000100000000001110010011;
ROM[6633] <= 32'b00000000011100010010000000100011;
ROM[6634] <= 32'b00000000010000010000000100010011;
ROM[6635] <= 32'b11111111110000010000000100010011;
ROM[6636] <= 32'b00000000000000010010001110000011;
ROM[6637] <= 32'b11111111110000010000000100010011;
ROM[6638] <= 32'b00000000000000010010010000000011;
ROM[6639] <= 32'b00000000011101000000001110110011;
ROM[6640] <= 32'b00000000011100010010000000100011;
ROM[6641] <= 32'b00000000010000010000000100010011;
ROM[6642] <= 32'b11111111110000010000000100010011;
ROM[6643] <= 32'b00000000000000010010001110000011;
ROM[6644] <= 32'b00000000011100011010010000100011;
ROM[6645] <= 32'b00000000010000000000000011101111;
ROM[6646] <= 32'b10011101110111111111000011101111;
ROM[6647] <= 32'b00000000000000000000001110010011;
ROM[6648] <= 32'b00000000011100010010000000100011;
ROM[6649] <= 32'b00000000010000010000000100010011;
ROM[6650] <= 32'b00000001010000000000001110010011;
ROM[6651] <= 32'b01000000011100011000001110110011;
ROM[6652] <= 32'b00000000000000111010000010000011;
ROM[6653] <= 32'b11111111110000010000000100010011;
ROM[6654] <= 32'b00000000000000010010001110000011;
ROM[6655] <= 32'b00000000011100100010000000100011;
ROM[6656] <= 32'b00000000010000100000000100010011;
ROM[6657] <= 32'b00000001010000000000001110010011;
ROM[6658] <= 32'b01000000011100011000001110110011;
ROM[6659] <= 32'b00000000010000111010000110000011;
ROM[6660] <= 32'b00000000100000111010001000000011;
ROM[6661] <= 32'b00000000110000111010001010000011;
ROM[6662] <= 32'b00000001000000111010001100000011;
ROM[6663] <= 32'b00000000000000001000000011100111;
ROM[6664] <= 32'b00000000001100000000001110010011;
ROM[6665] <= 32'b00000000011100010010000000100011;
ROM[6666] <= 32'b00000000010000010000000100010011;
ROM[6667] <= 32'b00000000000000000111001110110111;
ROM[6668] <= 32'b10000111100000111000001110010011;
ROM[6669] <= 32'b00000000111000111000001110110011;
ROM[6670] <= 32'b00000000011100010010000000100011;
ROM[6671] <= 32'b00000000010000010000000100010011;
ROM[6672] <= 32'b00000000001100010010000000100011;
ROM[6673] <= 32'b00000000010000010000000100010011;
ROM[6674] <= 32'b00000000010000010010000000100011;
ROM[6675] <= 32'b00000000010000010000000100010011;
ROM[6676] <= 32'b00000000010100010010000000100011;
ROM[6677] <= 32'b00000000010000010000000100010011;
ROM[6678] <= 32'b00000000011000010010000000100011;
ROM[6679] <= 32'b00000000010000010000000100010011;
ROM[6680] <= 32'b00000001010000000000001110010011;
ROM[6681] <= 32'b00000000010000111000001110010011;
ROM[6682] <= 32'b01000000011100010000001110110011;
ROM[6683] <= 32'b00000000011100000000001000110011;
ROM[6684] <= 32'b00000000001000000000000110110011;
ROM[6685] <= 32'b10110110100111111100000011101111;
ROM[6686] <= 32'b11111111110000010000000100010011;
ROM[6687] <= 32'b00000000000000010010001110000011;
ROM[6688] <= 32'b00000000000000111000001010010011;
ROM[6689] <= 32'b00000000000000100010001110000011;
ROM[6690] <= 32'b00000000011100010010000000100011;
ROM[6691] <= 32'b00000000010000010000000100010011;
ROM[6692] <= 32'b00000000000000000000001110010011;
ROM[6693] <= 32'b00000000011100010010000000100011;
ROM[6694] <= 32'b00000000010000010000000100010011;
ROM[6695] <= 32'b11111111110000010000000100010011;
ROM[6696] <= 32'b00000000000000010010001110000011;
ROM[6697] <= 32'b11111111110000010000000100010011;
ROM[6698] <= 32'b00000000000000010010010000000011;
ROM[6699] <= 32'b00000000011101000010010010110011;
ROM[6700] <= 32'b00000000100000111010010100110011;
ROM[6701] <= 32'b00000000101001001000001110110011;
ROM[6702] <= 32'b00000000000100111000001110010011;
ROM[6703] <= 32'b00000000000100111111001110010011;
ROM[6704] <= 32'b00000000011100010010000000100011;
ROM[6705] <= 32'b00000000010000010000000100010011;
ROM[6706] <= 32'b11111111110000010000000100010011;
ROM[6707] <= 32'b00000000000000010010001110000011;
ROM[6708] <= 32'b00000000000000111000101001100011;
ROM[6709] <= 32'b00000000000000000111001110110111;
ROM[6710] <= 32'b10001110100000111000001110010011;
ROM[6711] <= 32'b00000000111000111000001110110011;
ROM[6712] <= 32'b00000000000000111000000011100111;
ROM[6713] <= 32'b00000010000000000000000011101111;
ROM[6714] <= 32'b00000000000100000000001110010011;
ROM[6715] <= 32'b00000000011100010010000000100011;
ROM[6716] <= 32'b00000000010000010000000100010011;
ROM[6717] <= 32'b11111111110000010000000100010011;
ROM[6718] <= 32'b00000000000000010010001110000011;
ROM[6719] <= 32'b00000000011100100010000000100011;
ROM[6720] <= 32'b00000000010000000000000011101111;
ROM[6721] <= 32'b00000000000000000000001110010011;
ROM[6722] <= 32'b00000000011100010010000000100011;
ROM[6723] <= 32'b00000000010000010000000100010011;
ROM[6724] <= 32'b11111111110000010000000100010011;
ROM[6725] <= 32'b00000000000000010010001110000011;
ROM[6726] <= 32'b00000000110100101000010000110011;
ROM[6727] <= 32'b00000000011101000010001000100011;
ROM[6728] <= 32'b00000000000000100010001110000011;
ROM[6729] <= 32'b00000000011100010010000000100011;
ROM[6730] <= 32'b00000000010000010000000100010011;
ROM[6731] <= 32'b11111111110000010000000100010011;
ROM[6732] <= 32'b00000000000000010010001110000011;
ROM[6733] <= 32'b00000000110100101000010000110011;
ROM[6734] <= 32'b00000000011101000010000000100011;
ROM[6735] <= 32'b00000000000000100010001110000011;
ROM[6736] <= 32'b00000000011100010010000000100011;
ROM[6737] <= 32'b00000000010000010000000100010011;
ROM[6738] <= 32'b00000000000000000111001110110111;
ROM[6739] <= 32'b10011001010000111000001110010011;
ROM[6740] <= 32'b00000000111000111000001110110011;
ROM[6741] <= 32'b00000000011100010010000000100011;
ROM[6742] <= 32'b00000000010000010000000100010011;
ROM[6743] <= 32'b00000000001100010010000000100011;
ROM[6744] <= 32'b00000000010000010000000100010011;
ROM[6745] <= 32'b00000000010000010010000000100011;
ROM[6746] <= 32'b00000000010000010000000100010011;
ROM[6747] <= 32'b00000000010100010010000000100011;
ROM[6748] <= 32'b00000000010000010000000100010011;
ROM[6749] <= 32'b00000000011000010010000000100011;
ROM[6750] <= 32'b00000000010000010000000100010011;
ROM[6751] <= 32'b00000001010000000000001110010011;
ROM[6752] <= 32'b00000000010000111000001110010011;
ROM[6753] <= 32'b01000000011100010000001110110011;
ROM[6754] <= 32'b00000000011100000000001000110011;
ROM[6755] <= 32'b00000000001000000000000110110011;
ROM[6756] <= 32'b10101011000111111001000011101111;
ROM[6757] <= 32'b11111111110000010000000100010011;
ROM[6758] <= 32'b00000000000000010010001110000011;
ROM[6759] <= 32'b00000000110100101000010000110011;
ROM[6760] <= 32'b00000000011101000010010000100011;
ROM[6761] <= 32'b00000000000000010010001010000011;
ROM[6762] <= 32'b00000000010000010000000100010011;
ROM[6763] <= 32'b00000001010000000000001110010011;
ROM[6764] <= 32'b01000000011100011000001110110011;
ROM[6765] <= 32'b00000000000000111010000010000011;
ROM[6766] <= 32'b11111111110000010000000100010011;
ROM[6767] <= 32'b00000000000000010010001110000011;
ROM[6768] <= 32'b00000000011100100010000000100011;
ROM[6769] <= 32'b00000000010000100000000100010011;
ROM[6770] <= 32'b00000001010000000000001110010011;
ROM[6771] <= 32'b01000000011100011000001110110011;
ROM[6772] <= 32'b00000000010000111010000110000011;
ROM[6773] <= 32'b00000000100000111010001000000011;
ROM[6774] <= 32'b00000000110000111010001010000011;
ROM[6775] <= 32'b00000001000000111010001100000011;
ROM[6776] <= 32'b00000000000000001000000011100111;
ROM[6777] <= 32'b00000000000000100010001110000011;
ROM[6778] <= 32'b00000000011100010010000000100011;
ROM[6779] <= 32'b00000000010000010000000100010011;
ROM[6780] <= 32'b11111111110000010000000100010011;
ROM[6781] <= 32'b00000000000000010010001110000011;
ROM[6782] <= 32'b00000000000000111000001010010011;
ROM[6783] <= 32'b00000000110100101000010000110011;
ROM[6784] <= 32'b00000000010001000010001110000011;
ROM[6785] <= 32'b00000000011100010010000000100011;
ROM[6786] <= 32'b00000000010000010000000100010011;
ROM[6787] <= 32'b00000001010000000000001110010011;
ROM[6788] <= 32'b01000000011100011000001110110011;
ROM[6789] <= 32'b00000000000000111010000010000011;
ROM[6790] <= 32'b11111111110000010000000100010011;
ROM[6791] <= 32'b00000000000000010010001110000011;
ROM[6792] <= 32'b00000000011100100010000000100011;
ROM[6793] <= 32'b00000000010000100000000100010011;
ROM[6794] <= 32'b00000001010000000000001110010011;
ROM[6795] <= 32'b01000000011100011000001110110011;
ROM[6796] <= 32'b00000000010000111010000110000011;
ROM[6797] <= 32'b00000000100000111010001000000011;
ROM[6798] <= 32'b00000000110000111010001010000011;
ROM[6799] <= 32'b00000001000000111010001100000011;
ROM[6800] <= 32'b00000000000000001000000011100111;
ROM[6801] <= 32'b00000000000000100010001110000011;
ROM[6802] <= 32'b00000000011100010010000000100011;
ROM[6803] <= 32'b00000000010000010000000100010011;
ROM[6804] <= 32'b11111111110000010000000100010011;
ROM[6805] <= 32'b00000000000000010010001110000011;
ROM[6806] <= 32'b00000000000000111000001010010011;
ROM[6807] <= 32'b00000000010000100010001110000011;
ROM[6808] <= 32'b00000000011100010010000000100011;
ROM[6809] <= 32'b00000000010000010000000100010011;
ROM[6810] <= 32'b00000000110100101000010000110011;
ROM[6811] <= 32'b00000000100001000010001110000011;
ROM[6812] <= 32'b00000000011100010010000000100011;
ROM[6813] <= 32'b00000000010000010000000100010011;
ROM[6814] <= 32'b11111111110000010000000100010011;
ROM[6815] <= 32'b00000000000000010010001110000011;
ROM[6816] <= 32'b11111111110000010000000100010011;
ROM[6817] <= 32'b00000000000000010010010000000011;
ROM[6818] <= 32'b00000000011101000000001110110011;
ROM[6819] <= 32'b00000000011100010010000000100011;
ROM[6820] <= 32'b00000000010000010000000100010011;
ROM[6821] <= 32'b11111111110000010000000100010011;
ROM[6822] <= 32'b00000000000000010010001110000011;
ROM[6823] <= 32'b00000000000000111000001100010011;
ROM[6824] <= 32'b00000000110100110000010000110011;
ROM[6825] <= 32'b00000000000001000010001110000011;
ROM[6826] <= 32'b00000000011100010010000000100011;
ROM[6827] <= 32'b00000000010000010000000100010011;
ROM[6828] <= 32'b00000001010000000000001110010011;
ROM[6829] <= 32'b01000000011100011000001110110011;
ROM[6830] <= 32'b00000000000000111010000010000011;
ROM[6831] <= 32'b11111111110000010000000100010011;
ROM[6832] <= 32'b00000000000000010010001110000011;
ROM[6833] <= 32'b00000000011100100010000000100011;
ROM[6834] <= 32'b00000000010000100000000100010011;
ROM[6835] <= 32'b00000001010000000000001110010011;
ROM[6836] <= 32'b01000000011100011000001110110011;
ROM[6837] <= 32'b00000000010000111010000110000011;
ROM[6838] <= 32'b00000000100000111010001000000011;
ROM[6839] <= 32'b00000000110000111010001010000011;
ROM[6840] <= 32'b00000001000000111010001100000011;
ROM[6841] <= 32'b00000000000000001000000011100111;
ROM[6842] <= 32'b00000000000000100010001110000011;
ROM[6843] <= 32'b00000000011100010010000000100011;
ROM[6844] <= 32'b00000000010000010000000100010011;
ROM[6845] <= 32'b11111111110000010000000100010011;
ROM[6846] <= 32'b00000000000000010010001110000011;
ROM[6847] <= 32'b00000000000000111000001010010011;
ROM[6848] <= 32'b00000000010000100010001110000011;
ROM[6849] <= 32'b00000000011100010010000000100011;
ROM[6850] <= 32'b00000000010000010000000100010011;
ROM[6851] <= 32'b00000000110100101000010000110011;
ROM[6852] <= 32'b00000000100001000010001110000011;
ROM[6853] <= 32'b00000000011100010010000000100011;
ROM[6854] <= 32'b00000000010000010000000100010011;
ROM[6855] <= 32'b11111111110000010000000100010011;
ROM[6856] <= 32'b00000000000000010010001110000011;
ROM[6857] <= 32'b11111111110000010000000100010011;
ROM[6858] <= 32'b00000000000000010010010000000011;
ROM[6859] <= 32'b00000000011101000000001110110011;
ROM[6860] <= 32'b00000000011100010010000000100011;
ROM[6861] <= 32'b00000000010000010000000100010011;
ROM[6862] <= 32'b00000000100000100010001110000011;
ROM[6863] <= 32'b00000000011100010010000000100011;
ROM[6864] <= 32'b00000000010000010000000100010011;
ROM[6865] <= 32'b11111111110000010000000100010011;
ROM[6866] <= 32'b00000000000000010010001110000011;
ROM[6867] <= 32'b00000000011101100010000000100011;
ROM[6868] <= 32'b11111111110000010000000100010011;
ROM[6869] <= 32'b00000000000000010010001110000011;
ROM[6870] <= 32'b00000000000000111000001100010011;
ROM[6871] <= 32'b00000000000001100010001110000011;
ROM[6872] <= 32'b00000000011100010010000000100011;
ROM[6873] <= 32'b00000000010000010000000100010011;
ROM[6874] <= 32'b11111111110000010000000100010011;
ROM[6875] <= 32'b00000000000000010010001110000011;
ROM[6876] <= 32'b00000000110100110000010000110011;
ROM[6877] <= 32'b00000000011101000010000000100011;
ROM[6878] <= 32'b00000000000000000000001110010011;
ROM[6879] <= 32'b00000000011100010010000000100011;
ROM[6880] <= 32'b00000000010000010000000100010011;
ROM[6881] <= 32'b00000001010000000000001110010011;
ROM[6882] <= 32'b01000000011100011000001110110011;
ROM[6883] <= 32'b00000000000000111010000010000011;
ROM[6884] <= 32'b11111111110000010000000100010011;
ROM[6885] <= 32'b00000000000000010010001110000011;
ROM[6886] <= 32'b00000000011100100010000000100011;
ROM[6887] <= 32'b00000000010000100000000100010011;
ROM[6888] <= 32'b00000001010000000000001110010011;
ROM[6889] <= 32'b01000000011100011000001110110011;
ROM[6890] <= 32'b00000000010000111010000110000011;
ROM[6891] <= 32'b00000000100000111010001000000011;
ROM[6892] <= 32'b00000000110000111010001010000011;
ROM[6893] <= 32'b00000001000000111010001100000011;
ROM[6894] <= 32'b00000000000000001000000011100111;
ROM[6895] <= 32'b00000000000000100010001110000011;
ROM[6896] <= 32'b00000000011100010010000000100011;
ROM[6897] <= 32'b00000000010000010000000100010011;
ROM[6898] <= 32'b11111111110000010000000100010011;
ROM[6899] <= 32'b00000000000000010010001110000011;
ROM[6900] <= 32'b00000000000000111000001010010011;
ROM[6901] <= 32'b00000000110100101000010000110011;
ROM[6902] <= 32'b00000000010001000010001110000011;
ROM[6903] <= 32'b00000000011100010010000000100011;
ROM[6904] <= 32'b00000000010000010000000100010011;
ROM[6905] <= 32'b00000000110100101000010000110011;
ROM[6906] <= 32'b00000000000001000010001110000011;
ROM[6907] <= 32'b00000000011100010010000000100011;
ROM[6908] <= 32'b00000000010000010000000100010011;
ROM[6909] <= 32'b11111111110000010000000100010011;
ROM[6910] <= 32'b00000000000000010010001110000011;
ROM[6911] <= 32'b11111111110000010000000100010011;
ROM[6912] <= 32'b00000000000000010010010000000011;
ROM[6913] <= 32'b00000000011101000010001110110011;
ROM[6914] <= 32'b00000000011100010010000000100011;
ROM[6915] <= 32'b00000000010000010000000100010011;
ROM[6916] <= 32'b11111111110000010000000100010011;
ROM[6917] <= 32'b00000000000000010010001110000011;
ROM[6918] <= 32'b00000000000000111000101001100011;
ROM[6919] <= 32'b00000000000000000111001110110111;
ROM[6920] <= 32'b11000011000000111000001110010011;
ROM[6921] <= 32'b00000000111000111000001110110011;
ROM[6922] <= 32'b00000000000000111000000011100111;
ROM[6923] <= 32'b00001100110000000000000011101111;
ROM[6924] <= 32'b00000000110100101000010000110011;
ROM[6925] <= 32'b00000000010001000010001110000011;
ROM[6926] <= 32'b00000000011100010010000000100011;
ROM[6927] <= 32'b00000000010000010000000100010011;
ROM[6928] <= 32'b00000000110100101000010000110011;
ROM[6929] <= 32'b00000000100001000010001110000011;
ROM[6930] <= 32'b00000000011100010010000000100011;
ROM[6931] <= 32'b00000000010000010000000100010011;
ROM[6932] <= 32'b11111111110000010000000100010011;
ROM[6933] <= 32'b00000000000000010010001110000011;
ROM[6934] <= 32'b11111111110000010000000100010011;
ROM[6935] <= 32'b00000000000000010010010000000011;
ROM[6936] <= 32'b00000000011101000000001110110011;
ROM[6937] <= 32'b00000000011100010010000000100011;
ROM[6938] <= 32'b00000000010000010000000100010011;
ROM[6939] <= 32'b00000000010000100010001110000011;
ROM[6940] <= 32'b00000000011100010010000000100011;
ROM[6941] <= 32'b00000000010000010000000100010011;
ROM[6942] <= 32'b11111111110000010000000100010011;
ROM[6943] <= 32'b00000000000000010010001110000011;
ROM[6944] <= 32'b00000000011101100010000000100011;
ROM[6945] <= 32'b11111111110000010000000100010011;
ROM[6946] <= 32'b00000000000000010010001110000011;
ROM[6947] <= 32'b00000000000000111000001100010011;
ROM[6948] <= 32'b00000000000001100010001110000011;
ROM[6949] <= 32'b00000000011100010010000000100011;
ROM[6950] <= 32'b00000000010000010000000100010011;
ROM[6951] <= 32'b11111111110000010000000100010011;
ROM[6952] <= 32'b00000000000000010010001110000011;
ROM[6953] <= 32'b00000000110100110000010000110011;
ROM[6954] <= 32'b00000000011101000010000000100011;
ROM[6955] <= 32'b00000000110100101000010000110011;
ROM[6956] <= 32'b00000000010001000010001110000011;
ROM[6957] <= 32'b00000000011100010010000000100011;
ROM[6958] <= 32'b00000000010000010000000100010011;
ROM[6959] <= 32'b00000000000100000000001110010011;
ROM[6960] <= 32'b00000000011100010010000000100011;
ROM[6961] <= 32'b00000000010000010000000100010011;
ROM[6962] <= 32'b11111111110000010000000100010011;
ROM[6963] <= 32'b00000000000000010010001110000011;
ROM[6964] <= 32'b11111111110000010000000100010011;
ROM[6965] <= 32'b00000000000000010010010000000011;
ROM[6966] <= 32'b00000000011101000000001110110011;
ROM[6967] <= 32'b00000000011100010010000000100011;
ROM[6968] <= 32'b00000000010000010000000100010011;
ROM[6969] <= 32'b11111111110000010000000100010011;
ROM[6970] <= 32'b00000000000000010010001110000011;
ROM[6971] <= 32'b00000000110100101000010000110011;
ROM[6972] <= 32'b00000000011101000010001000100011;
ROM[6973] <= 32'b00000000010000000000000011101111;
ROM[6974] <= 32'b00000000110100101000010000110011;
ROM[6975] <= 32'b00000000100001000010001110000011;
ROM[6976] <= 32'b00000000011100010010000000100011;
ROM[6977] <= 32'b00000000010000010000000100010011;
ROM[6978] <= 32'b00000001010000000000001110010011;
ROM[6979] <= 32'b01000000011100011000001110110011;
ROM[6980] <= 32'b00000000000000111010000010000011;
ROM[6981] <= 32'b11111111110000010000000100010011;
ROM[6982] <= 32'b00000000000000010010001110000011;
ROM[6983] <= 32'b00000000011100100010000000100011;
ROM[6984] <= 32'b00000000010000100000000100010011;
ROM[6985] <= 32'b00000001010000000000001110010011;
ROM[6986] <= 32'b01000000011100011000001110110011;
ROM[6987] <= 32'b00000000010000111010000110000011;
ROM[6988] <= 32'b00000000100000111010001000000011;
ROM[6989] <= 32'b00000000110000111010001010000011;
ROM[6990] <= 32'b00000001000000111010001100000011;
ROM[6991] <= 32'b00000000000000001000000011100111;
ROM[6992] <= 32'b00000000000000100010001110000011;
ROM[6993] <= 32'b00000000011100010010000000100011;
ROM[6994] <= 32'b00000000010000010000000100010011;
ROM[6995] <= 32'b11111111110000010000000100010011;
ROM[6996] <= 32'b00000000000000010010001110000011;
ROM[6997] <= 32'b00000000000000111000001010010011;
ROM[6998] <= 32'b00000000110100101000010000110011;
ROM[6999] <= 32'b00000000010001000010001110000011;
ROM[7000] <= 32'b00000000011100010010000000100011;
ROM[7001] <= 32'b00000000010000010000000100010011;
ROM[7002] <= 32'b00000000000000000000001110010011;
ROM[7003] <= 32'b00000000011100010010000000100011;
ROM[7004] <= 32'b00000000010000010000000100010011;
ROM[7005] <= 32'b11111111110000010000000100010011;
ROM[7006] <= 32'b00000000000000010010001110000011;
ROM[7007] <= 32'b11111111110000010000000100010011;
ROM[7008] <= 32'b00000000000000010010010000000011;
ROM[7009] <= 32'b00000000100000111010001110110011;
ROM[7010] <= 32'b00000000011100010010000000100011;
ROM[7011] <= 32'b00000000010000010000000100010011;
ROM[7012] <= 32'b11111111110000010000000100010011;
ROM[7013] <= 32'b00000000000000010010001110000011;
ROM[7014] <= 32'b00000000000000111000101001100011;
ROM[7015] <= 32'b00000000000000000111001110110111;
ROM[7016] <= 32'b11011011000000111000001110010011;
ROM[7017] <= 32'b00000000111000111000001110110011;
ROM[7018] <= 32'b00000000000000111000000011100111;
ROM[7019] <= 32'b00000101000000000000000011101111;
ROM[7020] <= 32'b00000000110100101000010000110011;
ROM[7021] <= 32'b00000000010001000010001110000011;
ROM[7022] <= 32'b00000000011100010010000000100011;
ROM[7023] <= 32'b00000000010000010000000100010011;
ROM[7024] <= 32'b00000000000100000000001110010011;
ROM[7025] <= 32'b00000000011100010010000000100011;
ROM[7026] <= 32'b00000000010000010000000100010011;
ROM[7027] <= 32'b11111111110000010000000100010011;
ROM[7028] <= 32'b00000000000000010010001110000011;
ROM[7029] <= 32'b11111111110000010000000100010011;
ROM[7030] <= 32'b00000000000000010010010000000011;
ROM[7031] <= 32'b01000000011101000000001110110011;
ROM[7032] <= 32'b00000000011100010010000000100011;
ROM[7033] <= 32'b00000000010000010000000100010011;
ROM[7034] <= 32'b11111111110000010000000100010011;
ROM[7035] <= 32'b00000000000000010010001110000011;
ROM[7036] <= 32'b00000000110100101000010000110011;
ROM[7037] <= 32'b00000000011101000010001000100011;
ROM[7038] <= 32'b00000000010000000000000011101111;
ROM[7039] <= 32'b00000000000000000000001110010011;
ROM[7040] <= 32'b00000000011100010010000000100011;
ROM[7041] <= 32'b00000000010000010000000100010011;
ROM[7042] <= 32'b00000001010000000000001110010011;
ROM[7043] <= 32'b01000000011100011000001110110011;
ROM[7044] <= 32'b00000000000000111010000010000011;
ROM[7045] <= 32'b11111111110000010000000100010011;
ROM[7046] <= 32'b00000000000000010010001110000011;
ROM[7047] <= 32'b00000000011100100010000000100011;
ROM[7048] <= 32'b00000000010000100000000100010011;
ROM[7049] <= 32'b00000001010000000000001110010011;
ROM[7050] <= 32'b01000000011100011000001110110011;
ROM[7051] <= 32'b00000000010000111010000110000011;
ROM[7052] <= 32'b00000000100000111010001000000011;
ROM[7053] <= 32'b00000000110000111010001010000011;
ROM[7054] <= 32'b00000001000000111010001100000011;
ROM[7055] <= 32'b00000000000000001000000011100111;
ROM[7056] <= 32'b00000000000000010010000000100011;
ROM[7057] <= 32'b00000000010000010000000100010011;
ROM[7058] <= 32'b00000000000000010010000000100011;
ROM[7059] <= 32'b00000000010000010000000100010011;
ROM[7060] <= 32'b00000000000000010010000000100011;
ROM[7061] <= 32'b00000000010000010000000100010011;
ROM[7062] <= 32'b00000000000000100010001110000011;
ROM[7063] <= 32'b00000000011100010010000000100011;
ROM[7064] <= 32'b00000000010000010000000100010011;
ROM[7065] <= 32'b11111111110000010000000100010011;
ROM[7066] <= 32'b00000000000000010010001110000011;
ROM[7067] <= 32'b00000000000000111000001010010011;
ROM[7068] <= 32'b00000000000000000000001110010011;
ROM[7069] <= 32'b00000000011100010010000000100011;
ROM[7070] <= 32'b00000000010000010000000100010011;
ROM[7071] <= 32'b11111111110000010000000100010011;
ROM[7072] <= 32'b00000000000000010010001110000011;
ROM[7073] <= 32'b00000000011100011010000000100011;
ROM[7074] <= 32'b00000000110100101000010000110011;
ROM[7075] <= 32'b00000000010001000010001110000011;
ROM[7076] <= 32'b00000000011100010010000000100011;
ROM[7077] <= 32'b00000000010000010000000100010011;
ROM[7078] <= 32'b00000000000000000000001110010011;
ROM[7079] <= 32'b00000000011100010010000000100011;
ROM[7080] <= 32'b00000000010000010000000100010011;
ROM[7081] <= 32'b11111111110000010000000100010011;
ROM[7082] <= 32'b00000000000000010010001110000011;
ROM[7083] <= 32'b11111111110000010000000100010011;
ROM[7084] <= 32'b00000000000000010010010000000011;
ROM[7085] <= 32'b00000000100000111010001110110011;
ROM[7086] <= 32'b00000000011100010010000000100011;
ROM[7087] <= 32'b00000000010000010000000100010011;
ROM[7088] <= 32'b00000000000000000000001110010011;
ROM[7089] <= 32'b00000000011100010010000000100011;
ROM[7090] <= 32'b00000000010000010000000100010011;
ROM[7091] <= 32'b00000000110100101000010000110011;
ROM[7092] <= 32'b00000000100001000010001110000011;
ROM[7093] <= 32'b00000000011100010010000000100011;
ROM[7094] <= 32'b00000000010000010000000100010011;
ROM[7095] <= 32'b11111111110000010000000100010011;
ROM[7096] <= 32'b00000000000000010010001110000011;
ROM[7097] <= 32'b11111111110000010000000100010011;
ROM[7098] <= 32'b00000000000000010010010000000011;
ROM[7099] <= 32'b00000000011101000000001110110011;
ROM[7100] <= 32'b00000000011100010010000000100011;
ROM[7101] <= 32'b00000000010000010000000100010011;
ROM[7102] <= 32'b11111111110000010000000100010011;
ROM[7103] <= 32'b00000000000000010010001110000011;
ROM[7104] <= 32'b00000000000000111000001100010011;
ROM[7105] <= 32'b00000000110100110000010000110011;
ROM[7106] <= 32'b00000000000001000010001110000011;
ROM[7107] <= 32'b00000000011100010010000000100011;
ROM[7108] <= 32'b00000000010000010000000100010011;
ROM[7109] <= 32'b00000010110100000000001110010011;
ROM[7110] <= 32'b00000000011100010010000000100011;
ROM[7111] <= 32'b00000000010000010000000100010011;
ROM[7112] <= 32'b11111111110000010000000100010011;
ROM[7113] <= 32'b00000000000000010010001110000011;
ROM[7114] <= 32'b11111111110000010000000100010011;
ROM[7115] <= 32'b00000000000000010010010000000011;
ROM[7116] <= 32'b00000000011101000010010010110011;
ROM[7117] <= 32'b00000000100000111010010100110011;
ROM[7118] <= 32'b00000000101001001000001110110011;
ROM[7119] <= 32'b00000000000100111000001110010011;
ROM[7120] <= 32'b00000000000100111111001110010011;
ROM[7121] <= 32'b00000000011100010010000000100011;
ROM[7122] <= 32'b00000000010000010000000100010011;
ROM[7123] <= 32'b11111111110000010000000100010011;
ROM[7124] <= 32'b00000000000000010010001110000011;
ROM[7125] <= 32'b11111111110000010000000100010011;
ROM[7126] <= 32'b00000000000000010010010000000011;
ROM[7127] <= 32'b00000000011101000111001110110011;
ROM[7128] <= 32'b00000000011100010010000000100011;
ROM[7129] <= 32'b00000000010000010000000100010011;
ROM[7130] <= 32'b11111111110000010000000100010011;
ROM[7131] <= 32'b00000000000000010010001110000011;
ROM[7132] <= 32'b00000000000000111000101001100011;
ROM[7133] <= 32'b00000000000000000111001110110111;
ROM[7134] <= 32'b11111000100000111000001110010011;
ROM[7135] <= 32'b00000000111000111000001110110011;
ROM[7136] <= 32'b00000000000000111000000011100111;
ROM[7137] <= 32'b00000101000000000000000011101111;
ROM[7138] <= 32'b00000000000000000000001110010011;
ROM[7139] <= 32'b00000000011100010010000000100011;
ROM[7140] <= 32'b00000000010000010000000100010011;
ROM[7141] <= 32'b11111111110000010000000100010011;
ROM[7142] <= 32'b00000000000000010010001110000011;
ROM[7143] <= 32'b01000000011100000000001110110011;
ROM[7144] <= 32'b00000000000100111000001110010011;
ROM[7145] <= 32'b00000000011100010010000000100011;
ROM[7146] <= 32'b00000000010000010000000100010011;
ROM[7147] <= 32'b11111111110000010000000100010011;
ROM[7148] <= 32'b00000000000000010010001110000011;
ROM[7149] <= 32'b00000000011100011010010000100011;
ROM[7150] <= 32'b00000000000100000000001110010011;
ROM[7151] <= 32'b00000000011100010010000000100011;
ROM[7152] <= 32'b00000000010000010000000100010011;
ROM[7153] <= 32'b11111111110000010000000100010011;
ROM[7154] <= 32'b00000000000000010010001110000011;
ROM[7155] <= 32'b00000000011100011010001000100011;
ROM[7156] <= 32'b00000011010000000000000011101111;
ROM[7157] <= 32'b00000000000000000000001110010011;
ROM[7158] <= 32'b00000000011100010010000000100011;
ROM[7159] <= 32'b00000000010000010000000100010011;
ROM[7160] <= 32'b11111111110000010000000100010011;
ROM[7161] <= 32'b00000000000000010010001110000011;
ROM[7162] <= 32'b00000000011100011010010000100011;
ROM[7163] <= 32'b00000000000000000000001110010011;
ROM[7164] <= 32'b00000000011100010010000000100011;
ROM[7165] <= 32'b00000000010000010000000100010011;
ROM[7166] <= 32'b11111111110000010000000100010011;
ROM[7167] <= 32'b00000000000000010010001110000011;
ROM[7168] <= 32'b00000000011100011010001000100011;
ROM[7169] <= 32'b00000000010000011010001110000011;
ROM[7170] <= 32'b00000000011100010010000000100011;
ROM[7171] <= 32'b00000000010000010000000100010011;
ROM[7172] <= 32'b00000000110100101000010000110011;
ROM[7173] <= 32'b00000000010001000010001110000011;
ROM[7174] <= 32'b00000000011100010010000000100011;
ROM[7175] <= 32'b00000000010000010000000100010011;
ROM[7176] <= 32'b11111111110000010000000100010011;
ROM[7177] <= 32'b00000000000000010010001110000011;
ROM[7178] <= 32'b11111111110000010000000100010011;
ROM[7179] <= 32'b00000000000000010010010000000011;
ROM[7180] <= 32'b00000000011101000010001110110011;
ROM[7181] <= 32'b00000000011100010010000000100011;
ROM[7182] <= 32'b00000000010000010000000100010011;
ROM[7183] <= 32'b00000000010000011010001110000011;
ROM[7184] <= 32'b00000000011100010010000000100011;
ROM[7185] <= 32'b00000000010000010000000100010011;
ROM[7186] <= 32'b00000000110100101000010000110011;
ROM[7187] <= 32'b00000000100001000010001110000011;
ROM[7188] <= 32'b00000000011100010010000000100011;
ROM[7189] <= 32'b00000000010000010000000100010011;
ROM[7190] <= 32'b11111111110000010000000100010011;
ROM[7191] <= 32'b00000000000000010010001110000011;
ROM[7192] <= 32'b11111111110000010000000100010011;
ROM[7193] <= 32'b00000000000000010010010000000011;
ROM[7194] <= 32'b00000000011101000000001110110011;
ROM[7195] <= 32'b00000000011100010010000000100011;
ROM[7196] <= 32'b00000000010000010000000100010011;
ROM[7197] <= 32'b11111111110000010000000100010011;
ROM[7198] <= 32'b00000000000000010010001110000011;
ROM[7199] <= 32'b00000000000000111000001100010011;
ROM[7200] <= 32'b00000000110100110000010000110011;
ROM[7201] <= 32'b00000000000001000010001110000011;
ROM[7202] <= 32'b00000000011100010010000000100011;
ROM[7203] <= 32'b00000000010000010000000100010011;
ROM[7204] <= 32'b00000000000000000111001110110111;
ROM[7205] <= 32'b00001101110000111000001110010011;
ROM[7206] <= 32'b00000000111000111000001110110011;
ROM[7207] <= 32'b00000000011100010010000000100011;
ROM[7208] <= 32'b00000000010000010000000100010011;
ROM[7209] <= 32'b00000000001100010010000000100011;
ROM[7210] <= 32'b00000000010000010000000100010011;
ROM[7211] <= 32'b00000000010000010010000000100011;
ROM[7212] <= 32'b00000000010000010000000100010011;
ROM[7213] <= 32'b00000000010100010010000000100011;
ROM[7214] <= 32'b00000000010000010000000100010011;
ROM[7215] <= 32'b00000000011000010010000000100011;
ROM[7216] <= 32'b00000000010000010000000100010011;
ROM[7217] <= 32'b00000001010000000000001110010011;
ROM[7218] <= 32'b00000000010000111000001110010011;
ROM[7219] <= 32'b01000000011100010000001110110011;
ROM[7220] <= 32'b00000000011100000000001000110011;
ROM[7221] <= 32'b00000000001000000000000110110011;
ROM[7222] <= 32'b00101001000000000000000011101111;
ROM[7223] <= 32'b11111111110000010000000100010011;
ROM[7224] <= 32'b00000000000000010010001110000011;
ROM[7225] <= 32'b11111111110000010000000100010011;
ROM[7226] <= 32'b00000000000000010010010000000011;
ROM[7227] <= 32'b00000000011101000111001110110011;
ROM[7228] <= 32'b00000000011100010010000000100011;
ROM[7229] <= 32'b00000000010000010000000100010011;
ROM[7230] <= 32'b11111111110000010000000100010011;
ROM[7231] <= 32'b00000000000000010010001110000011;
ROM[7232] <= 32'b01000000011100000000001110110011;
ROM[7233] <= 32'b00000000000100111000001110010011;
ROM[7234] <= 32'b00000000011100010010000000100011;
ROM[7235] <= 32'b00000000010000010000000100010011;
ROM[7236] <= 32'b11111111110000010000000100010011;
ROM[7237] <= 32'b00000000000000010010001110000011;
ROM[7238] <= 32'b00000000000000111000101001100011;
ROM[7239] <= 32'b00000000000000001000001110110111;
ROM[7240] <= 32'b11001110010000111000001110010011;
ROM[7241] <= 32'b00000000111000111000001110110011;
ROM[7242] <= 32'b00000000000000111000000011100111;
ROM[7243] <= 32'b00000000000000011010001110000011;
ROM[7244] <= 32'b00000000011100010010000000100011;
ROM[7245] <= 32'b00000000010000010000000100010011;
ROM[7246] <= 32'b00000000101000000000001110010011;
ROM[7247] <= 32'b00000000011100010010000000100011;
ROM[7248] <= 32'b00000000010000010000000100010011;
ROM[7249] <= 32'b00000000000000000111001110110111;
ROM[7250] <= 32'b00011001000000111000001110010011;
ROM[7251] <= 32'b00000000111000111000001110110011;
ROM[7252] <= 32'b00000000011100010010000000100011;
ROM[7253] <= 32'b00000000010000010000000100010011;
ROM[7254] <= 32'b00000000001100010010000000100011;
ROM[7255] <= 32'b00000000010000010000000100010011;
ROM[7256] <= 32'b00000000010000010010000000100011;
ROM[7257] <= 32'b00000000010000010000000100010011;
ROM[7258] <= 32'b00000000010100010010000000100011;
ROM[7259] <= 32'b00000000010000010000000100010011;
ROM[7260] <= 32'b00000000011000010010000000100011;
ROM[7261] <= 32'b00000000010000010000000100010011;
ROM[7262] <= 32'b00000001010000000000001110010011;
ROM[7263] <= 32'b00000000100000111000001110010011;
ROM[7264] <= 32'b01000000011100010000001110110011;
ROM[7265] <= 32'b00000000011100000000001000110011;
ROM[7266] <= 32'b00000000001000000000000110110011;
ROM[7267] <= 32'b11011011110111111010000011101111;
ROM[7268] <= 32'b00000000010000011010001110000011;
ROM[7269] <= 32'b00000000011100010010000000100011;
ROM[7270] <= 32'b00000000010000010000000100010011;
ROM[7271] <= 32'b00000000110100101000010000110011;
ROM[7272] <= 32'b00000000100001000010001110000011;
ROM[7273] <= 32'b00000000011100010010000000100011;
ROM[7274] <= 32'b00000000010000010000000100010011;
ROM[7275] <= 32'b11111111110000010000000100010011;
ROM[7276] <= 32'b00000000000000010010001110000011;
ROM[7277] <= 32'b11111111110000010000000100010011;
ROM[7278] <= 32'b00000000000000010010010000000011;
ROM[7279] <= 32'b00000000011101000000001110110011;
ROM[7280] <= 32'b00000000011100010010000000100011;
ROM[7281] <= 32'b00000000010000010000000100010011;
ROM[7282] <= 32'b11111111110000010000000100010011;
ROM[7283] <= 32'b00000000000000010010001110000011;
ROM[7284] <= 32'b00000000000000111000001100010011;
ROM[7285] <= 32'b00000000110100110000010000110011;
ROM[7286] <= 32'b00000000000001000010001110000011;
ROM[7287] <= 32'b00000000011100010010000000100011;
ROM[7288] <= 32'b00000000010000010000000100010011;
ROM[7289] <= 32'b00000000000000000111001110110111;
ROM[7290] <= 32'b00100011000000111000001110010011;
ROM[7291] <= 32'b00000000111000111000001110110011;
ROM[7292] <= 32'b00000000011100010010000000100011;
ROM[7293] <= 32'b00000000010000010000000100010011;
ROM[7294] <= 32'b00000000001100010010000000100011;
ROM[7295] <= 32'b00000000010000010000000100010011;
ROM[7296] <= 32'b00000000010000010010000000100011;
ROM[7297] <= 32'b00000000010000010000000100010011;
ROM[7298] <= 32'b00000000010100010010000000100011;
ROM[7299] <= 32'b00000000010000010000000100010011;
ROM[7300] <= 32'b00000000011000010010000000100011;
ROM[7301] <= 32'b00000000010000010000000100010011;
ROM[7302] <= 32'b00000001010000000000001110010011;
ROM[7303] <= 32'b00000000010000111000001110010011;
ROM[7304] <= 32'b01000000011100010000001110110011;
ROM[7305] <= 32'b00000000011100000000001000110011;
ROM[7306] <= 32'b00000000001000000000000110110011;
ROM[7307] <= 32'b00100010100000000000000011101111;
ROM[7308] <= 32'b11111111110000010000000100010011;
ROM[7309] <= 32'b00000000000000010010001110000011;
ROM[7310] <= 32'b11111111110000010000000100010011;
ROM[7311] <= 32'b00000000000000010010010000000011;
ROM[7312] <= 32'b00000000011101000000001110110011;
ROM[7313] <= 32'b00000000011100010010000000100011;
ROM[7314] <= 32'b00000000010000010000000100010011;
ROM[7315] <= 32'b11111111110000010000000100010011;
ROM[7316] <= 32'b00000000000000010010001110000011;
ROM[7317] <= 32'b00000000011100011010000000100011;
ROM[7318] <= 32'b00000000010000011010001110000011;
ROM[7319] <= 32'b00000000011100010010000000100011;
ROM[7320] <= 32'b00000000010000010000000100010011;
ROM[7321] <= 32'b00000000000100000000001110010011;
ROM[7322] <= 32'b00000000011100010010000000100011;
ROM[7323] <= 32'b00000000010000010000000100010011;
ROM[7324] <= 32'b11111111110000010000000100010011;
ROM[7325] <= 32'b00000000000000010010001110000011;
ROM[7326] <= 32'b11111111110000010000000100010011;
ROM[7327] <= 32'b00000000000000010010010000000011;
ROM[7328] <= 32'b00000000011101000000001110110011;
ROM[7329] <= 32'b00000000011100010010000000100011;
ROM[7330] <= 32'b00000000010000010000000100010011;
ROM[7331] <= 32'b11111111110000010000000100010011;
ROM[7332] <= 32'b00000000000000010010001110000011;
ROM[7333] <= 32'b00000000011100011010001000100011;
ROM[7334] <= 32'b00011111000100000000000011101111;
ROM[7335] <= 32'b00000000100000011010001110000011;
ROM[7336] <= 32'b00000000011100010010000000100011;
ROM[7337] <= 32'b00000000010000010000000100010011;
ROM[7338] <= 32'b11111111110000010000000100010011;
ROM[7339] <= 32'b00000000000000010010001110000011;
ROM[7340] <= 32'b00000000000000111000101001100011;
ROM[7341] <= 32'b00000000000000000111001110110111;
ROM[7342] <= 32'b00101100100000111000001110010011;
ROM[7343] <= 32'b00000000111000111000001110110011;
ROM[7344] <= 32'b00000000000000111000000011100111;
ROM[7345] <= 32'b00000110000000000000000011101111;
ROM[7346] <= 32'b00000000000000011010001110000011;
ROM[7347] <= 32'b00000000011100010010000000100011;
ROM[7348] <= 32'b00000000010000010000000100010011;
ROM[7349] <= 32'b11111111110000010000000100010011;
ROM[7350] <= 32'b00000000000000010010001110000011;
ROM[7351] <= 32'b01000000011100000000001110110011;
ROM[7352] <= 32'b00000000011100010010000000100011;
ROM[7353] <= 32'b00000000010000010000000100010011;
ROM[7354] <= 32'b00000001010000000000001110010011;
ROM[7355] <= 32'b01000000011100011000001110110011;
ROM[7356] <= 32'b00000000000000111010000010000011;
ROM[7357] <= 32'b11111111110000010000000100010011;
ROM[7358] <= 32'b00000000000000010010001110000011;
ROM[7359] <= 32'b00000000011100100010000000100011;
ROM[7360] <= 32'b00000000010000100000000100010011;
ROM[7361] <= 32'b00000001010000000000001110010011;
ROM[7362] <= 32'b01000000011100011000001110110011;
ROM[7363] <= 32'b00000000010000111010000110000011;
ROM[7364] <= 32'b00000000100000111010001000000011;
ROM[7365] <= 32'b00000000110000111010001010000011;
ROM[7366] <= 32'b00000001000000111010001100000011;
ROM[7367] <= 32'b00000000000000001000000011100111;
ROM[7368] <= 32'b00000100100000000000000011101111;
ROM[7369] <= 32'b00000000000000011010001110000011;
ROM[7370] <= 32'b00000000011100010010000000100011;
ROM[7371] <= 32'b00000000010000010000000100010011;
ROM[7372] <= 32'b00000001010000000000001110010011;
ROM[7373] <= 32'b01000000011100011000001110110011;
ROM[7374] <= 32'b00000000000000111010000010000011;
ROM[7375] <= 32'b11111111110000010000000100010011;
ROM[7376] <= 32'b00000000000000010010001110000011;
ROM[7377] <= 32'b00000000011100100010000000100011;
ROM[7378] <= 32'b00000000010000100000000100010011;
ROM[7379] <= 32'b00000001010000000000001110010011;
ROM[7380] <= 32'b01000000011100011000001110110011;
ROM[7381] <= 32'b00000000010000111010000110000011;
ROM[7382] <= 32'b00000000100000111010001000000011;
ROM[7383] <= 32'b00000000110000111010001010000011;
ROM[7384] <= 32'b00000001000000111010001100000011;
ROM[7385] <= 32'b00000000000000001000000011100111;
ROM[7386] <= 32'b00000000000000100010001110000011;
ROM[7387] <= 32'b00000000011100010010000000100011;
ROM[7388] <= 32'b00000000010000010000000100010011;
ROM[7389] <= 32'b00000011000000000000001110010011;
ROM[7390] <= 32'b00000000011100010010000000100011;
ROM[7391] <= 32'b00000000010000010000000100010011;
ROM[7392] <= 32'b11111111110000010000000100010011;
ROM[7393] <= 32'b00000000000000010010001110000011;
ROM[7394] <= 32'b11111111110000010000000100010011;
ROM[7395] <= 32'b00000000000000010010010000000011;
ROM[7396] <= 32'b00000000011101000010001110110011;
ROM[7397] <= 32'b00000000011100010010000000100011;
ROM[7398] <= 32'b00000000010000010000000100010011;
ROM[7399] <= 32'b11111111110000010000000100010011;
ROM[7400] <= 32'b00000000000000010010001110000011;
ROM[7401] <= 32'b01000000011100000000001110110011;
ROM[7402] <= 32'b00000000000100111000001110010011;
ROM[7403] <= 32'b00000000011100010010000000100011;
ROM[7404] <= 32'b00000000010000010000000100010011;
ROM[7405] <= 32'b00000000000000100010001110000011;
ROM[7406] <= 32'b00000000011100010010000000100011;
ROM[7407] <= 32'b00000000010000010000000100010011;
ROM[7408] <= 32'b00000011100100000000001110010011;
ROM[7409] <= 32'b00000000011100010010000000100011;
ROM[7410] <= 32'b00000000010000010000000100010011;
ROM[7411] <= 32'b11111111110000010000000100010011;
ROM[7412] <= 32'b00000000000000010010001110000011;
ROM[7413] <= 32'b11111111110000010000000100010011;
ROM[7414] <= 32'b00000000000000010010010000000011;
ROM[7415] <= 32'b00000000100000111010001110110011;
ROM[7416] <= 32'b00000000011100010010000000100011;
ROM[7417] <= 32'b00000000010000010000000100010011;
ROM[7418] <= 32'b11111111110000010000000100010011;
ROM[7419] <= 32'b00000000000000010010001110000011;
ROM[7420] <= 32'b01000000011100000000001110110011;
ROM[7421] <= 32'b00000000000100111000001110010011;
ROM[7422] <= 32'b00000000011100010010000000100011;
ROM[7423] <= 32'b00000000010000010000000100010011;
ROM[7424] <= 32'b11111111110000010000000100010011;
ROM[7425] <= 32'b00000000000000010010001110000011;
ROM[7426] <= 32'b11111111110000010000000100010011;
ROM[7427] <= 32'b00000000000000010010010000000011;
ROM[7428] <= 32'b00000000011101000111001110110011;
ROM[7429] <= 32'b00000000011100010010000000100011;
ROM[7430] <= 32'b00000000010000010000000100010011;
ROM[7431] <= 32'b00000001010000000000001110010011;
ROM[7432] <= 32'b01000000011100011000001110110011;
ROM[7433] <= 32'b00000000000000111010000010000011;
ROM[7434] <= 32'b11111111110000010000000100010011;
ROM[7435] <= 32'b00000000000000010010001110000011;
ROM[7436] <= 32'b00000000011100100010000000100011;
ROM[7437] <= 32'b00000000010000100000000100010011;
ROM[7438] <= 32'b00000001010000000000001110010011;
ROM[7439] <= 32'b01000000011100011000001110110011;
ROM[7440] <= 32'b00000000010000111010000110000011;
ROM[7441] <= 32'b00000000100000111010001000000011;
ROM[7442] <= 32'b00000000110000111010001010000011;
ROM[7443] <= 32'b00000001000000111010001100000011;
ROM[7444] <= 32'b00000000000000001000000011100111;
ROM[7445] <= 32'b00000000000000100010001110000011;
ROM[7446] <= 32'b00000000011100010010000000100011;
ROM[7447] <= 32'b00000000010000010000000100010011;
ROM[7448] <= 32'b00000011000000000000001110010011;
ROM[7449] <= 32'b00000000011100010010000000100011;
ROM[7450] <= 32'b00000000010000010000000100010011;
ROM[7451] <= 32'b11111111110000010000000100010011;
ROM[7452] <= 32'b00000000000000010010001110000011;
ROM[7453] <= 32'b11111111110000010000000100010011;
ROM[7454] <= 32'b00000000000000010010010000000011;
ROM[7455] <= 32'b01000000011101000000001110110011;
ROM[7456] <= 32'b00000000011100010010000000100011;
ROM[7457] <= 32'b00000000010000010000000100010011;
ROM[7458] <= 32'b00000001010000000000001110010011;
ROM[7459] <= 32'b01000000011100011000001110110011;
ROM[7460] <= 32'b00000000000000111010000010000011;
ROM[7461] <= 32'b11111111110000010000000100010011;
ROM[7462] <= 32'b00000000000000010010001110000011;
ROM[7463] <= 32'b00000000011100100010000000100011;
ROM[7464] <= 32'b00000000010000100000000100010011;
ROM[7465] <= 32'b00000001010000000000001110010011;
ROM[7466] <= 32'b01000000011100011000001110110011;
ROM[7467] <= 32'b00000000010000111010000110000011;
ROM[7468] <= 32'b00000000100000111010001000000011;
ROM[7469] <= 32'b00000000110000111010001010000011;
ROM[7470] <= 32'b00000001000000111010001100000011;
ROM[7471] <= 32'b00000000000000001000000011100111;
ROM[7472] <= 32'b00000000000000100010001110000011;
ROM[7473] <= 32'b00000000011100010010000000100011;
ROM[7474] <= 32'b00000000010000010000000100010011;
ROM[7475] <= 32'b00000011000000000000001110010011;
ROM[7476] <= 32'b00000000011100010010000000100011;
ROM[7477] <= 32'b00000000010000010000000100010011;
ROM[7478] <= 32'b11111111110000010000000100010011;
ROM[7479] <= 32'b00000000000000010010001110000011;
ROM[7480] <= 32'b11111111110000010000000100010011;
ROM[7481] <= 32'b00000000000000010010010000000011;
ROM[7482] <= 32'b00000000011101000000001110110011;
ROM[7483] <= 32'b00000000011100010010000000100011;
ROM[7484] <= 32'b00000000010000010000000100010011;
ROM[7485] <= 32'b00000001010000000000001110010011;
ROM[7486] <= 32'b01000000011100011000001110110011;
ROM[7487] <= 32'b00000000000000111010000010000011;
ROM[7488] <= 32'b11111111110000010000000100010011;
ROM[7489] <= 32'b00000000000000010010001110000011;
ROM[7490] <= 32'b00000000011100100010000000100011;
ROM[7491] <= 32'b00000000010000100000000100010011;
ROM[7492] <= 32'b00000001010000000000001110010011;
ROM[7493] <= 32'b01000000011100011000001110110011;
ROM[7494] <= 32'b00000000010000111010000110000011;
ROM[7495] <= 32'b00000000100000111010001000000011;
ROM[7496] <= 32'b00000000110000111010001010000011;
ROM[7497] <= 32'b00000001000000111010001100000011;
ROM[7498] <= 32'b00000000000000001000000011100111;
ROM[7499] <= 32'b00000000000000100010001110000011;
ROM[7500] <= 32'b00000000011100010010000000100011;
ROM[7501] <= 32'b00000000010000010000000100010011;
ROM[7502] <= 32'b11111111110000010000000100010011;
ROM[7503] <= 32'b00000000000000010010001110000011;
ROM[7504] <= 32'b00000000000000111000001010010011;
ROM[7505] <= 32'b00000000000000000000001110010011;
ROM[7506] <= 32'b00000000011100010010000000100011;
ROM[7507] <= 32'b00000000010000010000000100010011;
ROM[7508] <= 32'b11111111110000010000000100010011;
ROM[7509] <= 32'b00000000000000010010001110000011;
ROM[7510] <= 32'b00000000110100101000010000110011;
ROM[7511] <= 32'b00000000011101000010001000100011;
ROM[7512] <= 32'b00000000010000100010001110000011;
ROM[7513] <= 32'b00000000011100010010000000100011;
ROM[7514] <= 32'b00000000010000010000000100010011;
ROM[7515] <= 32'b00000000000000000000001110010011;
ROM[7516] <= 32'b00000000011100010010000000100011;
ROM[7517] <= 32'b00000000010000010000000100010011;
ROM[7518] <= 32'b11111111110000010000000100010011;
ROM[7519] <= 32'b00000000000000010010001110000011;
ROM[7520] <= 32'b11111111110000010000000100010011;
ROM[7521] <= 32'b00000000000000010010010000000011;
ROM[7522] <= 32'b00000000011101000010001110110011;
ROM[7523] <= 32'b00000000011100010010000000100011;
ROM[7524] <= 32'b00000000010000010000000100010011;
ROM[7525] <= 32'b11111111110000010000000100010011;
ROM[7526] <= 32'b00000000000000010010001110000011;
ROM[7527] <= 32'b00000000000000111000101001100011;
ROM[7528] <= 32'b00000000000000000111001110110111;
ROM[7529] <= 32'b01011011010000111000001110010011;
ROM[7530] <= 32'b00000000111000111000001110110011;
ROM[7531] <= 32'b00000000000000111000000011100111;
ROM[7532] <= 32'b00001010000000000000000011101111;
ROM[7533] <= 32'b00000000010000100010001110000011;
ROM[7534] <= 32'b00000000011100010010000000100011;
ROM[7535] <= 32'b00000000010000010000000100010011;
ROM[7536] <= 32'b11111111110000010000000100010011;
ROM[7537] <= 32'b00000000000000010010001110000011;
ROM[7538] <= 32'b01000000011100000000001110110011;
ROM[7539] <= 32'b00000000011100010010000000100011;
ROM[7540] <= 32'b00000000010000010000000100010011;
ROM[7541] <= 32'b11111111110000010000000100010011;
ROM[7542] <= 32'b00000000000000010010001110000011;
ROM[7543] <= 32'b00000000011100100010001000100011;
ROM[7544] <= 32'b00000000000000010010001010000011;
ROM[7545] <= 32'b00000000010000010000000100010011;
ROM[7546] <= 32'b00000010110100000000001110010011;
ROM[7547] <= 32'b00000000011100010010000000100011;
ROM[7548] <= 32'b00000000010000010000000100010011;
ROM[7549] <= 32'b00000000000000000111001110110111;
ROM[7550] <= 32'b01100100000000111000001110010011;
ROM[7551] <= 32'b00000000111000111000001110110011;
ROM[7552] <= 32'b00000000011100010010000000100011;
ROM[7553] <= 32'b00000000010000010000000100010011;
ROM[7554] <= 32'b00000000001100010010000000100011;
ROM[7555] <= 32'b00000000010000010000000100010011;
ROM[7556] <= 32'b00000000010000010010000000100011;
ROM[7557] <= 32'b00000000010000010000000100010011;
ROM[7558] <= 32'b00000000010100010010000000100011;
ROM[7559] <= 32'b00000000010000010000000100010011;
ROM[7560] <= 32'b00000000011000010010000000100011;
ROM[7561] <= 32'b00000000010000010000000100010011;
ROM[7562] <= 32'b00000001010000000000001110010011;
ROM[7563] <= 32'b00000000100000111000001110010011;
ROM[7564] <= 32'b01000000011100010000001110110011;
ROM[7565] <= 32'b00000000011100000000001000110011;
ROM[7566] <= 32'b00000000001000000000000110110011;
ROM[7567] <= 32'b11011000000011111111000011101111;
ROM[7568] <= 32'b11111111110000010000000100010011;
ROM[7569] <= 32'b00000000000000010010001110000011;
ROM[7570] <= 32'b00000000011101100010000000100011;
ROM[7571] <= 32'b00000000010000000000000011101111;
ROM[7572] <= 32'b00000000000000010010001010000011;
ROM[7573] <= 32'b00000000010000010000000100010011;
ROM[7574] <= 32'b00000000010000100010001110000011;
ROM[7575] <= 32'b00000000011100010010000000100011;
ROM[7576] <= 32'b00000000010000010000000100010011;
ROM[7577] <= 32'b00000000000000000111001110110111;
ROM[7578] <= 32'b01101011000000111000001110010011;
ROM[7579] <= 32'b00000000111000111000001110110011;
ROM[7580] <= 32'b00000000011100010010000000100011;
ROM[7581] <= 32'b00000000010000010000000100010011;
ROM[7582] <= 32'b00000000001100010010000000100011;
ROM[7583] <= 32'b00000000010000010000000100010011;
ROM[7584] <= 32'b00000000010000010010000000100011;
ROM[7585] <= 32'b00000000010000010000000100010011;
ROM[7586] <= 32'b00000000010100010010000000100011;
ROM[7587] <= 32'b00000000010000010000000100010011;
ROM[7588] <= 32'b00000000011000010010000000100011;
ROM[7589] <= 32'b00000000010000010000000100010011;
ROM[7590] <= 32'b00000001010000000000001110010011;
ROM[7591] <= 32'b00000000100000111000001110010011;
ROM[7592] <= 32'b01000000011100010000001110110011;
ROM[7593] <= 32'b00000000011100000000001000110011;
ROM[7594] <= 32'b00000000001000000000000110110011;
ROM[7595] <= 32'b00000101010000000000000011101111;
ROM[7596] <= 32'b11111111110000010000000100010011;
ROM[7597] <= 32'b00000000000000010010001110000011;
ROM[7598] <= 32'b00000000011101100010000000100011;
ROM[7599] <= 32'b00000000000000000000001110010011;
ROM[7600] <= 32'b00000000011100010010000000100011;
ROM[7601] <= 32'b00000000010000010000000100010011;
ROM[7602] <= 32'b00000001010000000000001110010011;
ROM[7603] <= 32'b01000000011100011000001110110011;
ROM[7604] <= 32'b00000000000000111010000010000011;
ROM[7605] <= 32'b11111111110000010000000100010011;
ROM[7606] <= 32'b00000000000000010010001110000011;
ROM[7607] <= 32'b00000000011100100010000000100011;
ROM[7608] <= 32'b00000000010000100000000100010011;
ROM[7609] <= 32'b00000001010000000000001110010011;
ROM[7610] <= 32'b01000000011100011000001110110011;
ROM[7611] <= 32'b00000000010000111010000110000011;
ROM[7612] <= 32'b00000000100000111010001000000011;
ROM[7613] <= 32'b00000000110000111010001010000011;
ROM[7614] <= 32'b00000001000000111010001100000011;
ROM[7615] <= 32'b00000000000000001000000011100111;
ROM[7616] <= 32'b00000000000000010010000000100011;
ROM[7617] <= 32'b00000000010000010000000100010011;
ROM[7618] <= 32'b00000000000000100010001110000011;
ROM[7619] <= 32'b00000000011100010010000000100011;
ROM[7620] <= 32'b00000000010000010000000100010011;
ROM[7621] <= 32'b11111111110000010000000100010011;
ROM[7622] <= 32'b00000000000000010010001110000011;
ROM[7623] <= 32'b00000000000000111000001010010011;
ROM[7624] <= 32'b00000000010000100010001110000011;
ROM[7625] <= 32'b00000000011100010010000000100011;
ROM[7626] <= 32'b00000000010000010000000100010011;
ROM[7627] <= 32'b00000000101000000000001110010011;
ROM[7628] <= 32'b00000000011100010010000000100011;
ROM[7629] <= 32'b00000000010000010000000100010011;
ROM[7630] <= 32'b11111111110000010000000100010011;
ROM[7631] <= 32'b00000000000000010010001110000011;
ROM[7632] <= 32'b11111111110000010000000100010011;
ROM[7633] <= 32'b00000000000000010010010000000011;
ROM[7634] <= 32'b00000000011101000010001110110011;
ROM[7635] <= 32'b00000000011100010010000000100011;
ROM[7636] <= 32'b00000000010000010000000100010011;
ROM[7637] <= 32'b11111111110000010000000100010011;
ROM[7638] <= 32'b00000000000000010010001110000011;
ROM[7639] <= 32'b00000000000000111000101001100011;
ROM[7640] <= 32'b00000000000000000111001110110111;
ROM[7641] <= 32'b01110111010000111000001110010011;
ROM[7642] <= 32'b00000000111000111000001110110011;
ROM[7643] <= 32'b00000000000000111000000011100111;
ROM[7644] <= 32'b00001100000000000000000011101111;
ROM[7645] <= 32'b00000000000000010010001010000011;
ROM[7646] <= 32'b00000000010000010000000100010011;
ROM[7647] <= 32'b00000000010000100010001110000011;
ROM[7648] <= 32'b00000000011100010010000000100011;
ROM[7649] <= 32'b00000000010000010000000100010011;
ROM[7650] <= 32'b00000000000000000111001110110111;
ROM[7651] <= 32'b01111101010000111000001110010011;
ROM[7652] <= 32'b00000000111000111000001110110011;
ROM[7653] <= 32'b00000000011100010010000000100011;
ROM[7654] <= 32'b00000000010000010000000100010011;
ROM[7655] <= 32'b00000000001100010010000000100011;
ROM[7656] <= 32'b00000000010000010000000100010011;
ROM[7657] <= 32'b00000000010000010010000000100011;
ROM[7658] <= 32'b00000000010000010000000100010011;
ROM[7659] <= 32'b00000000010100010010000000100011;
ROM[7660] <= 32'b00000000010000010000000100010011;
ROM[7661] <= 32'b00000000011000010010000000100011;
ROM[7662] <= 32'b00000000010000010000000100010011;
ROM[7663] <= 32'b00000001010000000000001110010011;
ROM[7664] <= 32'b00000000010000111000001110010011;
ROM[7665] <= 32'b01000000011100010000001110110011;
ROM[7666] <= 32'b00000000011100000000001000110011;
ROM[7667] <= 32'b00000000001000000000000110110011;
ROM[7668] <= 32'b11001111000111111111000011101111;
ROM[7669] <= 32'b00000000000000001000001110110111;
ROM[7670] <= 32'b10000010000000111000001110010011;
ROM[7671] <= 32'b00000000111000111000001110110011;
ROM[7672] <= 32'b00000000011100010010000000100011;
ROM[7673] <= 32'b00000000010000010000000100010011;
ROM[7674] <= 32'b00000000001100010010000000100011;
ROM[7675] <= 32'b00000000010000010000000100010011;
ROM[7676] <= 32'b00000000010000010010000000100011;
ROM[7677] <= 32'b00000000010000010000000100010011;
ROM[7678] <= 32'b00000000010100010010000000100011;
ROM[7679] <= 32'b00000000010000010000000100010011;
ROM[7680] <= 32'b00000000011000010010000000100011;
ROM[7681] <= 32'b00000000010000010000000100010011;
ROM[7682] <= 32'b00000001010000000000001110010011;
ROM[7683] <= 32'b00000000100000111000001110010011;
ROM[7684] <= 32'b01000000011100010000001110110011;
ROM[7685] <= 32'b00000000011100000000001000110011;
ROM[7686] <= 32'b00000000001000000000000110110011;
ROM[7687] <= 32'b10111010000011111111000011101111;
ROM[7688] <= 32'b11111111110000010000000100010011;
ROM[7689] <= 32'b00000000000000010010001110000011;
ROM[7690] <= 32'b00000000011101100010000000100011;
ROM[7691] <= 32'b00100001100000000000000011101111;
ROM[7692] <= 32'b00000000010000100010001110000011;
ROM[7693] <= 32'b00000000011100010010000000100011;
ROM[7694] <= 32'b00000000010000010000000100010011;
ROM[7695] <= 32'b00000000101000000000001110010011;
ROM[7696] <= 32'b00000000011100010010000000100011;
ROM[7697] <= 32'b00000000010000010000000100010011;
ROM[7698] <= 32'b00000000000000001000001110110111;
ROM[7699] <= 32'b10001001010000111000001110010011;
ROM[7700] <= 32'b00000000111000111000001110110011;
ROM[7701] <= 32'b00000000011100010010000000100011;
ROM[7702] <= 32'b00000000010000010000000100010011;
ROM[7703] <= 32'b00000000001100010010000000100011;
ROM[7704] <= 32'b00000000010000010000000100010011;
ROM[7705] <= 32'b00000000010000010010000000100011;
ROM[7706] <= 32'b00000000010000010000000100010011;
ROM[7707] <= 32'b00000000010100010010000000100011;
ROM[7708] <= 32'b00000000010000010000000100010011;
ROM[7709] <= 32'b00000000011000010010000000100011;
ROM[7710] <= 32'b00000000010000010000000100010011;
ROM[7711] <= 32'b00000001010000000000001110010011;
ROM[7712] <= 32'b00000000100000111000001110010011;
ROM[7713] <= 32'b01000000011100010000001110110011;
ROM[7714] <= 32'b00000000011100000000001000110011;
ROM[7715] <= 32'b00000000001000000000000110110011;
ROM[7716] <= 32'b10100011110111111010000011101111;
ROM[7717] <= 32'b11111111110000010000000100010011;
ROM[7718] <= 32'b00000000000000010010001110000011;
ROM[7719] <= 32'b00000000011100011010000000100011;
ROM[7720] <= 32'b00000000000000010010001010000011;
ROM[7721] <= 32'b00000000010000010000000100010011;
ROM[7722] <= 32'b00000000000000011010001110000011;
ROM[7723] <= 32'b00000000011100010010000000100011;
ROM[7724] <= 32'b00000000010000010000000100010011;
ROM[7725] <= 32'b00000000000000001000001110110111;
ROM[7726] <= 32'b10010000000000111000001110010011;
ROM[7727] <= 32'b00000000111000111000001110110011;
ROM[7728] <= 32'b00000000011100010010000000100011;
ROM[7729] <= 32'b00000000010000010000000100010011;
ROM[7730] <= 32'b00000000001100010010000000100011;
ROM[7731] <= 32'b00000000010000010000000100010011;
ROM[7732] <= 32'b00000000010000010010000000100011;
ROM[7733] <= 32'b00000000010000010000000100010011;
ROM[7734] <= 32'b00000000010100010010000000100011;
ROM[7735] <= 32'b00000000010000010000000100010011;
ROM[7736] <= 32'b00000000011000010010000000100011;
ROM[7737] <= 32'b00000000010000010000000100010011;
ROM[7738] <= 32'b00000001010000000000001110010011;
ROM[7739] <= 32'b00000000100000111000001110010011;
ROM[7740] <= 32'b01000000011100010000001110110011;
ROM[7741] <= 32'b00000000011100000000001000110011;
ROM[7742] <= 32'b00000000001000000000000110110011;
ROM[7743] <= 32'b11100000010111111111000011101111;
ROM[7744] <= 32'b11111111110000010000000100010011;
ROM[7745] <= 32'b00000000000000010010001110000011;
ROM[7746] <= 32'b00000000011101100010000000100011;
ROM[7747] <= 32'b00000000000000010010001010000011;
ROM[7748] <= 32'b00000000010000010000000100010011;
ROM[7749] <= 32'b00000000010000100010001110000011;
ROM[7750] <= 32'b00000000011100010010000000100011;
ROM[7751] <= 32'b00000000010000010000000100010011;
ROM[7752] <= 32'b00000000000000011010001110000011;
ROM[7753] <= 32'b00000000011100010010000000100011;
ROM[7754] <= 32'b00000000010000010000000100010011;
ROM[7755] <= 32'b00000000101000000000001110010011;
ROM[7756] <= 32'b00000000011100010010000000100011;
ROM[7757] <= 32'b00000000010000010000000100010011;
ROM[7758] <= 32'b00000000000000001000001110110111;
ROM[7759] <= 32'b10011000010000111000001110010011;
ROM[7760] <= 32'b00000000111000111000001110110011;
ROM[7761] <= 32'b00000000011100010010000000100011;
ROM[7762] <= 32'b00000000010000010000000100010011;
ROM[7763] <= 32'b00000000001100010010000000100011;
ROM[7764] <= 32'b00000000010000010000000100010011;
ROM[7765] <= 32'b00000000010000010010000000100011;
ROM[7766] <= 32'b00000000010000010000000100010011;
ROM[7767] <= 32'b00000000010100010010000000100011;
ROM[7768] <= 32'b00000000010000010000000100010011;
ROM[7769] <= 32'b00000000011000010010000000100011;
ROM[7770] <= 32'b00000000010000010000000100010011;
ROM[7771] <= 32'b00000001010000000000001110010011;
ROM[7772] <= 32'b00000000100000111000001110010011;
ROM[7773] <= 32'b01000000011100010000001110110011;
ROM[7774] <= 32'b00000000011100000000001000110011;
ROM[7775] <= 32'b00000000001000000000000110110011;
ROM[7776] <= 32'b11011100100011111010000011101111;
ROM[7777] <= 32'b11111111110000010000000100010011;
ROM[7778] <= 32'b00000000000000010010001110000011;
ROM[7779] <= 32'b11111111110000010000000100010011;
ROM[7780] <= 32'b00000000000000010010010000000011;
ROM[7781] <= 32'b01000000011101000000001110110011;
ROM[7782] <= 32'b00000000011100010010000000100011;
ROM[7783] <= 32'b00000000010000010000000100010011;
ROM[7784] <= 32'b00000000000000001000001110110111;
ROM[7785] <= 32'b10011110110000111000001110010011;
ROM[7786] <= 32'b00000000111000111000001110110011;
ROM[7787] <= 32'b00000000011100010010000000100011;
ROM[7788] <= 32'b00000000010000010000000100010011;
ROM[7789] <= 32'b00000000001100010010000000100011;
ROM[7790] <= 32'b00000000010000010000000100010011;
ROM[7791] <= 32'b00000000010000010010000000100011;
ROM[7792] <= 32'b00000000010000010000000100010011;
ROM[7793] <= 32'b00000000010100010010000000100011;
ROM[7794] <= 32'b00000000010000010000000100010011;
ROM[7795] <= 32'b00000000011000010010000000100011;
ROM[7796] <= 32'b00000000010000010000000100010011;
ROM[7797] <= 32'b00000001010000000000001110010011;
ROM[7798] <= 32'b00000000010000111000001110010011;
ROM[7799] <= 32'b01000000011100010000001110110011;
ROM[7800] <= 32'b00000000011100000000001000110011;
ROM[7801] <= 32'b00000000001000000000000110110011;
ROM[7802] <= 32'b10101101100111111111000011101111;
ROM[7803] <= 32'b00000000000000001000001110110111;
ROM[7804] <= 32'b10100011100000111000001110010011;
ROM[7805] <= 32'b00000000111000111000001110110011;
ROM[7806] <= 32'b00000000011100010010000000100011;
ROM[7807] <= 32'b00000000010000010000000100010011;
ROM[7808] <= 32'b00000000001100010010000000100011;
ROM[7809] <= 32'b00000000010000010000000100010011;
ROM[7810] <= 32'b00000000010000010010000000100011;
ROM[7811] <= 32'b00000000010000010000000100010011;
ROM[7812] <= 32'b00000000010100010010000000100011;
ROM[7813] <= 32'b00000000010000010000000100010011;
ROM[7814] <= 32'b00000000011000010010000000100011;
ROM[7815] <= 32'b00000000010000010000000100010011;
ROM[7816] <= 32'b00000001010000000000001110010011;
ROM[7817] <= 32'b00000000100000111000001110010011;
ROM[7818] <= 32'b01000000011100010000001110110011;
ROM[7819] <= 32'b00000000011100000000001000110011;
ROM[7820] <= 32'b00000000001000000000000110110011;
ROM[7821] <= 32'b10011000100011111111000011101111;
ROM[7822] <= 32'b11111111110000010000000100010011;
ROM[7823] <= 32'b00000000000000010010001110000011;
ROM[7824] <= 32'b00000000011101100010000000100011;
ROM[7825] <= 32'b00000000000000000000001110010011;
ROM[7826] <= 32'b00000000011100010010000000100011;
ROM[7827] <= 32'b00000000010000010000000100010011;
ROM[7828] <= 32'b00000001010000000000001110010011;
ROM[7829] <= 32'b01000000011100011000001110110011;
ROM[7830] <= 32'b00000000000000111010000010000011;
ROM[7831] <= 32'b11111111110000010000000100010011;
ROM[7832] <= 32'b00000000000000010010001110000011;
ROM[7833] <= 32'b00000000011100100010000000100011;
ROM[7834] <= 32'b00000000010000100000000100010011;
ROM[7835] <= 32'b00000001010000000000001110010011;
ROM[7836] <= 32'b01000000011100011000001110110011;
ROM[7837] <= 32'b00000000010000111010000110000011;
ROM[7838] <= 32'b00000000100000111010001000000011;
ROM[7839] <= 32'b00000000110000111010001010000011;
ROM[7840] <= 32'b00000001000000111010001100000011;
ROM[7841] <= 32'b00000000000000001000000011100111;
ROM[7842] <= 32'b00001000000000000000001110010011;
ROM[7843] <= 32'b00000000011100010010000000100011;
ROM[7844] <= 32'b00000000010000010000000100010011;
ROM[7845] <= 32'b00000001010000000000001110010011;
ROM[7846] <= 32'b01000000011100011000001110110011;
ROM[7847] <= 32'b00000000000000111010000010000011;
ROM[7848] <= 32'b11111111110000010000000100010011;
ROM[7849] <= 32'b00000000000000010010001110000011;
ROM[7850] <= 32'b00000000011100100010000000100011;
ROM[7851] <= 32'b00000000010000100000000100010011;
ROM[7852] <= 32'b00000001010000000000001110010011;
ROM[7853] <= 32'b01000000011100011000001110110011;
ROM[7854] <= 32'b00000000010000111010000110000011;
ROM[7855] <= 32'b00000000100000111010001000000011;
ROM[7856] <= 32'b00000000110000111010001010000011;
ROM[7857] <= 32'b00000001000000111010001100000011;
ROM[7858] <= 32'b00000000000000001000000011100111;
ROM[7859] <= 32'b00001000000100000000001110010011;
ROM[7860] <= 32'b00000000011100010010000000100011;
ROM[7861] <= 32'b00000000010000010000000100010011;
ROM[7862] <= 32'b00000001010000000000001110010011;
ROM[7863] <= 32'b01000000011100011000001110110011;
ROM[7864] <= 32'b00000000000000111010000010000011;
ROM[7865] <= 32'b11111111110000010000000100010011;
ROM[7866] <= 32'b00000000000000010010001110000011;
ROM[7867] <= 32'b00000000011100100010000000100011;
ROM[7868] <= 32'b00000000010000100000000100010011;
ROM[7869] <= 32'b00000001010000000000001110010011;
ROM[7870] <= 32'b01000000011100011000001110110011;
ROM[7871] <= 32'b00000000010000111010000110000011;
ROM[7872] <= 32'b00000000100000111010001000000011;
ROM[7873] <= 32'b00000000110000111010001010000011;
ROM[7874] <= 32'b00000001000000111010001100000011;
ROM[7875] <= 32'b00000000000000001000000011100111;
ROM[7876] <= 32'b00000010001000000000001110010011;
ROM[7877] <= 32'b00000000011100010010000000100011;
ROM[7878] <= 32'b00000000010000010000000100010011;
ROM[7879] <= 32'b00000001010000000000001110010011;
ROM[7880] <= 32'b01000000011100011000001110110011;
ROM[7881] <= 32'b00000000000000111010000010000011;
ROM[7882] <= 32'b11111111110000010000000100010011;
ROM[7883] <= 32'b00000000000000010010001110000011;
ROM[7884] <= 32'b00000000011100100010000000100011;
ROM[7885] <= 32'b00000000010000100000000100010011;
ROM[7886] <= 32'b00000001010000000000001110010011;
ROM[7887] <= 32'b01000000011100011000001110110011;
ROM[7888] <= 32'b00000000010000111010000110000011;
ROM[7889] <= 32'b00000000100000111010001000000011;
ROM[7890] <= 32'b00000000110000111010001010000011;
ROM[7891] <= 32'b00000001000000111010001100000011;
ROM[7892] <= 32'b00000000000000001000000011100111;
ROM[7893] <= 32'b00000000000000001000001110110111;
ROM[7894] <= 32'b10111010000000111000001110010011;
ROM[7895] <= 32'b00000000111000111000001110110011;
ROM[7896] <= 32'b00000000011100010010000000100011;
ROM[7897] <= 32'b00000000010000010000000100010011;
ROM[7898] <= 32'b00000000001100010010000000100011;
ROM[7899] <= 32'b00000000010000010000000100010011;
ROM[7900] <= 32'b00000000010000010010000000100011;
ROM[7901] <= 32'b00000000010000010000000100010011;
ROM[7902] <= 32'b00000000010100010010000000100011;
ROM[7903] <= 32'b00000000010000010000000100010011;
ROM[7904] <= 32'b00000000011000010010000000100011;
ROM[7905] <= 32'b00000000010000010000000100010011;
ROM[7906] <= 32'b00000001010000000000001110010011;
ROM[7907] <= 32'b00000000000000111000001110010011;
ROM[7908] <= 32'b01000000011100010000001110110011;
ROM[7909] <= 32'b00000000011100000000001000110011;
ROM[7910] <= 32'b00000000001000000000000110110011;
ROM[7911] <= 32'b11111000100111111010000011101111;
ROM[7912] <= 32'b11111111110000010000000100010011;
ROM[7913] <= 32'b00000000000000010010001110000011;
ROM[7914] <= 32'b00000000011101100010000000100011;
ROM[7915] <= 32'b00000000000000001000001110110111;
ROM[7916] <= 32'b10111111100000111000001110010011;
ROM[7917] <= 32'b00000000111000111000001110110011;
ROM[7918] <= 32'b00000000011100010010000000100011;
ROM[7919] <= 32'b00000000010000010000000100010011;
ROM[7920] <= 32'b00000000001100010010000000100011;
ROM[7921] <= 32'b00000000010000010000000100010011;
ROM[7922] <= 32'b00000000010000010010000000100011;
ROM[7923] <= 32'b00000000010000010000000100010011;
ROM[7924] <= 32'b00000000010100010010000000100011;
ROM[7925] <= 32'b00000000010000010000000100010011;
ROM[7926] <= 32'b00000000011000010010000000100011;
ROM[7927] <= 32'b00000000010000010000000100010011;
ROM[7928] <= 32'b00000001010000000000001110010011;
ROM[7929] <= 32'b00000000000000111000001110010011;
ROM[7930] <= 32'b01000000011100010000001110110011;
ROM[7931] <= 32'b00000000011100000000001000110011;
ROM[7932] <= 32'b00000000001000000000000110110011;
ROM[7933] <= 32'b10100001000111111000000011101111;
ROM[7934] <= 32'b11111111110000010000000100010011;
ROM[7935] <= 32'b00000000000000010010001110000011;
ROM[7936] <= 32'b00000000011101100010000000100011;
ROM[7937] <= 32'b00000000000000001000001110110111;
ROM[7938] <= 32'b11000101000000111000001110010011;
ROM[7939] <= 32'b00000000111000111000001110110011;
ROM[7940] <= 32'b00000000011100010010000000100011;
ROM[7941] <= 32'b00000000010000010000000100010011;
ROM[7942] <= 32'b00000000001100010010000000100011;
ROM[7943] <= 32'b00000000010000010000000100010011;
ROM[7944] <= 32'b00000000010000010010000000100011;
ROM[7945] <= 32'b00000000010000010000000100010011;
ROM[7946] <= 32'b00000000010100010010000000100011;
ROM[7947] <= 32'b00000000010000010000000100010011;
ROM[7948] <= 32'b00000000011000010010000000100011;
ROM[7949] <= 32'b00000000010000010000000100010011;
ROM[7950] <= 32'b00000001010000000000001110010011;
ROM[7951] <= 32'b00000000000000111000001110010011;
ROM[7952] <= 32'b01000000011100010000001110110011;
ROM[7953] <= 32'b00000000011100000000001000110011;
ROM[7954] <= 32'b00000000001000000000000110110011;
ROM[7955] <= 32'b10001000010111111000000011101111;
ROM[7956] <= 32'b00000001010000000000001110010011;
ROM[7957] <= 32'b01000000011100011000001110110011;
ROM[7958] <= 32'b00000000000000111010000010000011;
ROM[7959] <= 32'b11111111110000010000000100010011;
ROM[7960] <= 32'b00000000000000010010001110000011;
ROM[7961] <= 32'b00000000011100100010000000100011;
ROM[7962] <= 32'b00000000010000100000000100010011;
ROM[7963] <= 32'b00000001010000000000001110010011;
ROM[7964] <= 32'b01000000011100011000001110110011;
ROM[7965] <= 32'b00000000010000111010000110000011;
ROM[7966] <= 32'b00000000100000111010001000000011;
ROM[7967] <= 32'b00000000110000111010001010000011;
ROM[7968] <= 32'b00000001000000111010001100000011;
ROM[7969] <= 32'b00000000000000001000000011100111;
ROM[7970] <= 32'b00000000000000000000001110010011;
ROM[7971] <= 32'b00000000011100010010000000100011;
ROM[7972] <= 32'b00000000010000010000000100010011;
ROM[7973] <= 32'b11111111110000010000000100010011;
ROM[7974] <= 32'b00000000000000010010001110000011;
ROM[7975] <= 32'b01000000011100000000001110110011;
ROM[7976] <= 32'b00000000000100111000001110010011;
ROM[7977] <= 32'b00000000011100010010000000100011;
ROM[7978] <= 32'b00000000010000010000000100010011;
ROM[7979] <= 32'b11111111110000010000000100010011;
ROM[7980] <= 32'b00000000000000010010001110000011;
ROM[7981] <= 32'b01000000011100000000001110110011;
ROM[7982] <= 32'b00000000000100111000001110010011;
ROM[7983] <= 32'b00000000011100010010000000100011;
ROM[7984] <= 32'b00000000010000010000000100010011;
ROM[7985] <= 32'b11111111110000010000000100010011;
ROM[7986] <= 32'b00000000000000010010001110000011;
ROM[7987] <= 32'b00000000000000111000101001100011;
ROM[7988] <= 32'b00000000000000001000001110110111;
ROM[7989] <= 32'b11001110010000111000001110010011;
ROM[7990] <= 32'b00000000111000111000001110110011;
ROM[7991] <= 32'b00000000000000111000000011100111;
ROM[7992] <= 32'b11111010100111111111000011101111;
ROM[7993] <= 32'b00000000000000000000001110010011;
ROM[7994] <= 32'b00000000011100010010000000100011;
ROM[7995] <= 32'b00000000010000010000000100010011;
ROM[7996] <= 32'b00000001010000000000001110010011;
ROM[7997] <= 32'b01000000011100011000001110110011;
ROM[7998] <= 32'b00000000000000111010000010000011;
ROM[7999] <= 32'b11111111110000010000000100010011;
ROM[8000] <= 32'b00000000000000010010001110000011;
ROM[8001] <= 32'b00000000011100100010000000100011;
ROM[8002] <= 32'b00000000010000100000000100010011;
ROM[8003] <= 32'b00000001010000000000001110010011;
ROM[8004] <= 32'b01000000011100011000001110110011;
ROM[8005] <= 32'b00000000010000111010000110000011;
ROM[8006] <= 32'b00000000100000111010001000000011;
ROM[8007] <= 32'b00000000110000111010001010000011;
ROM[8008] <= 32'b00000001000000111010001100000011;
ROM[8009] <= 32'b00000000000000001000000011100111;
ROM[8010] <= 32'b00000000000000010010000000100011;
ROM[8011] <= 32'b00000000010000010000000100010011;
ROM[8012] <= 32'b00000000000000010010000000100011;
ROM[8013] <= 32'b00000000010000010000000100010011;
ROM[8014] <= 32'b00000000000000000000001110010011;
ROM[8015] <= 32'b00000000011100010010000000100011;
ROM[8016] <= 32'b00000000010000010000000100010011;
ROM[8017] <= 32'b11111111110000010000000100010011;
ROM[8018] <= 32'b00000000000000010010001110000011;
ROM[8019] <= 32'b00000000011100011010000000100011;
ROM[8020] <= 32'b00000000000000011010001110000011;
ROM[8021] <= 32'b00000000011100010010000000100011;
ROM[8022] <= 32'b00000000010000010000000100010011;
ROM[8023] <= 32'b00000000000000100010001110000011;
ROM[8024] <= 32'b00000000011100010010000000100011;
ROM[8025] <= 32'b00000000010000010000000100010011;
ROM[8026] <= 32'b11111111110000010000000100010011;
ROM[8027] <= 32'b00000000000000010010001110000011;
ROM[8028] <= 32'b11111111110000010000000100010011;
ROM[8029] <= 32'b00000000000000010010010000000011;
ROM[8030] <= 32'b00000000011101000010001110110011;
ROM[8031] <= 32'b00000000011100010010000000100011;
ROM[8032] <= 32'b00000000010000010000000100010011;
ROM[8033] <= 32'b11111111110000010000000100010011;
ROM[8034] <= 32'b00000000000000010010001110000011;
ROM[8035] <= 32'b01000000011100000000001110110011;
ROM[8036] <= 32'b00000000000100111000001110010011;
ROM[8037] <= 32'b00000000011100010010000000100011;
ROM[8038] <= 32'b00000000010000010000000100010011;
ROM[8039] <= 32'b11111111110000010000000100010011;
ROM[8040] <= 32'b00000000000000010010001110000011;
ROM[8041] <= 32'b00000000000000111000101001100011;
ROM[8042] <= 32'b00000000000000001000001110110111;
ROM[8043] <= 32'b11101100000000111000001110010011;
ROM[8044] <= 32'b00000000111000111000001110110011;
ROM[8045] <= 32'b00000000000000111000000011100111;
ROM[8046] <= 32'b00000000000000000000001110010011;
ROM[8047] <= 32'b00000000011100010010000000100011;
ROM[8048] <= 32'b00000000010000010000000100010011;
ROM[8049] <= 32'b11111111110000010000000100010011;
ROM[8050] <= 32'b00000000000000010010001110000011;
ROM[8051] <= 32'b00000000011100011010001000100011;
ROM[8052] <= 32'b00000000010000011010001110000011;
ROM[8053] <= 32'b00000000011100010010000000100011;
ROM[8054] <= 32'b00000000010000010000000100010011;
ROM[8055] <= 32'b00000110010000000000001110010011;
ROM[8056] <= 32'b00000000011100010010000000100011;
ROM[8057] <= 32'b00000000010000010000000100010011;
ROM[8058] <= 32'b11111111110000010000000100010011;
ROM[8059] <= 32'b00000000000000010010001110000011;
ROM[8060] <= 32'b11111111110000010000000100010011;
ROM[8061] <= 32'b00000000000000010010010000000011;
ROM[8062] <= 32'b00000000011101000010001110110011;
ROM[8063] <= 32'b00000000011100010010000000100011;
ROM[8064] <= 32'b00000000010000010000000100010011;
ROM[8065] <= 32'b11111111110000010000000100010011;
ROM[8066] <= 32'b00000000000000010010001110000011;
ROM[8067] <= 32'b01000000011100000000001110110011;
ROM[8068] <= 32'b00000000000100111000001110010011;
ROM[8069] <= 32'b00000000011100010010000000100011;
ROM[8070] <= 32'b00000000010000010000000100010011;
ROM[8071] <= 32'b11111111110000010000000100010011;
ROM[8072] <= 32'b00000000000000010010001110000011;
ROM[8073] <= 32'b00000000000000111000101001100011;
ROM[8074] <= 32'b00000000000000001000001110110111;
ROM[8075] <= 32'b11100111110000111000001110010011;
ROM[8076] <= 32'b00000000111000111000001110110011;
ROM[8077] <= 32'b00000000000000111000000011100111;
ROM[8078] <= 32'b00000000010000011010001110000011;
ROM[8079] <= 32'b00000000011100010010000000100011;
ROM[8080] <= 32'b00000000010000010000000100010011;
ROM[8081] <= 32'b00000000000100000000001110010011;
ROM[8082] <= 32'b00000000011100010010000000100011;
ROM[8083] <= 32'b00000000010000010000000100010011;
ROM[8084] <= 32'b11111111110000010000000100010011;
ROM[8085] <= 32'b00000000000000010010001110000011;
ROM[8086] <= 32'b11111111110000010000000100010011;
ROM[8087] <= 32'b00000000000000010010010000000011;
ROM[8088] <= 32'b00000000011101000000001110110011;
ROM[8089] <= 32'b00000000011100010010000000100011;
ROM[8090] <= 32'b00000000010000010000000100010011;
ROM[8091] <= 32'b11111111110000010000000100010011;
ROM[8092] <= 32'b00000000000000010010001110000011;
ROM[8093] <= 32'b00000000011100011010001000100011;
ROM[8094] <= 32'b11110101100111111111000011101111;
ROM[8095] <= 32'b00000000000000011010001110000011;
ROM[8096] <= 32'b00000000011100010010000000100011;
ROM[8097] <= 32'b00000000010000010000000100010011;
ROM[8098] <= 32'b00000000000100000000001110010011;
ROM[8099] <= 32'b00000000011100010010000000100011;
ROM[8100] <= 32'b00000000010000010000000100010011;
ROM[8101] <= 32'b11111111110000010000000100010011;
ROM[8102] <= 32'b00000000000000010010001110000011;
ROM[8103] <= 32'b11111111110000010000000100010011;
ROM[8104] <= 32'b00000000000000010010010000000011;
ROM[8105] <= 32'b00000000011101000000001110110011;
ROM[8106] <= 32'b00000000011100010010000000100011;
ROM[8107] <= 32'b00000000010000010000000100010011;
ROM[8108] <= 32'b11111111110000010000000100010011;
ROM[8109] <= 32'b00000000000000010010001110000011;
ROM[8110] <= 32'b00000000011100011010000000100011;
ROM[8111] <= 32'b11101001010111111111000011101111;
ROM[8112] <= 32'b00000000000000000000001110010011;
ROM[8113] <= 32'b00000000011100010010000000100011;
ROM[8114] <= 32'b00000000010000010000000100010011;
ROM[8115] <= 32'b00000001010000000000001110010011;
ROM[8116] <= 32'b01000000011100011000001110110011;
ROM[8117] <= 32'b00000000000000111010000010000011;
ROM[8118] <= 32'b11111111110000010000000100010011;
ROM[8119] <= 32'b00000000000000010010001110000011;
ROM[8120] <= 32'b00000000011100100010000000100011;
ROM[8121] <= 32'b00000000010000100000000100010011;
ROM[8122] <= 32'b00000001010000000000001110010011;
ROM[8123] <= 32'b01000000011100011000001110110011;
ROM[8124] <= 32'b00000000010000111010000110000011;
ROM[8125] <= 32'b00000000100000111010001000000011;
ROM[8126] <= 32'b00000000110000111010001010000011;
ROM[8127] <= 32'b00000001000000111010001100000011;
ROM[8128] <= 32'b00000000000000001000000011100111;
ROM[8129] <= 32'b00000000000000111000000010010011;
        end
    assign address = addr[16:2];
    assign Inst = ROM[address];
        
endmodule