module ROM (                    //Instruction Memory
    input [16:0] addr,
    input clock,
    output [31:0] Inst
    );
    wire [14:0] address;
    
    (* ram_style="block" *)
    reg [31:0] ROM[32767:0];

    initial
        begin
ROM[0] <= 32'b00000000000000000010011100110111;
ROM[1] <= 32'b01011000000001110000011100010011;
ROM[2] <= 32'b00000000000000100010011010110111;
ROM[3] <= 32'b01011000000001101000011010010011;
ROM[4] <= 32'b00010000000001101000000100010011;
ROM[5] <= 32'b00000000000000010000000110010011;
ROM[6] <= 32'b00000000000001101000011000010011;
ROM[7] <= 32'b00000000000000010010000000100011;
ROM[8] <= 32'b00000000010000010000000100010011;
ROM[9] <= 32'b00000000101000000000001110010011;
ROM[10] <= 32'b00000000011100010010000000100011;
ROM[11] <= 32'b00000000010000010000000100010011;
ROM[12] <= 32'b00000000000000000000001110110111;
ROM[13] <= 32'b00000111110000111000001110010011;
ROM[14] <= 32'b00000000111000111000001110110011;
ROM[15] <= 32'b00000000011100010010000000100011;
ROM[16] <= 32'b00000000010000010000000100010011;
ROM[17] <= 32'b00000000001100010010000000100011;
ROM[18] <= 32'b00000000010000010000000100010011;
ROM[19] <= 32'b00000000010000010010000000100011;
ROM[20] <= 32'b00000000010000010000000100010011;
ROM[21] <= 32'b00000000010100010010000000100011;
ROM[22] <= 32'b00000000010000010000000100010011;
ROM[23] <= 32'b00000000011000010010000000100011;
ROM[24] <= 32'b00000000010000010000000100010011;
ROM[25] <= 32'b00000001010000000000001110010011;
ROM[26] <= 32'b00000000010000111000001110010011;
ROM[27] <= 32'b01000000011100010000001110110011;
ROM[28] <= 32'b00000000011100000000001000110011;
ROM[29] <= 32'b00000000001000000000000110110011;
ROM[30] <= 32'b00000001010000000000000011101111;
ROM[31] <= 32'b11111111110000010000000100010011;
ROM[32] <= 32'b00000000000000010010001110000011;
ROM[33] <= 32'b00000000011100011010000000100011;
ROM[34] <= 32'b00100110010000000000000011101111;
ROM[35] <= 32'b00000000000000010010000000100011;
ROM[36] <= 32'b00000000010000010000000100010011;
ROM[37] <= 32'b00000000000000010010000000100011;
ROM[38] <= 32'b00000000010000010000000100010011;
ROM[39] <= 32'b00000000000000010010000000100011;
ROM[40] <= 32'b00000000010000010000000100010011;
ROM[41] <= 32'b00000000000000010010000000100011;
ROM[42] <= 32'b00000000010000010000000100010011;
ROM[43] <= 32'b00000000001000000000001110010011;
ROM[44] <= 32'b00000000011100010010000000100011;
ROM[45] <= 32'b00000000010000010000000100010011;
ROM[46] <= 32'b11111111110000010000000100010011;
ROM[47] <= 32'b00000000000000010010001110000011;
ROM[48] <= 32'b00000000011100011010011000100011;
ROM[49] <= 32'b00000000000000000000001110010011;
ROM[50] <= 32'b00000000011100010010000000100011;
ROM[51] <= 32'b00000000010000010000000100010011;
ROM[52] <= 32'b11111111110000010000000100010011;
ROM[53] <= 32'b00000000000000010010001110000011;
ROM[54] <= 32'b00000000011100011010000000100011;
ROM[55] <= 32'b00000000000100000000001110010011;
ROM[56] <= 32'b00000000011100010010000000100011;
ROM[57] <= 32'b00000000010000010000000100010011;
ROM[58] <= 32'b11111111110000010000000100010011;
ROM[59] <= 32'b00000000000000010010001110000011;
ROM[60] <= 32'b00000000011100011010001000100011;
ROM[61] <= 32'b00000000000000100010001110000011;
ROM[62] <= 32'b00000000011100010010000000100011;
ROM[63] <= 32'b00000000010000010000000100010011;
ROM[64] <= 32'b00000000000100000000001110010011;
ROM[65] <= 32'b00000000011100010010000000100011;
ROM[66] <= 32'b00000000010000010000000100010011;
ROM[67] <= 32'b11111111110000010000000100010011;
ROM[68] <= 32'b00000000000000010010001110000011;
ROM[69] <= 32'b11111111110000010000000100010011;
ROM[70] <= 32'b00000000000000010010010000000011;
ROM[71] <= 32'b00000000011101000010010010110011;
ROM[72] <= 32'b00000000100000111010010100110011;
ROM[73] <= 32'b00000000101001001000001110110011;
ROM[74] <= 32'b00000000000100111000001110010011;
ROM[75] <= 32'b00000000000100111111001110010011;
ROM[76] <= 32'b00000000011100010010000000100011;
ROM[77] <= 32'b00000000010000010000000100010011;
ROM[78] <= 32'b11111111110000010000000100010011;
ROM[79] <= 32'b00000000000000010010001110000011;
ROM[80] <= 32'b00000000000000111000101001100011;
ROM[81] <= 32'b00000000000000000000001110110111;
ROM[82] <= 32'b00010101100000111000001110010011;
ROM[83] <= 32'b00000000111000111000001110110011;
ROM[84] <= 32'b00000000000000111000000011100111;
ROM[85] <= 32'b00000100000000000000000011101111;
ROM[86] <= 32'b00000000000000000000001110010011;
ROM[87] <= 32'b00000000011100010010000000100011;
ROM[88] <= 32'b00000000010000010000000100010011;
ROM[89] <= 32'b11111111110000010000000100010011;
ROM[90] <= 32'b00000000000000010010001110000011;
ROM[91] <= 32'b00000000011100100010000000100011;
ROM[92] <= 32'b00000000010000100000000100010011;
ROM[93] <= 32'b00000001010000000000001110010011;
ROM[94] <= 32'b01000000011100011000001110110011;
ROM[95] <= 32'b00000000000000111010000010000011;
ROM[96] <= 32'b00000000010000111010000110000011;
ROM[97] <= 32'b00000000100000111010001000000011;
ROM[98] <= 32'b00000000110000111010001010000011;
ROM[99] <= 32'b00000001000000111010001100000011;
ROM[100] <= 32'b00000000000000001000000011100111;
ROM[101] <= 32'b00000000110000011010001110000011;
ROM[102] <= 32'b00000000011100010010000000100011;
ROM[103] <= 32'b00000000010000010000000100010011;
ROM[104] <= 32'b00000000000000100010001110000011;
ROM[105] <= 32'b00000000011100010010000000100011;
ROM[106] <= 32'b00000000010000010000000100010011;
ROM[107] <= 32'b11111111110000010000000100010011;
ROM[108] <= 32'b00000000000000010010001110000011;
ROM[109] <= 32'b11111111110000010000000100010011;
ROM[110] <= 32'b00000000000000010010010000000011;
ROM[111] <= 32'b00000000011101000010001110110011;
ROM[112] <= 32'b00000000011100010010000000100011;
ROM[113] <= 32'b00000000010000010000000100010011;
ROM[114] <= 32'b11111111110000010000000100010011;
ROM[115] <= 32'b00000000000000010010001110000011;
ROM[116] <= 32'b01000000011100000000001110110011;
ROM[117] <= 32'b00000000000100111000001110010011;
ROM[118] <= 32'b00000000011100010010000000100011;
ROM[119] <= 32'b00000000010000010000000100010011;
ROM[120] <= 32'b11111111110000010000000100010011;
ROM[121] <= 32'b00000000000000010010001110000011;
ROM[122] <= 32'b00000000000000111000101001100011;
ROM[123] <= 32'b00000000000000000000001110110111;
ROM[124] <= 32'b00101011000000111000001110010011;
ROM[125] <= 32'b00000000111000111000001110110011;
ROM[126] <= 32'b00000000000000111000000011100111;
ROM[127] <= 32'b00000000000000011010001110000011;
ROM[128] <= 32'b00000000011100010010000000100011;
ROM[129] <= 32'b00000000010000010000000100010011;
ROM[130] <= 32'b00000000010000011010001110000011;
ROM[131] <= 32'b00000000011100010010000000100011;
ROM[132] <= 32'b00000000010000010000000100010011;
ROM[133] <= 32'b11111111110000010000000100010011;
ROM[134] <= 32'b00000000000000010010001110000011;
ROM[135] <= 32'b11111111110000010000000100010011;
ROM[136] <= 32'b00000000000000010010010000000011;
ROM[137] <= 32'b00000000100000111000001110110011;
ROM[138] <= 32'b00000000011100010010000000100011;
ROM[139] <= 32'b00000000010000010000000100010011;
ROM[140] <= 32'b11111111110000010000000100010011;
ROM[141] <= 32'b00000000000000010010001110000011;
ROM[142] <= 32'b00000000011100011010010000100011;
ROM[143] <= 32'b00000000010000011010001110000011;
ROM[144] <= 32'b00000000011100010010000000100011;
ROM[145] <= 32'b00000000010000010000000100010011;
ROM[146] <= 32'b11111111110000010000000100010011;
ROM[147] <= 32'b00000000000000010010001110000011;
ROM[148] <= 32'b00000000011100011010000000100011;
ROM[149] <= 32'b00000000100000011010001110000011;
ROM[150] <= 32'b00000000011100010010000000100011;
ROM[151] <= 32'b00000000010000010000000100010011;
ROM[152] <= 32'b11111111110000010000000100010011;
ROM[153] <= 32'b00000000000000010010001110000011;
ROM[154] <= 32'b00000000011100011010001000100011;
ROM[155] <= 32'b00000000110000011010001110000011;
ROM[156] <= 32'b00000000011100010010000000100011;
ROM[157] <= 32'b00000000010000010000000100010011;
ROM[158] <= 32'b00000000000100000000001110010011;
ROM[159] <= 32'b00000000011100010010000000100011;
ROM[160] <= 32'b00000000010000010000000100010011;
ROM[161] <= 32'b11111111110000010000000100010011;
ROM[162] <= 32'b00000000000000010010001110000011;
ROM[163] <= 32'b11111111110000010000000100010011;
ROM[164] <= 32'b00000000000000010010010000000011;
ROM[165] <= 32'b00000000100000111000001110110011;
ROM[166] <= 32'b00000000011100010010000000100011;
ROM[167] <= 32'b00000000010000010000000100010011;
ROM[168] <= 32'b11111111110000010000000100010011;
ROM[169] <= 32'b00000000000000010010001110000011;
ROM[170] <= 32'b00000000011100011010011000100011;
ROM[171] <= 32'b11101110100111111111000011101111;
ROM[172] <= 32'b00000000010000011010001110000011;
ROM[173] <= 32'b00000000011100010010000000100011;
ROM[174] <= 32'b00000000010000010000000100010011;
ROM[175] <= 32'b11111111110000010000000100010011;
ROM[176] <= 32'b00000000000000010010001110000011;
ROM[177] <= 32'b00000000011100100010000000100011;
ROM[178] <= 32'b00000000010000100000000100010011;
ROM[179] <= 32'b00000001010000000000001110010011;
ROM[180] <= 32'b01000000011100011000001110110011;
ROM[181] <= 32'b00000000000000111010000010000011;
ROM[182] <= 32'b00000000010000111010000110000011;
ROM[183] <= 32'b00000000100000111010001000000011;
ROM[184] <= 32'b00000000110000111010001010000011;
ROM[185] <= 32'b00000001000000111010001100000011;
ROM[186] <= 32'b00000000000000001000000011100111;
ROM[187] <= 32'b00000000000000111000000010010011;

        end
    assign address = addr[16:2];
    assign Inst = ROM[address];
        
endmodule


						
						

// module ROM ( //Instruction Memory
//     input [15:0] address,
//     input clock,
//     input IRWrite,
//     output reg [31:0] IR
//     );
    
//     (* ram_style="block" *)
//     reg [31:0] ROM[16383:0];

//     initial
//         begin
//             $readmemb("os.mem", ROM, 0, 16383);
//             IR <= 32'd15;
//         end
    
//     always @(posedge clock)
//         begin
//             if( IRWrite )
//                 IR <= ROM[address];
//         end
        
// endmodule

						
						


						
						
