module ROM ( //Instruction Memory
    input [16:0] addr,
    input clock,
    output [31:0] Inst
    );
    wire [14:0] address;
    
    (* ram_style="block" *)
    reg [31:0] ROM[32767:0];

    initial
        begin
    ROM[0] <= 32'b00000000000000000010011100110111;
ROM[1] <= 32'b01011000000001110000011100010011;
ROM[2] <= 32'b00000000000000100010011010110111;
ROM[3] <= 32'b01011000000001101000011010010011;
ROM[4] <= 32'b00000100000001101010000000100011;
ROM[5] <= 32'b00000100000001101010001000100011;
ROM[6] <= 32'b00000100000001101010010000100011;
ROM[7] <= 32'b00000100000001101010011000100011;
ROM[8] <= 32'b00000100000001101010100000100011;
ROM[9] <= 32'b00000100000001101010101000100011;
ROM[10] <= 32'b00000100000001101010110000100011;
ROM[11] <= 32'b00000100000001101010111000100011;
ROM[12] <= 32'b00000110000001101010000000100011;
ROM[13] <= 32'b00000110000001101010001000100011;
ROM[14] <= 32'b00000110000001101010010000100011;
ROM[15] <= 32'b00000110000001101010011000100011;
ROM[16] <= 32'b00000110000001101010100000100011;
ROM[17] <= 32'b00000110000001101010101000100011;
ROM[18] <= 32'b00000110000001101010110000100011;
ROM[19] <= 32'b00000110000001101010111000100011;
ROM[20] <= 32'b00001000000001101010000000100011;
ROM[21] <= 32'b00001000000001101010001000100011;
ROM[22] <= 32'b00001000000001101010010000100011;
ROM[23] <= 32'b00001000000001101010011000100011;
ROM[24] <= 32'b00001000000001101010100000100011;
ROM[25] <= 32'b00001000000001101010101000100011;
ROM[26] <= 32'b00001000000001101010110000100011;
ROM[27] <= 32'b00001000000001101010111000100011;
ROM[28] <= 32'b00001010000001101010000000100011;
ROM[29] <= 32'b00001010000001101010001000100011;
ROM[30] <= 32'b00001010000001101010010000100011;
ROM[31] <= 32'b00001010000001101010011000100011;
ROM[32] <= 32'b00001010000001101010100000100011;
ROM[33] <= 32'b00001010000001101010101000100011;
ROM[34] <= 32'b00001010000001101010110000100011;
ROM[35] <= 32'b00001010000001101010111000100011;
ROM[36] <= 32'b00001100000001101010000000100011;
ROM[37] <= 32'b00001100000001101010001000100011;
ROM[38] <= 32'b00001100000001101010010000100011;
ROM[39] <= 32'b00001100000001101010011000100011;
ROM[40] <= 32'b00001100000001101010100000100011;
ROM[41] <= 32'b00001100000001101010101000100011;
ROM[42] <= 32'b00001100000001101010110000100011;
ROM[43] <= 32'b00001100000001101010111000100011;
ROM[44] <= 32'b00001110000001101010000000100011;
ROM[45] <= 32'b00001110000001101010001000100011;
ROM[46] <= 32'b00001110000001101010010000100011;
ROM[47] <= 32'b00001110000001101010011000100011;
ROM[48] <= 32'b00001110000001101010100000100011;
ROM[49] <= 32'b00001110000001101010101000100011;
ROM[50] <= 32'b00001110000001101010110000100011;
ROM[51] <= 32'b00001110000001101010111000100011;
ROM[52] <= 32'b00010000000001101010000000100011;
ROM[53] <= 32'b00010000000001101010001000100011;
ROM[54] <= 32'b00010000000001101010010000100011;
ROM[55] <= 32'b00010000000001101010011000100011;
ROM[56] <= 32'b00010000000001101010100000100011;
ROM[57] <= 32'b00010000000001101010101000100011;
ROM[58] <= 32'b00010000000001101010110000100011;
ROM[59] <= 32'b00010000000001101010111000100011;
ROM[60] <= 32'b00010010000001101010000000100011;
ROM[61] <= 32'b00010010000001101010001000100011;
ROM[62] <= 32'b00010010000001101010010000100011;
ROM[63] <= 32'b00010010000001101010011000100011;
ROM[64] <= 32'b00010010000001101010100000100011;
ROM[65] <= 32'b00010010000001101010101000100011;
ROM[66] <= 32'b00010010000001101010110000100011;
ROM[67] <= 32'b00010010000001101010111000100011;
ROM[68] <= 32'b00010100000001101010000000100011;
ROM[69] <= 32'b00010100000001101010001000100011;
ROM[70] <= 32'b00010100000001101010010000100011;
ROM[71] <= 32'b00010100000001101010011000100011;
ROM[72] <= 32'b00010100000001101010100000100011;
ROM[73] <= 32'b00010100000001101010101000100011;
ROM[74] <= 32'b00010100000001101010110000100011;
ROM[75] <= 32'b00010100000001101010111000100011;
ROM[76] <= 32'b00010110000001101010000000100011;
ROM[77] <= 32'b00010110000001101010001000100011;
ROM[78] <= 32'b00010110000001101010010000100011;
ROM[79] <= 32'b00010110000001101010011000100011;
ROM[80] <= 32'b00010110000001101010100000100011;
ROM[81] <= 32'b00010110000001101010101000100011;
ROM[82] <= 32'b00010110000001101010110000100011;
ROM[83] <= 32'b00010110000001101010111000100011;
ROM[84] <= 32'b00011000000001101010000000100011;
ROM[85] <= 32'b00011000000001101010001000100011;
ROM[86] <= 32'b00011000000001101010010000100011;
ROM[87] <= 32'b00011000000001101010011000100011;
ROM[88] <= 32'b00011000000001101010100000100011;
ROM[89] <= 32'b00011000000001101010101000100011;
ROM[90] <= 32'b00011000000001101010110000100011;
ROM[91] <= 32'b00011000000001101010111000100011;
ROM[92] <= 32'b00011010000001101010000000100011;
ROM[93] <= 32'b00011010000001101010001000100011;
ROM[94] <= 32'b00011010000001101010010000100011;
ROM[95] <= 32'b00011010000001101010011000100011;
ROM[96] <= 32'b00011010000001101010100000100011;
ROM[97] <= 32'b00011010000001101010101000100011;
ROM[98] <= 32'b00011010000001101010110000100011;
ROM[99] <= 32'b00011010000001101010111000100011;
ROM[100] <= 32'b00011100000001101010000000100011;
ROM[101] <= 32'b00011100000001101010001000100011;
ROM[102] <= 32'b00011100000001101010010000100011;
ROM[103] <= 32'b00011100000001101010011000100011;
ROM[104] <= 32'b00011100000001101010100000100011;
ROM[105] <= 32'b00011100000001101010101000100011;
ROM[106] <= 32'b00011100000001101010110000100011;
ROM[107] <= 32'b00011100000001101010111000100011;
ROM[108] <= 32'b00011110000001101010000000100011;
ROM[109] <= 32'b00011110000001101010001000100011;
ROM[110] <= 32'b00011110000001101010010000100011;
ROM[111] <= 32'b00011110000001101010011000100011;
ROM[112] <= 32'b00011110000001101010100000100011;
ROM[113] <= 32'b00011110000001101010101000100011;
ROM[114] <= 32'b00011110000001101010110000100011;
ROM[115] <= 32'b00011110000001101010111000100011;
ROM[116] <= 32'b00100000000001101010000000100011;
ROM[117] <= 32'b00100000000001101010001000100011;
ROM[118] <= 32'b00100000000001101010010000100011;
ROM[119] <= 32'b00100000000001101010011000100011;
ROM[120] <= 32'b00100000000001101010100000100011;
ROM[121] <= 32'b00100000000001101010101000100011;
ROM[122] <= 32'b00100000000001101010110000100011;
ROM[123] <= 32'b00100000000001101010111000100011;
ROM[124] <= 32'b00100010000001101010000000100011;
ROM[125] <= 32'b00100010000001101010001000100011;
ROM[126] <= 32'b00100010000001101010010000100011;
ROM[127] <= 32'b00100010000001101010011000100011;
ROM[128] <= 32'b00100010000001101010100000100011;
ROM[129] <= 32'b00100010000001101010101000100011;
ROM[130] <= 32'b00100010000001101010110000100011;
ROM[131] <= 32'b00100010000001101010111000100011;
ROM[132] <= 32'b00100100000001101010000000100011;
ROM[133] <= 32'b00100100000001101010001000100011;
ROM[134] <= 32'b00100100000001101010010000100011;
ROM[135] <= 32'b00100100000001101010011000100011;
ROM[136] <= 32'b00100100000001101010100000100011;
ROM[137] <= 32'b00100100000001101010101000100011;
ROM[138] <= 32'b00100100000001101010110000100011;
ROM[139] <= 32'b00100100000001101010111000100011;
ROM[140] <= 32'b00100110000001101010000000100011;
ROM[141] <= 32'b00100110000001101010001000100011;
ROM[142] <= 32'b00100110000001101010010000100011;
ROM[143] <= 32'b00100110000001101010011000100011;
ROM[144] <= 32'b00100110000001101010100000100011;
ROM[145] <= 32'b00100110000001101010101000100011;
ROM[146] <= 32'b00100110000001101010110000100011;
ROM[147] <= 32'b00100110000001101010111000100011;
ROM[148] <= 32'b00101000000001101010000000100011;
ROM[149] <= 32'b00101000000001101010001000100011;
ROM[150] <= 32'b00101000000001101010010000100011;
ROM[151] <= 32'b00101000000001101010011000100011;
ROM[152] <= 32'b00101000000001101010100000100011;
ROM[153] <= 32'b00101000000001101010101000100011;
ROM[154] <= 32'b00101000000001101010110000100011;
ROM[155] <= 32'b00101000000001101010111000100011;
ROM[156] <= 32'b00101010000001101010000000100011;
ROM[157] <= 32'b00101010000001101010001000100011;
ROM[158] <= 32'b00101010000001101010010000100011;
ROM[159] <= 32'b00101010000001101010011000100011;
ROM[160] <= 32'b00101010000001101010100000100011;
ROM[161] <= 32'b00101010000001101010101000100011;
ROM[162] <= 32'b00101010000001101010110000100011;
ROM[163] <= 32'b00101010000001101010111000100011;
ROM[164] <= 32'b00101100000001101010000000100011;
ROM[165] <= 32'b00101100000001101010001000100011;
ROM[166] <= 32'b00101100000001101010010000100011;
ROM[167] <= 32'b00101100000001101010011000100011;
ROM[168] <= 32'b00101100000001101010100000100011;
ROM[169] <= 32'b00101100000001101010101000100011;
ROM[170] <= 32'b00101100000001101010110000100011;
ROM[171] <= 32'b00101100000001101010111000100011;
ROM[172] <= 32'b00101110000001101010000000100011;
ROM[173] <= 32'b00101110000001101010001000100011;
ROM[174] <= 32'b00101110000001101010010000100011;
ROM[175] <= 32'b00101110000001101010011000100011;
ROM[176] <= 32'b00101110000001101010100000100011;
ROM[177] <= 32'b00101110000001101010101000100011;
ROM[178] <= 32'b00101110000001101010110000100011;
ROM[179] <= 32'b00101110000001101010111000100011;
ROM[180] <= 32'b00110000000001101010000000100011;
ROM[181] <= 32'b00110000000001101010001000100011;
ROM[182] <= 32'b00110000000001101010010000100011;
ROM[183] <= 32'b00110000000001101010011000100011;
ROM[184] <= 32'b00110000000001101010100000100011;
ROM[185] <= 32'b00110000000001101010101000100011;
ROM[186] <= 32'b00110000000001101010110000100011;
ROM[187] <= 32'b00110000000001101010111000100011;
ROM[188] <= 32'b00110010000001101010000000100011;
ROM[189] <= 32'b00110010000001101010001000100011;
ROM[190] <= 32'b00110010000001101010010000100011;
ROM[191] <= 32'b00110010000001101010011000100011;
ROM[192] <= 32'b00110010000001101010100000100011;
ROM[193] <= 32'b00110010000001101010101000100011;
ROM[194] <= 32'b00110010000001101010110000100011;
ROM[195] <= 32'b00110010000001101010111000100011;
ROM[196] <= 32'b00110100000001101010000000100011;
ROM[197] <= 32'b00110100000001101010001000100011;
ROM[198] <= 32'b00110100000001101010010000100011;
ROM[199] <= 32'b00110100000001101010011000100011;
ROM[200] <= 32'b00110100000001101010100000100011;
ROM[201] <= 32'b00110100000001101010101000100011;
ROM[202] <= 32'b00110100000001101010110000100011;
ROM[203] <= 32'b00110100000001101010111000100011;
ROM[204] <= 32'b00110110000001101010000000100011;
ROM[205] <= 32'b00110110000001101010001000100011;
ROM[206] <= 32'b00110110000001101010010000100011;
ROM[207] <= 32'b00110110000001101010011000100011;
ROM[208] <= 32'b00110110000001101010100000100011;
ROM[209] <= 32'b00110110000001101010101000100011;
ROM[210] <= 32'b00110110000001101010110000100011;
ROM[211] <= 32'b00110110000001101010111000100011;
ROM[212] <= 32'b00111000000001101010000000100011;
ROM[213] <= 32'b00111000000001101010001000100011;
ROM[214] <= 32'b00111000000001101010010000100011;
ROM[215] <= 32'b00111000000001101010011000100011;
ROM[216] <= 32'b00111000000001101010100000100011;
ROM[217] <= 32'b00111000000001101010101000100011;
ROM[218] <= 32'b00111000000001101010110000100011;
ROM[219] <= 32'b00111000000001101010111000100011;
ROM[220] <= 32'b00111010000001101010000000100011;
ROM[221] <= 32'b00111010000001101010001000100011;
ROM[222] <= 32'b00111010000001101010010000100011;
ROM[223] <= 32'b00111010000001101010011000100011;
ROM[224] <= 32'b00111010000001101010100000100011;
ROM[225] <= 32'b00111010000001101010101000100011;
ROM[226] <= 32'b00111010000001101010110000100011;
ROM[227] <= 32'b00111010000001101010111000100011;
ROM[228] <= 32'b00111100000001101010000000100011;
ROM[229] <= 32'b00111100000001101010001000100011;
ROM[230] <= 32'b00111100000001101010010000100011;
ROM[231] <= 32'b00111100000001101010011000100011;
ROM[232] <= 32'b00111100000001101010100000100011;
ROM[233] <= 32'b00111100000001101010101000100011;
ROM[234] <= 32'b00111100000001101010110000100011;
ROM[235] <= 32'b00111100000001101010111000100011;
ROM[236] <= 32'b00111110000001101010000000100011;
ROM[237] <= 32'b00111110000001101010001000100011;
ROM[238] <= 32'b00111110000001101010010000100011;
ROM[239] <= 32'b00111110000001101010011000100011;
ROM[240] <= 32'b00111110000001101010100000100011;
ROM[241] <= 32'b00111110000001101010101000100011;
ROM[242] <= 32'b00111110000001101010110000100011;
ROM[243] <= 32'b00111110000001101010111000100011;
ROM[244] <= 32'b00000000000001101000011000010011;
ROM[245] <= 32'b01000000000001101000000100010011;
ROM[246] <= 32'b00000000000000010000000110010011;
ROM[247] <= 32'b00000000000000010000001000010011;
ROM[248] <= 32'b00000000000000010000001010010011;
ROM[249] <= 32'b00000000000000010000001100010011;
ROM[250] <= 32'b00000000000000000000001110110111;
ROM[251] <= 32'b01000011010000111000001110010011;
ROM[252] <= 32'b00000000111000111000001110110011;
ROM[253] <= 32'b00000000011100010010000000100011;
ROM[254] <= 32'b00000000010000010000000100010011;
ROM[255] <= 32'b00000000001100010010000000100011;
ROM[256] <= 32'b00000000010000010000000100010011;
ROM[257] <= 32'b00000000010000010010000000100011;
ROM[258] <= 32'b00000000010000010000000100010011;
ROM[259] <= 32'b00000000010100010010000000100011;
ROM[260] <= 32'b00000000010000010000000100010011;
ROM[261] <= 32'b00000000011000010010000000100011;
ROM[262] <= 32'b00000000010000010000000100010011;
ROM[263] <= 32'b00000001010000000000001110010011;
ROM[264] <= 32'b00000000000000111000001110010011;
ROM[265] <= 32'b01000000011100010000001110110011;
ROM[266] <= 32'b00000000011100000000001000110011;
ROM[267] <= 32'b00000000001000000000000110110011;
ROM[268] <= 32'b01110101100000010010000011101111;
ROM[269] <= 32'b11111111110000010000000100010011;
ROM[270] <= 32'b00000000000000010010001110000011;
ROM[271] <= 32'b00110010110100010010000011101111;
ROM[272] <= 32'b00000000000000100010001110000011;
ROM[273] <= 32'b00000000011100010010000000100011;
ROM[274] <= 32'b00000000010000010000000100010011;
ROM[275] <= 32'b00000000000000000000001110110111;
ROM[276] <= 32'b01001001100000111000001110010011;
ROM[277] <= 32'b00000000111000111000001110110011;
ROM[278] <= 32'b00000000011100010010000000100011;
ROM[279] <= 32'b00000000010000010000000100010011;
ROM[280] <= 32'b00000000001100010010000000100011;
ROM[281] <= 32'b00000000010000010000000100010011;
ROM[282] <= 32'b00000000010000010010000000100011;
ROM[283] <= 32'b00000000010000010000000100010011;
ROM[284] <= 32'b00000000010100010010000000100011;
ROM[285] <= 32'b00000000010000010000000100010011;
ROM[286] <= 32'b00000000011000010010000000100011;
ROM[287] <= 32'b00000000010000010000000100010011;
ROM[288] <= 32'b00000001010000000000001110010011;
ROM[289] <= 32'b00000000010000111000001110010011;
ROM[290] <= 32'b01000000011100010000001110110011;
ROM[291] <= 32'b00000000011100000000001000110011;
ROM[292] <= 32'b00000000001000000000000110110011;
ROM[293] <= 32'b01110111000100001001000011101111;
ROM[294] <= 32'b00000001010000000000001110010011;
ROM[295] <= 32'b01000000011100011000001110110011;
ROM[296] <= 32'b00000000000000111010000010000011;
ROM[297] <= 32'b11111111110000010000000100010011;
ROM[298] <= 32'b00000000000000010010001110000011;
ROM[299] <= 32'b00000000011100100010000000100011;
ROM[300] <= 32'b00000000010000100000000100010011;
ROM[301] <= 32'b00000001010000000000001110010011;
ROM[302] <= 32'b01000000011100011000001110110011;
ROM[303] <= 32'b00000000010000111010000110000011;
ROM[304] <= 32'b00000000100000111010001000000011;
ROM[305] <= 32'b00000000110000111010001010000011;
ROM[306] <= 32'b00000001000000111010001100000011;
ROM[307] <= 32'b00000000000000001000000011100111;
ROM[308] <= 32'b00000000000000100010001110000011;
ROM[309] <= 32'b00000000000000111000001010010011;
ROM[310] <= 32'b00000000010100010010000000100011;
ROM[311] <= 32'b00000000010000010000000100010011;
ROM[312] <= 32'b00000000000000000000001110110111;
ROM[313] <= 32'b01010010110000111000001110010011;
ROM[314] <= 32'b00000000111000111000001110110011;
ROM[315] <= 32'b00000000011100010010000000100011;
ROM[316] <= 32'b00000000010000010000000100010011;
ROM[317] <= 32'b00000000001100010010000000100011;
ROM[318] <= 32'b00000000010000010000000100010011;
ROM[319] <= 32'b00000000010000010010000000100011;
ROM[320] <= 32'b00000000010000010000000100010011;
ROM[321] <= 32'b00000000010100010010000000100011;
ROM[322] <= 32'b00000000010000010000000100010011;
ROM[323] <= 32'b00000000011000010010000000100011;
ROM[324] <= 32'b00000000010000010000000100010011;
ROM[325] <= 32'b00000001010000000000001110010011;
ROM[326] <= 32'b00000000010000111000001110010011;
ROM[327] <= 32'b01000000011100010000001110110011;
ROM[328] <= 32'b00000000011100000000001000110011;
ROM[329] <= 32'b00000000001000000000000110110011;
ROM[330] <= 32'b01110101010000001001000011101111;
ROM[331] <= 32'b11111111110000010000000100010011;
ROM[332] <= 32'b00000000000000010010001110000011;
ROM[333] <= 32'b00000000011101100010000000100011;
ROM[334] <= 32'b00000000000000000000001110010011;
ROM[335] <= 32'b00000000011100010010000000100011;
ROM[336] <= 32'b00000000010000010000000100010011;
ROM[337] <= 32'b00000001010000000000001110010011;
ROM[338] <= 32'b01000000011100011000001110110011;
ROM[339] <= 32'b00000000000000111010000010000011;
ROM[340] <= 32'b11111111110000010000000100010011;
ROM[341] <= 32'b00000000000000010010001110000011;
ROM[342] <= 32'b00000000011100100010000000100011;
ROM[343] <= 32'b00000000010000100000000100010011;
ROM[344] <= 32'b00000001010000000000001110010011;
ROM[345] <= 32'b01000000011100011000001110110011;
ROM[346] <= 32'b00000000010000111010000110000011;
ROM[347] <= 32'b00000000100000111010001000000011;
ROM[348] <= 32'b00000000110000111010001010000011;
ROM[349] <= 32'b00000001000000111010001100000011;
ROM[350] <= 32'b00000000000000001000000011100111;
ROM[351] <= 32'b00000000000000010010000000100011;
ROM[352] <= 32'b00000000010000010000000100010011;
ROM[353] <= 32'b00000000000000010010000000100011;
ROM[354] <= 32'b00000000010000010000000100010011;
ROM[355] <= 32'b00000000000000010010000000100011;
ROM[356] <= 32'b00000000010000010000000100010011;
ROM[357] <= 32'b00000000000000010010000000100011;
ROM[358] <= 32'b00000000010000010000000100010011;
ROM[359] <= 32'b00000000000000010010000000100011;
ROM[360] <= 32'b00000000010000010000000100010011;
ROM[361] <= 32'b00000000000000010010000000100011;
ROM[362] <= 32'b00000000010000010000000100010011;
ROM[363] <= 32'b00000000000000010010000000100011;
ROM[364] <= 32'b00000000010000010000000100010011;
ROM[365] <= 32'b00000000000000010010000000100011;
ROM[366] <= 32'b00000000010000010000000100010011;
ROM[367] <= 32'b00000000000000010010000000100011;
ROM[368] <= 32'b00000000010000010000000100010011;
ROM[369] <= 32'b00000000000000010010000000100011;
ROM[370] <= 32'b00000000010000010000000100010011;
ROM[371] <= 32'b00000000000000010010000000100011;
ROM[372] <= 32'b00000000010000010000000100010011;
ROM[373] <= 32'b00000000000000010010000000100011;
ROM[374] <= 32'b00000000010000010000000100010011;
ROM[375] <= 32'b00000000000000010010000000100011;
ROM[376] <= 32'b00000000010000010000000100010011;
ROM[377] <= 32'b00000000000000010010000000100011;
ROM[378] <= 32'b00000000010000010000000100010011;
ROM[379] <= 32'b00000000000000010010000000100011;
ROM[380] <= 32'b00000000010000010000000100010011;
ROM[381] <= 32'b00000000000000010010000000100011;
ROM[382] <= 32'b00000000010000010000000100010011;
ROM[383] <= 32'b00000000000000010010000000100011;
ROM[384] <= 32'b00000000010000010000000100010011;
ROM[385] <= 32'b00000000000000010010000000100011;
ROM[386] <= 32'b00000000010000010000000100010011;
ROM[387] <= 32'b00000000000000010010000000100011;
ROM[388] <= 32'b00000000010000010000000100010011;
ROM[389] <= 32'b00000000000000010010000000100011;
ROM[390] <= 32'b00000000010000010000000100010011;
ROM[391] <= 32'b00000000000000010010000000100011;
ROM[392] <= 32'b00000000010000010000000100010011;
ROM[393] <= 32'b00000000000000010010000000100011;
ROM[394] <= 32'b00000000010000010000000100010011;
ROM[395] <= 32'b00000000000000010010000000100011;
ROM[396] <= 32'b00000000010000010000000100010011;
ROM[397] <= 32'b00000000000000010010000000100011;
ROM[398] <= 32'b00000000010000010000000100010011;
ROM[399] <= 32'b00000000000000010010000000100011;
ROM[400] <= 32'b00000000010000010000000100010011;
ROM[401] <= 32'b00000000000000010010000000100011;
ROM[402] <= 32'b00000000010000010000000100010011;
ROM[403] <= 32'b00000000000000010010000000100011;
ROM[404] <= 32'b00000000010000010000000100010011;
ROM[405] <= 32'b00000000000000010010000000100011;
ROM[406] <= 32'b00000000010000010000000100010011;
ROM[407] <= 32'b00000000000000010010000000100011;
ROM[408] <= 32'b00000000010000010000000100010011;
ROM[409] <= 32'b00000000000000010010000000100011;
ROM[410] <= 32'b00000000010000010000000100010011;
ROM[411] <= 32'b00000000000000010010000000100011;
ROM[412] <= 32'b00000000010000010000000100010011;
ROM[413] <= 32'b00000000010100000000001110010011;
ROM[414] <= 32'b00000000011100010010000000100011;
ROM[415] <= 32'b00000000010000010000000100010011;
ROM[416] <= 32'b00000000000000000000001110110111;
ROM[417] <= 32'b01101100110000111000001110010011;
ROM[418] <= 32'b00000000111000111000001110110011;
ROM[419] <= 32'b00000000011100010010000000100011;
ROM[420] <= 32'b00000000010000010000000100010011;
ROM[421] <= 32'b00000000001100010010000000100011;
ROM[422] <= 32'b00000000010000010000000100010011;
ROM[423] <= 32'b00000000010000010010000000100011;
ROM[424] <= 32'b00000000010000010000000100010011;
ROM[425] <= 32'b00000000010100010010000000100011;
ROM[426] <= 32'b00000000010000010000000100010011;
ROM[427] <= 32'b00000000011000010010000000100011;
ROM[428] <= 32'b00000000010000010000000100010011;
ROM[429] <= 32'b00000001010000000000001110010011;
ROM[430] <= 32'b00000000010000111000001110010011;
ROM[431] <= 32'b01000000011100010000001110110011;
ROM[432] <= 32'b00000000011100000000001000110011;
ROM[433] <= 32'b00000000001000000000000110110011;
ROM[434] <= 32'b11010111100111111111000011101111;
ROM[435] <= 32'b11111111110000010000000100010011;
ROM[436] <= 32'b00000000000000010010001110000011;
ROM[437] <= 32'b00000000011100011010000000100011;
ROM[438] <= 32'b00000000010000000000001110010011;
ROM[439] <= 32'b00000000011100010010000000100011;
ROM[440] <= 32'b00000000010000010000000100010011;
ROM[441] <= 32'b00000000000000000000001110110111;
ROM[442] <= 32'b01110011000000111000001110010011;
ROM[443] <= 32'b00000000111000111000001110110011;
ROM[444] <= 32'b00000000011100010010000000100011;
ROM[445] <= 32'b00000000010000010000000100010011;
ROM[446] <= 32'b00000000001100010010000000100011;
ROM[447] <= 32'b00000000010000010000000100010011;
ROM[448] <= 32'b00000000010000010010000000100011;
ROM[449] <= 32'b00000000010000010000000100010011;
ROM[450] <= 32'b00000000010100010010000000100011;
ROM[451] <= 32'b00000000010000010000000100010011;
ROM[452] <= 32'b00000000011000010010000000100011;
ROM[453] <= 32'b00000000010000010000000100010011;
ROM[454] <= 32'b00000001010000000000001110010011;
ROM[455] <= 32'b00000000010000111000001110010011;
ROM[456] <= 32'b01000000011100010000001110110011;
ROM[457] <= 32'b00000000011100000000001000110011;
ROM[458] <= 32'b00000000001000000000000110110011;
ROM[459] <= 32'b00011101010000010001000011101111;
ROM[460] <= 32'b11111111110000010000000100010011;
ROM[461] <= 32'b00000000000000010010001110000011;
ROM[462] <= 32'b00000100011100011010100000100011;
ROM[463] <= 32'b00000101000000011010001110000011;
ROM[464] <= 32'b00000000011100010010000000100011;
ROM[465] <= 32'b00000000010000010000000100010011;
ROM[466] <= 32'b00000100101000000000001110010011;
ROM[467] <= 32'b00000000011100010010000000100011;
ROM[468] <= 32'b00000000010000010000000100010011;
ROM[469] <= 32'b00000000000000000000001110110111;
ROM[470] <= 32'b01111010000000111000001110010011;
ROM[471] <= 32'b00000000111000111000001110110011;
ROM[472] <= 32'b00000000011100010010000000100011;
ROM[473] <= 32'b00000000010000010000000100010011;
ROM[474] <= 32'b00000000001100010010000000100011;
ROM[475] <= 32'b00000000010000010000000100010011;
ROM[476] <= 32'b00000000010000010010000000100011;
ROM[477] <= 32'b00000000010000010000000100010011;
ROM[478] <= 32'b00000000010100010010000000100011;
ROM[479] <= 32'b00000000010000010000000100010011;
ROM[480] <= 32'b00000000011000010010000000100011;
ROM[481] <= 32'b00000000010000010000000100010011;
ROM[482] <= 32'b00000001010000000000001110010011;
ROM[483] <= 32'b00000000100000111000001110010011;
ROM[484] <= 32'b01000000011100010000001110110011;
ROM[485] <= 32'b00000000011100000000001000110011;
ROM[486] <= 32'b00000000001000000000000110110011;
ROM[487] <= 32'b01010010000000010001000011101111;
ROM[488] <= 32'b11111111110000010000000100010011;
ROM[489] <= 32'b00000000000000010010001110000011;
ROM[490] <= 32'b00000000011101100010000000100011;
ROM[491] <= 32'b00000101000000011010001110000011;
ROM[492] <= 32'b00000000011100010010000000100011;
ROM[493] <= 32'b00000000010000010000000100010011;
ROM[494] <= 32'b00000100000100000000001110010011;
ROM[495] <= 32'b00000000011100010010000000100011;
ROM[496] <= 32'b00000000010000010000000100010011;
ROM[497] <= 32'b00000000000000000001001110110111;
ROM[498] <= 32'b10000001000000111000001110010011;
ROM[499] <= 32'b00000000111000111000001110110011;
ROM[500] <= 32'b00000000011100010010000000100011;
ROM[501] <= 32'b00000000010000010000000100010011;
ROM[502] <= 32'b00000000001100010010000000100011;
ROM[503] <= 32'b00000000010000010000000100010011;
ROM[504] <= 32'b00000000010000010010000000100011;
ROM[505] <= 32'b00000000010000010000000100010011;
ROM[506] <= 32'b00000000010100010010000000100011;
ROM[507] <= 32'b00000000010000010000000100010011;
ROM[508] <= 32'b00000000011000010010000000100011;
ROM[509] <= 32'b00000000010000010000000100010011;
ROM[510] <= 32'b00000001010000000000001110010011;
ROM[511] <= 32'b00000000100000111000001110010011;
ROM[512] <= 32'b01000000011100010000001110110011;
ROM[513] <= 32'b00000000011100000000001000110011;
ROM[514] <= 32'b00000000001000000000000110110011;
ROM[515] <= 32'b01001011000000010001000011101111;
ROM[516] <= 32'b11111111110000010000000100010011;
ROM[517] <= 32'b00000000000000010010001110000011;
ROM[518] <= 32'b00000000011101100010000000100011;
ROM[519] <= 32'b00000101000000011010001110000011;
ROM[520] <= 32'b00000000011100010010000000100011;
ROM[521] <= 32'b00000000010000010000000100010011;
ROM[522] <= 32'b00000100001100000000001110010011;
ROM[523] <= 32'b00000000011100010010000000100011;
ROM[524] <= 32'b00000000010000010000000100010011;
ROM[525] <= 32'b00000000000000000001001110110111;
ROM[526] <= 32'b10001000000000111000001110010011;
ROM[527] <= 32'b00000000111000111000001110110011;
ROM[528] <= 32'b00000000011100010010000000100011;
ROM[529] <= 32'b00000000010000010000000100010011;
ROM[530] <= 32'b00000000001100010010000000100011;
ROM[531] <= 32'b00000000010000010000000100010011;
ROM[532] <= 32'b00000000010000010010000000100011;
ROM[533] <= 32'b00000000010000010000000100010011;
ROM[534] <= 32'b00000000010100010010000000100011;
ROM[535] <= 32'b00000000010000010000000100010011;
ROM[536] <= 32'b00000000011000010010000000100011;
ROM[537] <= 32'b00000000010000010000000100010011;
ROM[538] <= 32'b00000001010000000000001110010011;
ROM[539] <= 32'b00000000100000111000001110010011;
ROM[540] <= 32'b01000000011100010000001110110011;
ROM[541] <= 32'b00000000011100000000001000110011;
ROM[542] <= 32'b00000000001000000000000110110011;
ROM[543] <= 32'b01000100000000010001000011101111;
ROM[544] <= 32'b11111111110000010000000100010011;
ROM[545] <= 32'b00000000000000010010001110000011;
ROM[546] <= 32'b00000000011101100010000000100011;
ROM[547] <= 32'b00000101000000011010001110000011;
ROM[548] <= 32'b00000000011100010010000000100011;
ROM[549] <= 32'b00000000010000010000000100010011;
ROM[550] <= 32'b00000100101100000000001110010011;
ROM[551] <= 32'b00000000011100010010000000100011;
ROM[552] <= 32'b00000000010000010000000100010011;
ROM[553] <= 32'b00000000000000000001001110110111;
ROM[554] <= 32'b10001111000000111000001110010011;
ROM[555] <= 32'b00000000111000111000001110110011;
ROM[556] <= 32'b00000000011100010010000000100011;
ROM[557] <= 32'b00000000010000010000000100010011;
ROM[558] <= 32'b00000000001100010010000000100011;
ROM[559] <= 32'b00000000010000010000000100010011;
ROM[560] <= 32'b00000000010000010010000000100011;
ROM[561] <= 32'b00000000010000010000000100010011;
ROM[562] <= 32'b00000000010100010010000000100011;
ROM[563] <= 32'b00000000010000010000000100010011;
ROM[564] <= 32'b00000000011000010010000000100011;
ROM[565] <= 32'b00000000010000010000000100010011;
ROM[566] <= 32'b00000001010000000000001110010011;
ROM[567] <= 32'b00000000100000111000001110010011;
ROM[568] <= 32'b01000000011100010000001110110011;
ROM[569] <= 32'b00000000011100000000001000110011;
ROM[570] <= 32'b00000000001000000000000110110011;
ROM[571] <= 32'b00111101000000010001000011101111;
ROM[572] <= 32'b11111111110000010000000100010011;
ROM[573] <= 32'b00000000000000010010001110000011;
ROM[574] <= 32'b00000000011101100010000000100011;
ROM[575] <= 32'b00000101000000011010001110000011;
ROM[576] <= 32'b00000100011100011010100000100011;
ROM[577] <= 32'b00000000101100000000001110010011;
ROM[578] <= 32'b00000000011100010010000000100011;
ROM[579] <= 32'b00000000010000010000000100010011;
ROM[580] <= 32'b00000000000000000001001110110111;
ROM[581] <= 32'b10010101110000111000001110010011;
ROM[582] <= 32'b00000000111000111000001110110011;
ROM[583] <= 32'b00000000011100010010000000100011;
ROM[584] <= 32'b00000000010000010000000100010011;
ROM[585] <= 32'b00000000001100010010000000100011;
ROM[586] <= 32'b00000000010000010000000100010011;
ROM[587] <= 32'b00000000010000010010000000100011;
ROM[588] <= 32'b00000000010000010000000100010011;
ROM[589] <= 32'b00000000010100010010000000100011;
ROM[590] <= 32'b00000000010000010000000100010011;
ROM[591] <= 32'b00000000011000010010000000100011;
ROM[592] <= 32'b00000000010000010000000100010011;
ROM[593] <= 32'b00000001010000000000001110010011;
ROM[594] <= 32'b00000000010000111000001110010011;
ROM[595] <= 32'b01000000011100010000001110110011;
ROM[596] <= 32'b00000000011100000000001000110011;
ROM[597] <= 32'b00000000001000000000000110110011;
ROM[598] <= 32'b01111010100100010000000011101111;
ROM[599] <= 32'b11111111110000010000000100010011;
ROM[600] <= 32'b00000000000000010010001110000011;
ROM[601] <= 32'b00000100011100011010101000100011;
ROM[602] <= 32'b00000101010000011010001110000011;
ROM[603] <= 32'b00000000011100010010000000100011;
ROM[604] <= 32'b00000000010000010000000100010011;
ROM[605] <= 32'b00000101000000000000001110010011;
ROM[606] <= 32'b00000000011100010010000000100011;
ROM[607] <= 32'b00000000010000010000000100010011;
ROM[608] <= 32'b00000000000000000001001110110111;
ROM[609] <= 32'b10011100110000111000001110010011;
ROM[610] <= 32'b00000000111000111000001110110011;
ROM[611] <= 32'b00000000011100010010000000100011;
ROM[612] <= 32'b00000000010000010000000100010011;
ROM[613] <= 32'b00000000001100010010000000100011;
ROM[614] <= 32'b00000000010000010000000100010011;
ROM[615] <= 32'b00000000010000010010000000100011;
ROM[616] <= 32'b00000000010000010000000100010011;
ROM[617] <= 32'b00000000010100010010000000100011;
ROM[618] <= 32'b00000000010000010000000100010011;
ROM[619] <= 32'b00000000011000010010000000100011;
ROM[620] <= 32'b00000000010000010000000100010011;
ROM[621] <= 32'b00000001010000000000001110010011;
ROM[622] <= 32'b00000000100000111000001110010011;
ROM[623] <= 32'b01000000011100010000001110110011;
ROM[624] <= 32'b00000000011100000000001000110011;
ROM[625] <= 32'b00000000001000000000000110110011;
ROM[626] <= 32'b00101111010000010001000011101111;
ROM[627] <= 32'b11111111110000010000000100010011;
ROM[628] <= 32'b00000000000000010010001110000011;
ROM[629] <= 32'b00000000011101100010000000100011;
ROM[630] <= 32'b00000101010000011010001110000011;
ROM[631] <= 32'b00000000011100010010000000100011;
ROM[632] <= 32'b00000000010000010000000100010011;
ROM[633] <= 32'b00000101001000000000001110010011;
ROM[634] <= 32'b00000000011100010010000000100011;
ROM[635] <= 32'b00000000010000010000000100010011;
ROM[636] <= 32'b00000000000000000001001110110111;
ROM[637] <= 32'b10100011110000111000001110010011;
ROM[638] <= 32'b00000000111000111000001110110011;
ROM[639] <= 32'b00000000011100010010000000100011;
ROM[640] <= 32'b00000000010000010000000100010011;
ROM[641] <= 32'b00000000001100010010000000100011;
ROM[642] <= 32'b00000000010000010000000100010011;
ROM[643] <= 32'b00000000010000010010000000100011;
ROM[644] <= 32'b00000000010000010000000100010011;
ROM[645] <= 32'b00000000010100010010000000100011;
ROM[646] <= 32'b00000000010000010000000100010011;
ROM[647] <= 32'b00000000011000010010000000100011;
ROM[648] <= 32'b00000000010000010000000100010011;
ROM[649] <= 32'b00000001010000000000001110010011;
ROM[650] <= 32'b00000000100000111000001110010011;
ROM[651] <= 32'b01000000011100010000001110110011;
ROM[652] <= 32'b00000000011100000000001000110011;
ROM[653] <= 32'b00000000001000000000000110110011;
ROM[654] <= 32'b00101000010000010001000011101111;
ROM[655] <= 32'b11111111110000010000000100010011;
ROM[656] <= 32'b00000000000000010010001110000011;
ROM[657] <= 32'b00000000011101100010000000100011;
ROM[658] <= 32'b00000101010000011010001110000011;
ROM[659] <= 32'b00000000011100010010000000100011;
ROM[660] <= 32'b00000000010000010000000100010011;
ROM[661] <= 32'b00000100111100000000001110010011;
ROM[662] <= 32'b00000000011100010010000000100011;
ROM[663] <= 32'b00000000010000010000000100010011;
ROM[664] <= 32'b00000000000000000001001110110111;
ROM[665] <= 32'b10101010110000111000001110010011;
ROM[666] <= 32'b00000000111000111000001110110011;
ROM[667] <= 32'b00000000011100010010000000100011;
ROM[668] <= 32'b00000000010000010000000100010011;
ROM[669] <= 32'b00000000001100010010000000100011;
ROM[670] <= 32'b00000000010000010000000100010011;
ROM[671] <= 32'b00000000010000010010000000100011;
ROM[672] <= 32'b00000000010000010000000100010011;
ROM[673] <= 32'b00000000010100010010000000100011;
ROM[674] <= 32'b00000000010000010000000100010011;
ROM[675] <= 32'b00000000011000010010000000100011;
ROM[676] <= 32'b00000000010000010000000100010011;
ROM[677] <= 32'b00000001010000000000001110010011;
ROM[678] <= 32'b00000000100000111000001110010011;
ROM[679] <= 32'b01000000011100010000001110110011;
ROM[680] <= 32'b00000000011100000000001000110011;
ROM[681] <= 32'b00000000001000000000000110110011;
ROM[682] <= 32'b00100001010000010001000011101111;
ROM[683] <= 32'b11111111110000010000000100010011;
ROM[684] <= 32'b00000000000000010010001110000011;
ROM[685] <= 32'b00000000011101100010000000100011;
ROM[686] <= 32'b00000101010000011010001110000011;
ROM[687] <= 32'b00000000011100010010000000100011;
ROM[688] <= 32'b00000000010000010000000100010011;
ROM[689] <= 32'b00000100011100000000001110010011;
ROM[690] <= 32'b00000000011100010010000000100011;
ROM[691] <= 32'b00000000010000010000000100010011;
ROM[692] <= 32'b00000000000000000001001110110111;
ROM[693] <= 32'b10110001110000111000001110010011;
ROM[694] <= 32'b00000000111000111000001110110011;
ROM[695] <= 32'b00000000011100010010000000100011;
ROM[696] <= 32'b00000000010000010000000100010011;
ROM[697] <= 32'b00000000001100010010000000100011;
ROM[698] <= 32'b00000000010000010000000100010011;
ROM[699] <= 32'b00000000010000010010000000100011;
ROM[700] <= 32'b00000000010000010000000100010011;
ROM[701] <= 32'b00000000010100010010000000100011;
ROM[702] <= 32'b00000000010000010000000100010011;
ROM[703] <= 32'b00000000011000010010000000100011;
ROM[704] <= 32'b00000000010000010000000100010011;
ROM[705] <= 32'b00000001010000000000001110010011;
ROM[706] <= 32'b00000000100000111000001110010011;
ROM[707] <= 32'b01000000011100010000001110110011;
ROM[708] <= 32'b00000000011100000000001000110011;
ROM[709] <= 32'b00000000001000000000000110110011;
ROM[710] <= 32'b00011010010000010001000011101111;
ROM[711] <= 32'b11111111110000010000000100010011;
ROM[712] <= 32'b00000000000000010010001110000011;
ROM[713] <= 32'b00000000011101100010000000100011;
ROM[714] <= 32'b00000101010000011010001110000011;
ROM[715] <= 32'b00000000011100010010000000100011;
ROM[716] <= 32'b00000000010000010000000100010011;
ROM[717] <= 32'b00000101001000000000001110010011;
ROM[718] <= 32'b00000000011100010010000000100011;
ROM[719] <= 32'b00000000010000010000000100010011;
ROM[720] <= 32'b00000000000000000001001110110111;
ROM[721] <= 32'b10111000110000111000001110010011;
ROM[722] <= 32'b00000000111000111000001110110011;
ROM[723] <= 32'b00000000011100010010000000100011;
ROM[724] <= 32'b00000000010000010000000100010011;
ROM[725] <= 32'b00000000001100010010000000100011;
ROM[726] <= 32'b00000000010000010000000100010011;
ROM[727] <= 32'b00000000010000010010000000100011;
ROM[728] <= 32'b00000000010000010000000100010011;
ROM[729] <= 32'b00000000010100010010000000100011;
ROM[730] <= 32'b00000000010000010000000100010011;
ROM[731] <= 32'b00000000011000010010000000100011;
ROM[732] <= 32'b00000000010000010000000100010011;
ROM[733] <= 32'b00000001010000000000001110010011;
ROM[734] <= 32'b00000000100000111000001110010011;
ROM[735] <= 32'b01000000011100010000001110110011;
ROM[736] <= 32'b00000000011100000000001000110011;
ROM[737] <= 32'b00000000001000000000000110110011;
ROM[738] <= 32'b00010011010000010001000011101111;
ROM[739] <= 32'b11111111110000010000000100010011;
ROM[740] <= 32'b00000000000000010010001110000011;
ROM[741] <= 32'b00000000011101100010000000100011;
ROM[742] <= 32'b00000101010000011010001110000011;
ROM[743] <= 32'b00000000011100010010000000100011;
ROM[744] <= 32'b00000000010000010000000100010011;
ROM[745] <= 32'b00000100000100000000001110010011;
ROM[746] <= 32'b00000000011100010010000000100011;
ROM[747] <= 32'b00000000010000010000000100010011;
ROM[748] <= 32'b00000000000000000001001110110111;
ROM[749] <= 32'b10111111110000111000001110010011;
ROM[750] <= 32'b00000000111000111000001110110011;
ROM[751] <= 32'b00000000011100010010000000100011;
ROM[752] <= 32'b00000000010000010000000100010011;
ROM[753] <= 32'b00000000001100010010000000100011;
ROM[754] <= 32'b00000000010000010000000100010011;
ROM[755] <= 32'b00000000010000010010000000100011;
ROM[756] <= 32'b00000000010000010000000100010011;
ROM[757] <= 32'b00000000010100010010000000100011;
ROM[758] <= 32'b00000000010000010000000100010011;
ROM[759] <= 32'b00000000011000010010000000100011;
ROM[760] <= 32'b00000000010000010000000100010011;
ROM[761] <= 32'b00000001010000000000001110010011;
ROM[762] <= 32'b00000000100000111000001110010011;
ROM[763] <= 32'b01000000011100010000001110110011;
ROM[764] <= 32'b00000000011100000000001000110011;
ROM[765] <= 32'b00000000001000000000000110110011;
ROM[766] <= 32'b00001100010000010001000011101111;
ROM[767] <= 32'b11111111110000010000000100010011;
ROM[768] <= 32'b00000000000000010010001110000011;
ROM[769] <= 32'b00000000011101100010000000100011;
ROM[770] <= 32'b00000101010000011010001110000011;
ROM[771] <= 32'b00000000011100010010000000100011;
ROM[772] <= 32'b00000000010000010000000100010011;
ROM[773] <= 32'b00000100110100000000001110010011;
ROM[774] <= 32'b00000000011100010010000000100011;
ROM[775] <= 32'b00000000010000010000000100010011;
ROM[776] <= 32'b00000000000000000001001110110111;
ROM[777] <= 32'b11000110110000111000001110010011;
ROM[778] <= 32'b00000000111000111000001110110011;
ROM[779] <= 32'b00000000011100010010000000100011;
ROM[780] <= 32'b00000000010000010000000100010011;
ROM[781] <= 32'b00000000001100010010000000100011;
ROM[782] <= 32'b00000000010000010000000100010011;
ROM[783] <= 32'b00000000010000010010000000100011;
ROM[784] <= 32'b00000000010000010000000100010011;
ROM[785] <= 32'b00000000010100010010000000100011;
ROM[786] <= 32'b00000000010000010000000100010011;
ROM[787] <= 32'b00000000011000010010000000100011;
ROM[788] <= 32'b00000000010000010000000100010011;
ROM[789] <= 32'b00000001010000000000001110010011;
ROM[790] <= 32'b00000000100000111000001110010011;
ROM[791] <= 32'b01000000011100010000001110110011;
ROM[792] <= 32'b00000000011100000000001000110011;
ROM[793] <= 32'b00000000001000000000000110110011;
ROM[794] <= 32'b00000101010000010001000011101111;
ROM[795] <= 32'b11111111110000010000000100010011;
ROM[796] <= 32'b00000000000000010010001110000011;
ROM[797] <= 32'b00000000011101100010000000100011;
ROM[798] <= 32'b00000101010000011010001110000011;
ROM[799] <= 32'b00000000011100010010000000100011;
ROM[800] <= 32'b00000000010000010000000100010011;
ROM[801] <= 32'b00000100110100000000001110010011;
ROM[802] <= 32'b00000000011100010010000000100011;
ROM[803] <= 32'b00000000010000010000000100010011;
ROM[804] <= 32'b00000000000000000001001110110111;
ROM[805] <= 32'b11001101110000111000001110010011;
ROM[806] <= 32'b00000000111000111000001110110011;
ROM[807] <= 32'b00000000011100010010000000100011;
ROM[808] <= 32'b00000000010000010000000100010011;
ROM[809] <= 32'b00000000001100010010000000100011;
ROM[810] <= 32'b00000000010000010000000100010011;
ROM[811] <= 32'b00000000010000010010000000100011;
ROM[812] <= 32'b00000000010000010000000100010011;
ROM[813] <= 32'b00000000010100010010000000100011;
ROM[814] <= 32'b00000000010000010000000100010011;
ROM[815] <= 32'b00000000011000010010000000100011;
ROM[816] <= 32'b00000000010000010000000100010011;
ROM[817] <= 32'b00000001010000000000001110010011;
ROM[818] <= 32'b00000000100000111000001110010011;
ROM[819] <= 32'b01000000011100010000001110110011;
ROM[820] <= 32'b00000000011100000000001000110011;
ROM[821] <= 32'b00000000001000000000000110110011;
ROM[822] <= 32'b01111110010100010000000011101111;
ROM[823] <= 32'b11111111110000010000000100010011;
ROM[824] <= 32'b00000000000000010010001110000011;
ROM[825] <= 32'b00000000011101100010000000100011;
ROM[826] <= 32'b00000101010000011010001110000011;
ROM[827] <= 32'b00000000011100010010000000100011;
ROM[828] <= 32'b00000000010000010000000100010011;
ROM[829] <= 32'b00000100100100000000001110010011;
ROM[830] <= 32'b00000000011100010010000000100011;
ROM[831] <= 32'b00000000010000010000000100010011;
ROM[832] <= 32'b00000000000000000001001110110111;
ROM[833] <= 32'b11010100110000111000001110010011;
ROM[834] <= 32'b00000000111000111000001110110011;
ROM[835] <= 32'b00000000011100010010000000100011;
ROM[836] <= 32'b00000000010000010000000100010011;
ROM[837] <= 32'b00000000001100010010000000100011;
ROM[838] <= 32'b00000000010000010000000100010011;
ROM[839] <= 32'b00000000010000010010000000100011;
ROM[840] <= 32'b00000000010000010000000100010011;
ROM[841] <= 32'b00000000010100010010000000100011;
ROM[842] <= 32'b00000000010000010000000100010011;
ROM[843] <= 32'b00000000011000010010000000100011;
ROM[844] <= 32'b00000000010000010000000100010011;
ROM[845] <= 32'b00000001010000000000001110010011;
ROM[846] <= 32'b00000000100000111000001110010011;
ROM[847] <= 32'b01000000011100010000001110110011;
ROM[848] <= 32'b00000000011100000000001000110011;
ROM[849] <= 32'b00000000001000000000000110110011;
ROM[850] <= 32'b01110111010100010000000011101111;
ROM[851] <= 32'b11111111110000010000000100010011;
ROM[852] <= 32'b00000000000000010010001110000011;
ROM[853] <= 32'b00000000011101100010000000100011;
ROM[854] <= 32'b00000101010000011010001110000011;
ROM[855] <= 32'b00000000011100010010000000100011;
ROM[856] <= 32'b00000000010000010000000100010011;
ROM[857] <= 32'b00000100111000000000001110010011;
ROM[858] <= 32'b00000000011100010010000000100011;
ROM[859] <= 32'b00000000010000010000000100010011;
ROM[860] <= 32'b00000000000000000001001110110111;
ROM[861] <= 32'b11011011110000111000001110010011;
ROM[862] <= 32'b00000000111000111000001110110011;
ROM[863] <= 32'b00000000011100010010000000100011;
ROM[864] <= 32'b00000000010000010000000100010011;
ROM[865] <= 32'b00000000001100010010000000100011;
ROM[866] <= 32'b00000000010000010000000100010011;
ROM[867] <= 32'b00000000010000010010000000100011;
ROM[868] <= 32'b00000000010000010000000100010011;
ROM[869] <= 32'b00000000010100010010000000100011;
ROM[870] <= 32'b00000000010000010000000100010011;
ROM[871] <= 32'b00000000011000010010000000100011;
ROM[872] <= 32'b00000000010000010000000100010011;
ROM[873] <= 32'b00000001010000000000001110010011;
ROM[874] <= 32'b00000000100000111000001110010011;
ROM[875] <= 32'b01000000011100010000001110110011;
ROM[876] <= 32'b00000000011100000000001000110011;
ROM[877] <= 32'b00000000001000000000000110110011;
ROM[878] <= 32'b01110000010100010000000011101111;
ROM[879] <= 32'b11111111110000010000000100010011;
ROM[880] <= 32'b00000000000000010010001110000011;
ROM[881] <= 32'b00000000011101100010000000100011;
ROM[882] <= 32'b00000101010000011010001110000011;
ROM[883] <= 32'b00000000011100010010000000100011;
ROM[884] <= 32'b00000000010000010000000100010011;
ROM[885] <= 32'b00000100011100000000001110010011;
ROM[886] <= 32'b00000000011100010010000000100011;
ROM[887] <= 32'b00000000010000010000000100010011;
ROM[888] <= 32'b00000000000000000001001110110111;
ROM[889] <= 32'b11100010110000111000001110010011;
ROM[890] <= 32'b00000000111000111000001110110011;
ROM[891] <= 32'b00000000011100010010000000100011;
ROM[892] <= 32'b00000000010000010000000100010011;
ROM[893] <= 32'b00000000001100010010000000100011;
ROM[894] <= 32'b00000000010000010000000100010011;
ROM[895] <= 32'b00000000010000010010000000100011;
ROM[896] <= 32'b00000000010000010000000100010011;
ROM[897] <= 32'b00000000010100010010000000100011;
ROM[898] <= 32'b00000000010000010000000100010011;
ROM[899] <= 32'b00000000011000010010000000100011;
ROM[900] <= 32'b00000000010000010000000100010011;
ROM[901] <= 32'b00000001010000000000001110010011;
ROM[902] <= 32'b00000000100000111000001110010011;
ROM[903] <= 32'b01000000011100010000001110110011;
ROM[904] <= 32'b00000000011100000000001000110011;
ROM[905] <= 32'b00000000001000000000000110110011;
ROM[906] <= 32'b01101001010100010000000011101111;
ROM[907] <= 32'b11111111110000010000000100010011;
ROM[908] <= 32'b00000000000000010010001110000011;
ROM[909] <= 32'b00000000011101100010000000100011;
ROM[910] <= 32'b00000101010000011010001110000011;
ROM[911] <= 32'b00000100011100011010101000100011;
ROM[912] <= 32'b00000000100000000000001110010011;
ROM[913] <= 32'b00000000011100010010000000100011;
ROM[914] <= 32'b00000000010000010000000100010011;
ROM[915] <= 32'b00000000000000000001001110110111;
ROM[916] <= 32'b11101001100000111000001110010011;
ROM[917] <= 32'b00000000111000111000001110110011;
ROM[918] <= 32'b00000000011100010010000000100011;
ROM[919] <= 32'b00000000010000010000000100010011;
ROM[920] <= 32'b00000000001100010010000000100011;
ROM[921] <= 32'b00000000010000010000000100010011;
ROM[922] <= 32'b00000000010000010010000000100011;
ROM[923] <= 32'b00000000010000010000000100010011;
ROM[924] <= 32'b00000000010100010010000000100011;
ROM[925] <= 32'b00000000010000010000000100010011;
ROM[926] <= 32'b00000000011000010010000000100011;
ROM[927] <= 32'b00000000010000010000000100010011;
ROM[928] <= 32'b00000001010000000000001110010011;
ROM[929] <= 32'b00000000010000111000001110010011;
ROM[930] <= 32'b01000000011100010000001110110011;
ROM[931] <= 32'b00000000011100000000001000110011;
ROM[932] <= 32'b00000000001000000000000110110011;
ROM[933] <= 32'b00100110110100010000000011101111;
ROM[934] <= 32'b11111111110000010000000100010011;
ROM[935] <= 32'b00000000000000010010001110000011;
ROM[936] <= 32'b00000100011100011010110000100011;
ROM[937] <= 32'b00000101100000011010001110000011;
ROM[938] <= 32'b00000000011100010010000000100011;
ROM[939] <= 32'b00000000010000010000000100010011;
ROM[940] <= 32'b00000100110000000000001110010011;
ROM[941] <= 32'b00000000011100010010000000100011;
ROM[942] <= 32'b00000000010000010000000100010011;
ROM[943] <= 32'b00000000000000000001001110110111;
ROM[944] <= 32'b11110000100000111000001110010011;
ROM[945] <= 32'b00000000111000111000001110110011;
ROM[946] <= 32'b00000000011100010010000000100011;
ROM[947] <= 32'b00000000010000010000000100010011;
ROM[948] <= 32'b00000000001100010010000000100011;
ROM[949] <= 32'b00000000010000010000000100010011;
ROM[950] <= 32'b00000000010000010010000000100011;
ROM[951] <= 32'b00000000010000010000000100010011;
ROM[952] <= 32'b00000000010100010010000000100011;
ROM[953] <= 32'b00000000010000010000000100010011;
ROM[954] <= 32'b00000000011000010010000000100011;
ROM[955] <= 32'b00000000010000010000000100010011;
ROM[956] <= 32'b00000001010000000000001110010011;
ROM[957] <= 32'b00000000100000111000001110010011;
ROM[958] <= 32'b01000000011100010000001110110011;
ROM[959] <= 32'b00000000011100000000001000110011;
ROM[960] <= 32'b00000000001000000000000110110011;
ROM[961] <= 32'b01011011100100010000000011101111;
ROM[962] <= 32'b11111111110000010000000100010011;
ROM[963] <= 32'b00000000000000010010001110000011;
ROM[964] <= 32'b00000000011101100010000000100011;
ROM[965] <= 32'b00000101100000011010001110000011;
ROM[966] <= 32'b00000000011100010010000000100011;
ROM[967] <= 32'b00000000010000010000000100010011;
ROM[968] <= 32'b00000100000100000000001110010011;
ROM[969] <= 32'b00000000011100010010000000100011;
ROM[970] <= 32'b00000000010000010000000100010011;
ROM[971] <= 32'b00000000000000000001001110110111;
ROM[972] <= 32'b11110111100000111000001110010011;
ROM[973] <= 32'b00000000111000111000001110110011;
ROM[974] <= 32'b00000000011100010010000000100011;
ROM[975] <= 32'b00000000010000010000000100010011;
ROM[976] <= 32'b00000000001100010010000000100011;
ROM[977] <= 32'b00000000010000010000000100010011;
ROM[978] <= 32'b00000000010000010010000000100011;
ROM[979] <= 32'b00000000010000010000000100010011;
ROM[980] <= 32'b00000000010100010010000000100011;
ROM[981] <= 32'b00000000010000010000000100010011;
ROM[982] <= 32'b00000000011000010010000000100011;
ROM[983] <= 32'b00000000010000010000000100010011;
ROM[984] <= 32'b00000001010000000000001110010011;
ROM[985] <= 32'b00000000100000111000001110010011;
ROM[986] <= 32'b01000000011100010000001110110011;
ROM[987] <= 32'b00000000011100000000001000110011;
ROM[988] <= 32'b00000000001000000000000110110011;
ROM[989] <= 32'b01010100100100010000000011101111;
ROM[990] <= 32'b11111111110000010000000100010011;
ROM[991] <= 32'b00000000000000010010001110000011;
ROM[992] <= 32'b00000000011101100010000000100011;
ROM[993] <= 32'b00000101100000011010001110000011;
ROM[994] <= 32'b00000000011100010010000000100011;
ROM[995] <= 32'b00000000010000010000000100010011;
ROM[996] <= 32'b00000100111000000000001110010011;
ROM[997] <= 32'b00000000011100010010000000100011;
ROM[998] <= 32'b00000000010000010000000100010011;
ROM[999] <= 32'b00000000000000000001001110110111;
ROM[1000] <= 32'b11111110100000111000001110010011;
ROM[1001] <= 32'b00000000111000111000001110110011;
ROM[1002] <= 32'b00000000011100010010000000100011;
ROM[1003] <= 32'b00000000010000010000000100010011;
ROM[1004] <= 32'b00000000001100010010000000100011;
ROM[1005] <= 32'b00000000010000010000000100010011;
ROM[1006] <= 32'b00000000010000010010000000100011;
ROM[1007] <= 32'b00000000010000010000000100010011;
ROM[1008] <= 32'b00000000010100010010000000100011;
ROM[1009] <= 32'b00000000010000010000000100010011;
ROM[1010] <= 32'b00000000011000010010000000100011;
ROM[1011] <= 32'b00000000010000010000000100010011;
ROM[1012] <= 32'b00000001010000000000001110010011;
ROM[1013] <= 32'b00000000100000111000001110010011;
ROM[1014] <= 32'b01000000011100010000001110110011;
ROM[1015] <= 32'b00000000011100000000001000110011;
ROM[1016] <= 32'b00000000001000000000000110110011;
ROM[1017] <= 32'b01001101100100010000000011101111;
ROM[1018] <= 32'b11111111110000010000000100010011;
ROM[1019] <= 32'b00000000000000010010001110000011;
ROM[1020] <= 32'b00000000011101100010000000100011;
ROM[1021] <= 32'b00000101100000011010001110000011;
ROM[1022] <= 32'b00000000011100010010000000100011;
ROM[1023] <= 32'b00000000010000010000000100010011;
ROM[1024] <= 32'b00000100011100000000001110010011;
ROM[1025] <= 32'b00000000011100010010000000100011;
ROM[1026] <= 32'b00000000010000010000000100010011;
ROM[1027] <= 32'b00000000000000000001001110110111;
ROM[1028] <= 32'b00000101100000111000001110010011;
ROM[1029] <= 32'b00000000111000111000001110110011;
ROM[1030] <= 32'b00000000011100010010000000100011;
ROM[1031] <= 32'b00000000010000010000000100010011;
ROM[1032] <= 32'b00000000001100010010000000100011;
ROM[1033] <= 32'b00000000010000010000000100010011;
ROM[1034] <= 32'b00000000010000010010000000100011;
ROM[1035] <= 32'b00000000010000010000000100010011;
ROM[1036] <= 32'b00000000010100010010000000100011;
ROM[1037] <= 32'b00000000010000010000000100010011;
ROM[1038] <= 32'b00000000011000010010000000100011;
ROM[1039] <= 32'b00000000010000010000000100010011;
ROM[1040] <= 32'b00000001010000000000001110010011;
ROM[1041] <= 32'b00000000100000111000001110010011;
ROM[1042] <= 32'b01000000011100010000001110110011;
ROM[1043] <= 32'b00000000011100000000001000110011;
ROM[1044] <= 32'b00000000001000000000000110110011;
ROM[1045] <= 32'b01000110100100010000000011101111;
ROM[1046] <= 32'b11111111110000010000000100010011;
ROM[1047] <= 32'b00000000000000010010001110000011;
ROM[1048] <= 32'b00000000011101100010000000100011;
ROM[1049] <= 32'b00000101100000011010001110000011;
ROM[1050] <= 32'b00000000011100010010000000100011;
ROM[1051] <= 32'b00000000010000010000000100010011;
ROM[1052] <= 32'b00000101010100000000001110010011;
ROM[1053] <= 32'b00000000011100010010000000100011;
ROM[1054] <= 32'b00000000010000010000000100010011;
ROM[1055] <= 32'b00000000000000000001001110110111;
ROM[1056] <= 32'b00001100100000111000001110010011;
ROM[1057] <= 32'b00000000111000111000001110110011;
ROM[1058] <= 32'b00000000011100010010000000100011;
ROM[1059] <= 32'b00000000010000010000000100010011;
ROM[1060] <= 32'b00000000001100010010000000100011;
ROM[1061] <= 32'b00000000010000010000000100010011;
ROM[1062] <= 32'b00000000010000010010000000100011;
ROM[1063] <= 32'b00000000010000010000000100010011;
ROM[1064] <= 32'b00000000010100010010000000100011;
ROM[1065] <= 32'b00000000010000010000000100010011;
ROM[1066] <= 32'b00000000011000010010000000100011;
ROM[1067] <= 32'b00000000010000010000000100010011;
ROM[1068] <= 32'b00000001010000000000001110010011;
ROM[1069] <= 32'b00000000100000111000001110010011;
ROM[1070] <= 32'b01000000011100010000001110110011;
ROM[1071] <= 32'b00000000011100000000001000110011;
ROM[1072] <= 32'b00000000001000000000000110110011;
ROM[1073] <= 32'b00111111100100010000000011101111;
ROM[1074] <= 32'b11111111110000010000000100010011;
ROM[1075] <= 32'b00000000000000010010001110000011;
ROM[1076] <= 32'b00000000011101100010000000100011;
ROM[1077] <= 32'b00000101100000011010001110000011;
ROM[1078] <= 32'b00000000011100010010000000100011;
ROM[1079] <= 32'b00000000010000010000000100010011;
ROM[1080] <= 32'b00000100000100000000001110010011;
ROM[1081] <= 32'b00000000011100010010000000100011;
ROM[1082] <= 32'b00000000010000010000000100010011;
ROM[1083] <= 32'b00000000000000000001001110110111;
ROM[1084] <= 32'b00010011100000111000001110010011;
ROM[1085] <= 32'b00000000111000111000001110110011;
ROM[1086] <= 32'b00000000011100010010000000100011;
ROM[1087] <= 32'b00000000010000010000000100010011;
ROM[1088] <= 32'b00000000001100010010000000100011;
ROM[1089] <= 32'b00000000010000010000000100010011;
ROM[1090] <= 32'b00000000010000010010000000100011;
ROM[1091] <= 32'b00000000010000010000000100010011;
ROM[1092] <= 32'b00000000010100010010000000100011;
ROM[1093] <= 32'b00000000010000010000000100010011;
ROM[1094] <= 32'b00000000011000010010000000100011;
ROM[1095] <= 32'b00000000010000010000000100010011;
ROM[1096] <= 32'b00000001010000000000001110010011;
ROM[1097] <= 32'b00000000100000111000001110010011;
ROM[1098] <= 32'b01000000011100010000001110110011;
ROM[1099] <= 32'b00000000011100000000001000110011;
ROM[1100] <= 32'b00000000001000000000000110110011;
ROM[1101] <= 32'b00111000100100010000000011101111;
ROM[1102] <= 32'b11111111110000010000000100010011;
ROM[1103] <= 32'b00000000000000010010001110000011;
ROM[1104] <= 32'b00000000011101100010000000100011;
ROM[1105] <= 32'b00000101100000011010001110000011;
ROM[1106] <= 32'b00000000011100010010000000100011;
ROM[1107] <= 32'b00000000010000010000000100010011;
ROM[1108] <= 32'b00000100011100000000001110010011;
ROM[1109] <= 32'b00000000011100010010000000100011;
ROM[1110] <= 32'b00000000010000010000000100010011;
ROM[1111] <= 32'b00000000000000000001001110110111;
ROM[1112] <= 32'b00011010100000111000001110010011;
ROM[1113] <= 32'b00000000111000111000001110110011;
ROM[1114] <= 32'b00000000011100010010000000100011;
ROM[1115] <= 32'b00000000010000010000000100010011;
ROM[1116] <= 32'b00000000001100010010000000100011;
ROM[1117] <= 32'b00000000010000010000000100010011;
ROM[1118] <= 32'b00000000010000010010000000100011;
ROM[1119] <= 32'b00000000010000010000000100010011;
ROM[1120] <= 32'b00000000010100010010000000100011;
ROM[1121] <= 32'b00000000010000010000000100010011;
ROM[1122] <= 32'b00000000011000010010000000100011;
ROM[1123] <= 32'b00000000010000010000000100010011;
ROM[1124] <= 32'b00000001010000000000001110010011;
ROM[1125] <= 32'b00000000100000111000001110010011;
ROM[1126] <= 32'b01000000011100010000001110110011;
ROM[1127] <= 32'b00000000011100000000001000110011;
ROM[1128] <= 32'b00000000001000000000000110110011;
ROM[1129] <= 32'b00110001100100010000000011101111;
ROM[1130] <= 32'b11111111110000010000000100010011;
ROM[1131] <= 32'b00000000000000010010001110000011;
ROM[1132] <= 32'b00000000011101100010000000100011;
ROM[1133] <= 32'b00000101100000011010001110000011;
ROM[1134] <= 32'b00000000011100010010000000100011;
ROM[1135] <= 32'b00000000010000010000000100010011;
ROM[1136] <= 32'b00000100010100000000001110010011;
ROM[1137] <= 32'b00000000011100010010000000100011;
ROM[1138] <= 32'b00000000010000010000000100010011;
ROM[1139] <= 32'b00000000000000000001001110110111;
ROM[1140] <= 32'b00100001100000111000001110010011;
ROM[1141] <= 32'b00000000111000111000001110110011;
ROM[1142] <= 32'b00000000011100010010000000100011;
ROM[1143] <= 32'b00000000010000010000000100010011;
ROM[1144] <= 32'b00000000001100010010000000100011;
ROM[1145] <= 32'b00000000010000010000000100010011;
ROM[1146] <= 32'b00000000010000010010000000100011;
ROM[1147] <= 32'b00000000010000010000000100010011;
ROM[1148] <= 32'b00000000010100010010000000100011;
ROM[1149] <= 32'b00000000010000010000000100010011;
ROM[1150] <= 32'b00000000011000010010000000100011;
ROM[1151] <= 32'b00000000010000010000000100010011;
ROM[1152] <= 32'b00000001010000000000001110010011;
ROM[1153] <= 32'b00000000100000111000001110010011;
ROM[1154] <= 32'b01000000011100010000001110110011;
ROM[1155] <= 32'b00000000011100000000001000110011;
ROM[1156] <= 32'b00000000001000000000000110110011;
ROM[1157] <= 32'b00101010100100010000000011101111;
ROM[1158] <= 32'b11111111110000010000000100010011;
ROM[1159] <= 32'b00000000000000010010001110000011;
ROM[1160] <= 32'b00000000011101100010000000100011;
ROM[1161] <= 32'b00000101100000011010001110000011;
ROM[1162] <= 32'b00000100011100011010110000100011;
ROM[1163] <= 32'b00000000100000000000001110010011;
ROM[1164] <= 32'b00000000011100010010000000100011;
ROM[1165] <= 32'b00000000010000010000000100010011;
ROM[1166] <= 32'b00000000000000000001001110110111;
ROM[1167] <= 32'b00101000010000111000001110010011;
ROM[1168] <= 32'b00000000111000111000001110110011;
ROM[1169] <= 32'b00000000011100010010000000100011;
ROM[1170] <= 32'b00000000010000010000000100010011;
ROM[1171] <= 32'b00000000001100010010000000100011;
ROM[1172] <= 32'b00000000010000010000000100010011;
ROM[1173] <= 32'b00000000010000010010000000100011;
ROM[1174] <= 32'b00000000010000010000000100010011;
ROM[1175] <= 32'b00000000010100010010000000100011;
ROM[1176] <= 32'b00000000010000010000000100010011;
ROM[1177] <= 32'b00000000011000010010000000100011;
ROM[1178] <= 32'b00000000010000010000000100010011;
ROM[1179] <= 32'b00000001010000000000001110010011;
ROM[1180] <= 32'b00000000010000111000001110010011;
ROM[1181] <= 32'b01000000011100010000001110110011;
ROM[1182] <= 32'b00000000011100000000001000110011;
ROM[1183] <= 32'b00000000001000000000000110110011;
ROM[1184] <= 32'b01101000000000010000000011101111;
ROM[1185] <= 32'b11111111110000010000000100010011;
ROM[1186] <= 32'b00000000000000010010001110000011;
ROM[1187] <= 32'b00000100011100011010111000100011;
ROM[1188] <= 32'b00000101110000011010001110000011;
ROM[1189] <= 32'b00000000011100010010000000100011;
ROM[1190] <= 32'b00000000010000010000000100010011;
ROM[1191] <= 32'b00000100001100000000001110010011;
ROM[1192] <= 32'b00000000011100010010000000100011;
ROM[1193] <= 32'b00000000010000010000000100010011;
ROM[1194] <= 32'b00000000000000000001001110110111;
ROM[1195] <= 32'b00101111010000111000001110010011;
ROM[1196] <= 32'b00000000111000111000001110110011;
ROM[1197] <= 32'b00000000011100010010000000100011;
ROM[1198] <= 32'b00000000010000010000000100010011;
ROM[1199] <= 32'b00000000001100010010000000100011;
ROM[1200] <= 32'b00000000010000010000000100010011;
ROM[1201] <= 32'b00000000010000010010000000100011;
ROM[1202] <= 32'b00000000010000010000000100010011;
ROM[1203] <= 32'b00000000010100010010000000100011;
ROM[1204] <= 32'b00000000010000010000000100010011;
ROM[1205] <= 32'b00000000011000010010000000100011;
ROM[1206] <= 32'b00000000010000010000000100010011;
ROM[1207] <= 32'b00000001010000000000001110010011;
ROM[1208] <= 32'b00000000100000111000001110010011;
ROM[1209] <= 32'b01000000011100010000001110110011;
ROM[1210] <= 32'b00000000011100000000001000110011;
ROM[1211] <= 32'b00000000001000000000000110110011;
ROM[1212] <= 32'b00011100110100010000000011101111;
ROM[1213] <= 32'b11111111110000010000000100010011;
ROM[1214] <= 32'b00000000000000010010001110000011;
ROM[1215] <= 32'b00000000011101100010000000100011;
ROM[1216] <= 32'b00000101110000011010001110000011;
ROM[1217] <= 32'b00000000011100010010000000100011;
ROM[1218] <= 32'b00000000010000010000000100010011;
ROM[1219] <= 32'b00000100111100000000001110010011;
ROM[1220] <= 32'b00000000011100010010000000100011;
ROM[1221] <= 32'b00000000010000010000000100010011;
ROM[1222] <= 32'b00000000000000000001001110110111;
ROM[1223] <= 32'b00110110010000111000001110010011;
ROM[1224] <= 32'b00000000111000111000001110110011;
ROM[1225] <= 32'b00000000011100010010000000100011;
ROM[1226] <= 32'b00000000010000010000000100010011;
ROM[1227] <= 32'b00000000001100010010000000100011;
ROM[1228] <= 32'b00000000010000010000000100010011;
ROM[1229] <= 32'b00000000010000010010000000100011;
ROM[1230] <= 32'b00000000010000010000000100010011;
ROM[1231] <= 32'b00000000010100010010000000100011;
ROM[1232] <= 32'b00000000010000010000000100010011;
ROM[1233] <= 32'b00000000011000010010000000100011;
ROM[1234] <= 32'b00000000010000010000000100010011;
ROM[1235] <= 32'b00000001010000000000001110010011;
ROM[1236] <= 32'b00000000100000111000001110010011;
ROM[1237] <= 32'b01000000011100010000001110110011;
ROM[1238] <= 32'b00000000011100000000001000110011;
ROM[1239] <= 32'b00000000001000000000000110110011;
ROM[1240] <= 32'b00010101110100010000000011101111;
ROM[1241] <= 32'b11111111110000010000000100010011;
ROM[1242] <= 32'b00000000000000010010001110000011;
ROM[1243] <= 32'b00000000011101100010000000100011;
ROM[1244] <= 32'b00000101110000011010001110000011;
ROM[1245] <= 32'b00000000011100010010000000100011;
ROM[1246] <= 32'b00000000010000010000000100010011;
ROM[1247] <= 32'b00000100110100000000001110010011;
ROM[1248] <= 32'b00000000011100010010000000100011;
ROM[1249] <= 32'b00000000010000010000000100010011;
ROM[1250] <= 32'b00000000000000000001001110110111;
ROM[1251] <= 32'b00111101010000111000001110010011;
ROM[1252] <= 32'b00000000111000111000001110110011;
ROM[1253] <= 32'b00000000011100010010000000100011;
ROM[1254] <= 32'b00000000010000010000000100010011;
ROM[1255] <= 32'b00000000001100010010000000100011;
ROM[1256] <= 32'b00000000010000010000000100010011;
ROM[1257] <= 32'b00000000010000010010000000100011;
ROM[1258] <= 32'b00000000010000010000000100010011;
ROM[1259] <= 32'b00000000010100010010000000100011;
ROM[1260] <= 32'b00000000010000010000000100010011;
ROM[1261] <= 32'b00000000011000010010000000100011;
ROM[1262] <= 32'b00000000010000010000000100010011;
ROM[1263] <= 32'b00000001010000000000001110010011;
ROM[1264] <= 32'b00000000100000111000001110010011;
ROM[1265] <= 32'b01000000011100010000001110110011;
ROM[1266] <= 32'b00000000011100000000001000110011;
ROM[1267] <= 32'b00000000001000000000000110110011;
ROM[1268] <= 32'b00001110110100010000000011101111;
ROM[1269] <= 32'b11111111110000010000000100010011;
ROM[1270] <= 32'b00000000000000010010001110000011;
ROM[1271] <= 32'b00000000011101100010000000100011;
ROM[1272] <= 32'b00000101110000011010001110000011;
ROM[1273] <= 32'b00000000011100010010000000100011;
ROM[1274] <= 32'b00000000010000010000000100010011;
ROM[1275] <= 32'b00000101000000000000001110010011;
ROM[1276] <= 32'b00000000011100010010000000100011;
ROM[1277] <= 32'b00000000010000010000000100010011;
ROM[1278] <= 32'b00000000000000000001001110110111;
ROM[1279] <= 32'b01000100010000111000001110010011;
ROM[1280] <= 32'b00000000111000111000001110110011;
ROM[1281] <= 32'b00000000011100010010000000100011;
ROM[1282] <= 32'b00000000010000010000000100010011;
ROM[1283] <= 32'b00000000001100010010000000100011;
ROM[1284] <= 32'b00000000010000010000000100010011;
ROM[1285] <= 32'b00000000010000010010000000100011;
ROM[1286] <= 32'b00000000010000010000000100010011;
ROM[1287] <= 32'b00000000010100010010000000100011;
ROM[1288] <= 32'b00000000010000010000000100010011;
ROM[1289] <= 32'b00000000011000010010000000100011;
ROM[1290] <= 32'b00000000010000010000000100010011;
ROM[1291] <= 32'b00000001010000000000001110010011;
ROM[1292] <= 32'b00000000100000111000001110010011;
ROM[1293] <= 32'b01000000011100010000001110110011;
ROM[1294] <= 32'b00000000011100000000001000110011;
ROM[1295] <= 32'b00000000001000000000000110110011;
ROM[1296] <= 32'b00000111110100010000000011101111;
ROM[1297] <= 32'b11111111110000010000000100010011;
ROM[1298] <= 32'b00000000000000010010001110000011;
ROM[1299] <= 32'b00000000011101100010000000100011;
ROM[1300] <= 32'b00000101110000011010001110000011;
ROM[1301] <= 32'b00000000011100010010000000100011;
ROM[1302] <= 32'b00000000010000010000000100010011;
ROM[1303] <= 32'b00000100100100000000001110010011;
ROM[1304] <= 32'b00000000011100010010000000100011;
ROM[1305] <= 32'b00000000010000010000000100010011;
ROM[1306] <= 32'b00000000000000000001001110110111;
ROM[1307] <= 32'b01001011010000111000001110010011;
ROM[1308] <= 32'b00000000111000111000001110110011;
ROM[1309] <= 32'b00000000011100010010000000100011;
ROM[1310] <= 32'b00000000010000010000000100010011;
ROM[1311] <= 32'b00000000001100010010000000100011;
ROM[1312] <= 32'b00000000010000010000000100010011;
ROM[1313] <= 32'b00000000010000010010000000100011;
ROM[1314] <= 32'b00000000010000010000000100010011;
ROM[1315] <= 32'b00000000010100010010000000100011;
ROM[1316] <= 32'b00000000010000010000000100010011;
ROM[1317] <= 32'b00000000011000010010000000100011;
ROM[1318] <= 32'b00000000010000010000000100010011;
ROM[1319] <= 32'b00000001010000000000001110010011;
ROM[1320] <= 32'b00000000100000111000001110010011;
ROM[1321] <= 32'b01000000011100010000001110110011;
ROM[1322] <= 32'b00000000011100000000001000110011;
ROM[1323] <= 32'b00000000001000000000000110110011;
ROM[1324] <= 32'b00000000110100010000000011101111;
ROM[1325] <= 32'b11111111110000010000000100010011;
ROM[1326] <= 32'b00000000000000010010001110000011;
ROM[1327] <= 32'b00000000011101100010000000100011;
ROM[1328] <= 32'b00000101110000011010001110000011;
ROM[1329] <= 32'b00000000011100010010000000100011;
ROM[1330] <= 32'b00000000010000010000000100010011;
ROM[1331] <= 32'b00000100110000000000001110010011;
ROM[1332] <= 32'b00000000011100010010000000100011;
ROM[1333] <= 32'b00000000010000010000000100010011;
ROM[1334] <= 32'b00000000000000000001001110110111;
ROM[1335] <= 32'b01010010010000111000001110010011;
ROM[1336] <= 32'b00000000111000111000001110110011;
ROM[1337] <= 32'b00000000011100010010000000100011;
ROM[1338] <= 32'b00000000010000010000000100010011;
ROM[1339] <= 32'b00000000001100010010000000100011;
ROM[1340] <= 32'b00000000010000010000000100010011;
ROM[1341] <= 32'b00000000010000010010000000100011;
ROM[1342] <= 32'b00000000010000010000000100010011;
ROM[1343] <= 32'b00000000010100010010000000100011;
ROM[1344] <= 32'b00000000010000010000000100010011;
ROM[1345] <= 32'b00000000011000010010000000100011;
ROM[1346] <= 32'b00000000010000010000000100010011;
ROM[1347] <= 32'b00000001010000000000001110010011;
ROM[1348] <= 32'b00000000100000111000001110010011;
ROM[1349] <= 32'b01000000011100010000001110110011;
ROM[1350] <= 32'b00000000011100000000001000110011;
ROM[1351] <= 32'b00000000001000000000000110110011;
ROM[1352] <= 32'b01111001110000010000000011101111;
ROM[1353] <= 32'b11111111110000010000000100010011;
ROM[1354] <= 32'b00000000000000010010001110000011;
ROM[1355] <= 32'b00000000011101100010000000100011;
ROM[1356] <= 32'b00000101110000011010001110000011;
ROM[1357] <= 32'b00000000011100010010000000100011;
ROM[1358] <= 32'b00000000010000010000000100010011;
ROM[1359] <= 32'b00000100010100000000001110010011;
ROM[1360] <= 32'b00000000011100010010000000100011;
ROM[1361] <= 32'b00000000010000010000000100010011;
ROM[1362] <= 32'b00000000000000000001001110110111;
ROM[1363] <= 32'b01011001010000111000001110010011;
ROM[1364] <= 32'b00000000111000111000001110110011;
ROM[1365] <= 32'b00000000011100010010000000100011;
ROM[1366] <= 32'b00000000010000010000000100010011;
ROM[1367] <= 32'b00000000001100010010000000100011;
ROM[1368] <= 32'b00000000010000010000000100010011;
ROM[1369] <= 32'b00000000010000010010000000100011;
ROM[1370] <= 32'b00000000010000010000000100010011;
ROM[1371] <= 32'b00000000010100010010000000100011;
ROM[1372] <= 32'b00000000010000010000000100010011;
ROM[1373] <= 32'b00000000011000010010000000100011;
ROM[1374] <= 32'b00000000010000010000000100010011;
ROM[1375] <= 32'b00000001010000000000001110010011;
ROM[1376] <= 32'b00000000100000111000001110010011;
ROM[1377] <= 32'b01000000011100010000001110110011;
ROM[1378] <= 32'b00000000011100000000001000110011;
ROM[1379] <= 32'b00000000001000000000000110110011;
ROM[1380] <= 32'b01110010110000010000000011101111;
ROM[1381] <= 32'b11111111110000010000000100010011;
ROM[1382] <= 32'b00000000000000010010001110000011;
ROM[1383] <= 32'b00000000011101100010000000100011;
ROM[1384] <= 32'b00000101110000011010001110000011;
ROM[1385] <= 32'b00000000011100010010000000100011;
ROM[1386] <= 32'b00000000010000010000000100010011;
ROM[1387] <= 32'b00000101001000000000001110010011;
ROM[1388] <= 32'b00000000011100010010000000100011;
ROM[1389] <= 32'b00000000010000010000000100010011;
ROM[1390] <= 32'b00000000000000000001001110110111;
ROM[1391] <= 32'b01100000010000111000001110010011;
ROM[1392] <= 32'b00000000111000111000001110110011;
ROM[1393] <= 32'b00000000011100010010000000100011;
ROM[1394] <= 32'b00000000010000010000000100010011;
ROM[1395] <= 32'b00000000001100010010000000100011;
ROM[1396] <= 32'b00000000010000010000000100010011;
ROM[1397] <= 32'b00000000010000010010000000100011;
ROM[1398] <= 32'b00000000010000010000000100010011;
ROM[1399] <= 32'b00000000010100010010000000100011;
ROM[1400] <= 32'b00000000010000010000000100010011;
ROM[1401] <= 32'b00000000011000010010000000100011;
ROM[1402] <= 32'b00000000010000010000000100010011;
ROM[1403] <= 32'b00000001010000000000001110010011;
ROM[1404] <= 32'b00000000100000111000001110010011;
ROM[1405] <= 32'b01000000011100010000001110110011;
ROM[1406] <= 32'b00000000011100000000001000110011;
ROM[1407] <= 32'b00000000001000000000000110110011;
ROM[1408] <= 32'b01101011110000010000000011101111;
ROM[1409] <= 32'b11111111110000010000000100010011;
ROM[1410] <= 32'b00000000000000010010001110000011;
ROM[1411] <= 32'b00000000011101100010000000100011;
ROM[1412] <= 32'b00000101110000011010001110000011;
ROM[1413] <= 32'b00000100011100011010111000100011;
ROM[1414] <= 32'b00000000011100000000001110010011;
ROM[1415] <= 32'b00000000011100010010000000100011;
ROM[1416] <= 32'b00000000010000010000000100010011;
ROM[1417] <= 32'b00000000000000000001001110110111;
ROM[1418] <= 32'b01100111000000111000001110010011;
ROM[1419] <= 32'b00000000111000111000001110110011;
ROM[1420] <= 32'b00000000011100010010000000100011;
ROM[1421] <= 32'b00000000010000010000000100010011;
ROM[1422] <= 32'b00000000001100010010000000100011;
ROM[1423] <= 32'b00000000010000010000000100010011;
ROM[1424] <= 32'b00000000010000010010000000100011;
ROM[1425] <= 32'b00000000010000010000000100010011;
ROM[1426] <= 32'b00000000010100010010000000100011;
ROM[1427] <= 32'b00000000010000010000000100010011;
ROM[1428] <= 32'b00000000011000010010000000100011;
ROM[1429] <= 32'b00000000010000010000000100010011;
ROM[1430] <= 32'b00000001010000000000001110010011;
ROM[1431] <= 32'b00000000010000111000001110010011;
ROM[1432] <= 32'b01000000011100010000001110110011;
ROM[1433] <= 32'b00000000011100000000001000110011;
ROM[1434] <= 32'b00000000001000000000000110110011;
ROM[1435] <= 32'b00101001010000010000000011101111;
ROM[1436] <= 32'b11111111110000010000000100010011;
ROM[1437] <= 32'b00000000000000010010001110000011;
ROM[1438] <= 32'b00000110011100011010000000100011;
ROM[1439] <= 32'b00000110000000011010001110000011;
ROM[1440] <= 32'b00000000011100010010000000100011;
ROM[1441] <= 32'b00000000010000010000000100010011;
ROM[1442] <= 32'b00000101011000000000001110010011;
ROM[1443] <= 32'b00000000011100010010000000100011;
ROM[1444] <= 32'b00000000010000010000000100010011;
ROM[1445] <= 32'b00000000000000000001001110110111;
ROM[1446] <= 32'b01101110000000111000001110010011;
ROM[1447] <= 32'b00000000111000111000001110110011;
ROM[1448] <= 32'b00000000011100010010000000100011;
ROM[1449] <= 32'b00000000010000010000000100010011;
ROM[1450] <= 32'b00000000001100010010000000100011;
ROM[1451] <= 32'b00000000010000010000000100010011;
ROM[1452] <= 32'b00000000010000010010000000100011;
ROM[1453] <= 32'b00000000010000010000000100010011;
ROM[1454] <= 32'b00000000010100010010000000100011;
ROM[1455] <= 32'b00000000010000010000000100010011;
ROM[1456] <= 32'b00000000011000010010000000100011;
ROM[1457] <= 32'b00000000010000010000000100010011;
ROM[1458] <= 32'b00000001010000000000001110010011;
ROM[1459] <= 32'b00000000100000111000001110010011;
ROM[1460] <= 32'b01000000011100010000001110110011;
ROM[1461] <= 32'b00000000011100000000001000110011;
ROM[1462] <= 32'b00000000001000000000000110110011;
ROM[1463] <= 32'b01011110000000010000000011101111;
ROM[1464] <= 32'b11111111110000010000000100010011;
ROM[1465] <= 32'b00000000000000010010001110000011;
ROM[1466] <= 32'b00000000011101100010000000100011;
ROM[1467] <= 32'b00000110000000011010001110000011;
ROM[1468] <= 32'b00000000011100010010000000100011;
ROM[1469] <= 32'b00000000010000010000000100010011;
ROM[1470] <= 32'b00000100100100000000001110010011;
ROM[1471] <= 32'b00000000011100010010000000100011;
ROM[1472] <= 32'b00000000010000010000000100010011;
ROM[1473] <= 32'b00000000000000000001001110110111;
ROM[1474] <= 32'b01110101000000111000001110010011;
ROM[1475] <= 32'b00000000111000111000001110110011;
ROM[1476] <= 32'b00000000011100010010000000100011;
ROM[1477] <= 32'b00000000010000010000000100010011;
ROM[1478] <= 32'b00000000001100010010000000100011;
ROM[1479] <= 32'b00000000010000010000000100010011;
ROM[1480] <= 32'b00000000010000010010000000100011;
ROM[1481] <= 32'b00000000010000010000000100010011;
ROM[1482] <= 32'b00000000010100010010000000100011;
ROM[1483] <= 32'b00000000010000010000000100010011;
ROM[1484] <= 32'b00000000011000010010000000100011;
ROM[1485] <= 32'b00000000010000010000000100010011;
ROM[1486] <= 32'b00000001010000000000001110010011;
ROM[1487] <= 32'b00000000100000111000001110010011;
ROM[1488] <= 32'b01000000011100010000001110110011;
ROM[1489] <= 32'b00000000011100000000001000110011;
ROM[1490] <= 32'b00000000001000000000000110110011;
ROM[1491] <= 32'b01010111000000010000000011101111;
ROM[1492] <= 32'b11111111110000010000000100010011;
ROM[1493] <= 32'b00000000000000010010001110000011;
ROM[1494] <= 32'b00000000011101100010000000100011;
ROM[1495] <= 32'b00000110000000011010001110000011;
ROM[1496] <= 32'b00000000011100010010000000100011;
ROM[1497] <= 32'b00000000010000010000000100010011;
ROM[1498] <= 32'b00000101001000000000001110010011;
ROM[1499] <= 32'b00000000011100010010000000100011;
ROM[1500] <= 32'b00000000010000010000000100010011;
ROM[1501] <= 32'b00000000000000000001001110110111;
ROM[1502] <= 32'b01111100000000111000001110010011;
ROM[1503] <= 32'b00000000111000111000001110110011;
ROM[1504] <= 32'b00000000011100010010000000100011;
ROM[1505] <= 32'b00000000010000010000000100010011;
ROM[1506] <= 32'b00000000001100010010000000100011;
ROM[1507] <= 32'b00000000010000010000000100010011;
ROM[1508] <= 32'b00000000010000010010000000100011;
ROM[1509] <= 32'b00000000010000010000000100010011;
ROM[1510] <= 32'b00000000010100010010000000100011;
ROM[1511] <= 32'b00000000010000010000000100010011;
ROM[1512] <= 32'b00000000011000010010000000100011;
ROM[1513] <= 32'b00000000010000010000000100010011;
ROM[1514] <= 32'b00000001010000000000001110010011;
ROM[1515] <= 32'b00000000100000111000001110010011;
ROM[1516] <= 32'b01000000011100010000001110110011;
ROM[1517] <= 32'b00000000011100000000001000110011;
ROM[1518] <= 32'b00000000001000000000000110110011;
ROM[1519] <= 32'b01010000000000010000000011101111;
ROM[1520] <= 32'b11111111110000010000000100010011;
ROM[1521] <= 32'b00000000000000010010001110000011;
ROM[1522] <= 32'b00000000011101100010000000100011;
ROM[1523] <= 32'b00000110000000011010001110000011;
ROM[1524] <= 32'b00000000011100010010000000100011;
ROM[1525] <= 32'b00000000010000010000000100010011;
ROM[1526] <= 32'b00000101010000000000001110010011;
ROM[1527] <= 32'b00000000011100010010000000100011;
ROM[1528] <= 32'b00000000010000010000000100010011;
ROM[1529] <= 32'b00000000000000000010001110110111;
ROM[1530] <= 32'b10000011000000111000001110010011;
ROM[1531] <= 32'b00000000111000111000001110110011;
ROM[1532] <= 32'b00000000011100010010000000100011;
ROM[1533] <= 32'b00000000010000010000000100010011;
ROM[1534] <= 32'b00000000001100010010000000100011;
ROM[1535] <= 32'b00000000010000010000000100010011;
ROM[1536] <= 32'b00000000010000010010000000100011;
ROM[1537] <= 32'b00000000010000010000000100010011;
ROM[1538] <= 32'b00000000010100010010000000100011;
ROM[1539] <= 32'b00000000010000010000000100010011;
ROM[1540] <= 32'b00000000011000010010000000100011;
ROM[1541] <= 32'b00000000010000010000000100010011;
ROM[1542] <= 32'b00000001010000000000001110010011;
ROM[1543] <= 32'b00000000100000111000001110010011;
ROM[1544] <= 32'b01000000011100010000001110110011;
ROM[1545] <= 32'b00000000011100000000001000110011;
ROM[1546] <= 32'b00000000001000000000000110110011;
ROM[1547] <= 32'b01001001000000010000000011101111;
ROM[1548] <= 32'b11111111110000010000000100010011;
ROM[1549] <= 32'b00000000000000010010001110000011;
ROM[1550] <= 32'b00000000011101100010000000100011;
ROM[1551] <= 32'b00000110000000011010001110000011;
ROM[1552] <= 32'b00000000011100010010000000100011;
ROM[1553] <= 32'b00000000010000010000000100010011;
ROM[1554] <= 32'b00000101010100000000001110010011;
ROM[1555] <= 32'b00000000011100010010000000100011;
ROM[1556] <= 32'b00000000010000010000000100010011;
ROM[1557] <= 32'b00000000000000000010001110110111;
ROM[1558] <= 32'b10001010000000111000001110010011;
ROM[1559] <= 32'b00000000111000111000001110110011;
ROM[1560] <= 32'b00000000011100010010000000100011;
ROM[1561] <= 32'b00000000010000010000000100010011;
ROM[1562] <= 32'b00000000001100010010000000100011;
ROM[1563] <= 32'b00000000010000010000000100010011;
ROM[1564] <= 32'b00000000010000010010000000100011;
ROM[1565] <= 32'b00000000010000010000000100010011;
ROM[1566] <= 32'b00000000010100010010000000100011;
ROM[1567] <= 32'b00000000010000010000000100010011;
ROM[1568] <= 32'b00000000011000010010000000100011;
ROM[1569] <= 32'b00000000010000010000000100010011;
ROM[1570] <= 32'b00000001010000000000001110010011;
ROM[1571] <= 32'b00000000100000111000001110010011;
ROM[1572] <= 32'b01000000011100010000001110110011;
ROM[1573] <= 32'b00000000011100000000001000110011;
ROM[1574] <= 32'b00000000001000000000000110110011;
ROM[1575] <= 32'b01000010000000010000000011101111;
ROM[1576] <= 32'b11111111110000010000000100010011;
ROM[1577] <= 32'b00000000000000010010001110000011;
ROM[1578] <= 32'b00000000011101100010000000100011;
ROM[1579] <= 32'b00000110000000011010001110000011;
ROM[1580] <= 32'b00000000011100010010000000100011;
ROM[1581] <= 32'b00000000010000010000000100010011;
ROM[1582] <= 32'b00000100000100000000001110010011;
ROM[1583] <= 32'b00000000011100010010000000100011;
ROM[1584] <= 32'b00000000010000010000000100010011;
ROM[1585] <= 32'b00000000000000000010001110110111;
ROM[1586] <= 32'b10010001000000111000001110010011;
ROM[1587] <= 32'b00000000111000111000001110110011;
ROM[1588] <= 32'b00000000011100010010000000100011;
ROM[1589] <= 32'b00000000010000010000000100010011;
ROM[1590] <= 32'b00000000001100010010000000100011;
ROM[1591] <= 32'b00000000010000010000000100010011;
ROM[1592] <= 32'b00000000010000010010000000100011;
ROM[1593] <= 32'b00000000010000010000000100010011;
ROM[1594] <= 32'b00000000010100010010000000100011;
ROM[1595] <= 32'b00000000010000010000000100010011;
ROM[1596] <= 32'b00000000011000010010000000100011;
ROM[1597] <= 32'b00000000010000010000000100010011;
ROM[1598] <= 32'b00000001010000000000001110010011;
ROM[1599] <= 32'b00000000100000111000001110010011;
ROM[1600] <= 32'b01000000011100010000001110110011;
ROM[1601] <= 32'b00000000011100000000001000110011;
ROM[1602] <= 32'b00000000001000000000000110110011;
ROM[1603] <= 32'b00111011000000010000000011101111;
ROM[1604] <= 32'b11111111110000010000000100010011;
ROM[1605] <= 32'b00000000000000010010001110000011;
ROM[1606] <= 32'b00000000011101100010000000100011;
ROM[1607] <= 32'b00000110000000011010001110000011;
ROM[1608] <= 32'b00000000011100010010000000100011;
ROM[1609] <= 32'b00000000010000010000000100010011;
ROM[1610] <= 32'b00000100110000000000001110010011;
ROM[1611] <= 32'b00000000011100010010000000100011;
ROM[1612] <= 32'b00000000010000010000000100010011;
ROM[1613] <= 32'b00000000000000000010001110110111;
ROM[1614] <= 32'b10011000000000111000001110010011;
ROM[1615] <= 32'b00000000111000111000001110110011;
ROM[1616] <= 32'b00000000011100010010000000100011;
ROM[1617] <= 32'b00000000010000010000000100010011;
ROM[1618] <= 32'b00000000001100010010000000100011;
ROM[1619] <= 32'b00000000010000010000000100010011;
ROM[1620] <= 32'b00000000010000010010000000100011;
ROM[1621] <= 32'b00000000010000010000000100010011;
ROM[1622] <= 32'b00000000010100010010000000100011;
ROM[1623] <= 32'b00000000010000010000000100010011;
ROM[1624] <= 32'b00000000011000010010000000100011;
ROM[1625] <= 32'b00000000010000010000000100010011;
ROM[1626] <= 32'b00000001010000000000001110010011;
ROM[1627] <= 32'b00000000100000111000001110010011;
ROM[1628] <= 32'b01000000011100010000001110110011;
ROM[1629] <= 32'b00000000011100000000001000110011;
ROM[1630] <= 32'b00000000001000000000000110110011;
ROM[1631] <= 32'b00110100000000010000000011101111;
ROM[1632] <= 32'b11111111110000010000000100010011;
ROM[1633] <= 32'b00000000000000010010001110000011;
ROM[1634] <= 32'b00000000011101100010000000100011;
ROM[1635] <= 32'b00000110000000011010001110000011;
ROM[1636] <= 32'b00000110011100011010000000100011;
ROM[1637] <= 32'b00000000000000000000001110010011;
ROM[1638] <= 32'b00000000011100010010000000100011;
ROM[1639] <= 32'b00000000010000010000000100010011;
ROM[1640] <= 32'b00000000000000011010001110000011;
ROM[1641] <= 32'b11111111110000010000000100010011;
ROM[1642] <= 32'b00000000000000010010010000000011;
ROM[1643] <= 32'b00000000011101000000001110110011;
ROM[1644] <= 32'b00000000011100010010000000100011;
ROM[1645] <= 32'b00000000010000010000000100010011;
ROM[1646] <= 32'b00000101000000011010001110000011;
ROM[1647] <= 32'b00000000011101100010000000100011;
ROM[1648] <= 32'b11111111110000010000000100010011;
ROM[1649] <= 32'b00000000000000010010001110000011;
ROM[1650] <= 32'b00000000000000111000001100010011;
ROM[1651] <= 32'b00000000000001100010001110000011;
ROM[1652] <= 32'b00000000110100110000010000110011;
ROM[1653] <= 32'b00000000011101000010000000100011;
ROM[1654] <= 32'b00000000010000000000001110010011;
ROM[1655] <= 32'b00000000011100010010000000100011;
ROM[1656] <= 32'b00000000010000010000000100010011;
ROM[1657] <= 32'b00000000000000011010001110000011;
ROM[1658] <= 32'b11111111110000010000000100010011;
ROM[1659] <= 32'b00000000000000010010010000000011;
ROM[1660] <= 32'b00000000011101000000001110110011;
ROM[1661] <= 32'b00000000011100010010000000100011;
ROM[1662] <= 32'b00000000010000010000000100010011;
ROM[1663] <= 32'b00000101010000011010001110000011;
ROM[1664] <= 32'b00000000011101100010000000100011;
ROM[1665] <= 32'b11111111110000010000000100010011;
ROM[1666] <= 32'b00000000000000010010001110000011;
ROM[1667] <= 32'b00000000000000111000001100010011;
ROM[1668] <= 32'b00000000000001100010001110000011;
ROM[1669] <= 32'b00000000110100110000010000110011;
ROM[1670] <= 32'b00000000011101000010000000100011;
ROM[1671] <= 32'b00000000100000000000001110010011;
ROM[1672] <= 32'b00000000011100010010000000100011;
ROM[1673] <= 32'b00000000010000010000000100010011;
ROM[1674] <= 32'b00000000000000011010001110000011;
ROM[1675] <= 32'b11111111110000010000000100010011;
ROM[1676] <= 32'b00000000000000010010010000000011;
ROM[1677] <= 32'b00000000011101000000001110110011;
ROM[1678] <= 32'b00000000011100010010000000100011;
ROM[1679] <= 32'b00000000010000010000000100010011;
ROM[1680] <= 32'b00000101100000011010001110000011;
ROM[1681] <= 32'b00000000011101100010000000100011;
ROM[1682] <= 32'b11111111110000010000000100010011;
ROM[1683] <= 32'b00000000000000010010001110000011;
ROM[1684] <= 32'b00000000000000111000001100010011;
ROM[1685] <= 32'b00000000000001100010001110000011;
ROM[1686] <= 32'b00000000110100110000010000110011;
ROM[1687] <= 32'b00000000011101000010000000100011;
ROM[1688] <= 32'b00000000110000000000001110010011;
ROM[1689] <= 32'b00000000011100010010000000100011;
ROM[1690] <= 32'b00000000010000010000000100010011;
ROM[1691] <= 32'b00000000000000011010001110000011;
ROM[1692] <= 32'b11111111110000010000000100010011;
ROM[1693] <= 32'b00000000000000010010010000000011;
ROM[1694] <= 32'b00000000011101000000001110110011;
ROM[1695] <= 32'b00000000011100010010000000100011;
ROM[1696] <= 32'b00000000010000010000000100010011;
ROM[1697] <= 32'b00000101110000011010001110000011;
ROM[1698] <= 32'b00000000011101100010000000100011;
ROM[1699] <= 32'b11111111110000010000000100010011;
ROM[1700] <= 32'b00000000000000010010001110000011;
ROM[1701] <= 32'b00000000000000111000001100010011;
ROM[1702] <= 32'b00000000000001100010001110000011;
ROM[1703] <= 32'b00000000110100110000010000110011;
ROM[1704] <= 32'b00000000011101000010000000100011;
ROM[1705] <= 32'b00000001000000000000001110010011;
ROM[1706] <= 32'b00000000011100010010000000100011;
ROM[1707] <= 32'b00000000010000010000000100010011;
ROM[1708] <= 32'b00000000000000011010001110000011;
ROM[1709] <= 32'b11111111110000010000000100010011;
ROM[1710] <= 32'b00000000000000010010010000000011;
ROM[1711] <= 32'b00000000011101000000001110110011;
ROM[1712] <= 32'b00000000011100010010000000100011;
ROM[1713] <= 32'b00000000010000010000000100010011;
ROM[1714] <= 32'b00000110000000011010001110000011;
ROM[1715] <= 32'b00000000011101100010000000100011;
ROM[1716] <= 32'b11111111110000010000000100010011;
ROM[1717] <= 32'b00000000000000010010001110000011;
ROM[1718] <= 32'b00000000000000111000001100010011;
ROM[1719] <= 32'b00000000000001100010001110000011;
ROM[1720] <= 32'b00000000110100110000010000110011;
ROM[1721] <= 32'b00000000011101000010000000100011;
ROM[1722] <= 32'b00000000010100000000001110010011;
ROM[1723] <= 32'b00000000011100010010000000100011;
ROM[1724] <= 32'b00000000010000010000000100010011;
ROM[1725] <= 32'b00000000000000000010001110110111;
ROM[1726] <= 32'b10110100000000111000001110010011;
ROM[1727] <= 32'b00000000111000111000001110110011;
ROM[1728] <= 32'b00000000011100010010000000100011;
ROM[1729] <= 32'b00000000010000010000000100010011;
ROM[1730] <= 32'b00000000001100010010000000100011;
ROM[1731] <= 32'b00000000010000010000000100010011;
ROM[1732] <= 32'b00000000010000010010000000100011;
ROM[1733] <= 32'b00000000010000010000000100010011;
ROM[1734] <= 32'b00000000010100010010000000100011;
ROM[1735] <= 32'b00000000010000010000000100010011;
ROM[1736] <= 32'b00000000011000010010000000100011;
ROM[1737] <= 32'b00000000010000010000000100010011;
ROM[1738] <= 32'b00000001010000000000001110010011;
ROM[1739] <= 32'b00000000010000111000001110010011;
ROM[1740] <= 32'b01000000011100010000001110110011;
ROM[1741] <= 32'b00000000011100000000001000110011;
ROM[1742] <= 32'b00000000001000000000000110110011;
ROM[1743] <= 32'b10010000010111111110000011101111;
ROM[1744] <= 32'b11111111110000010000000100010011;
ROM[1745] <= 32'b00000000000000010010001110000011;
ROM[1746] <= 32'b00000100011100011010000000100011;
ROM[1747] <= 32'b00000000000000000000001110010011;
ROM[1748] <= 32'b00000000011100010010000000100011;
ROM[1749] <= 32'b00000000010000010000000100010011;
ROM[1750] <= 32'b00000100000000011010001110000011;
ROM[1751] <= 32'b11111111110000010000000100010011;
ROM[1752] <= 32'b00000000000000010010010000000011;
ROM[1753] <= 32'b00000000011101000000001110110011;
ROM[1754] <= 32'b00000000011100010010000000100011;
ROM[1755] <= 32'b00000000010000010000000100010011;
ROM[1756] <= 32'b00000000010000000000001110010011;
ROM[1757] <= 32'b00000000011101100010000000100011;
ROM[1758] <= 32'b11111111110000010000000100010011;
ROM[1759] <= 32'b00000000000000010010001110000011;
ROM[1760] <= 32'b00000000000000111000001100010011;
ROM[1761] <= 32'b00000000000001100010001110000011;
ROM[1762] <= 32'b00000000110100110000010000110011;
ROM[1763] <= 32'b00000000011101000010000000100011;
ROM[1764] <= 32'b00000000010000000000001110010011;
ROM[1765] <= 32'b00000000011100010010000000100011;
ROM[1766] <= 32'b00000000010000010000000100010011;
ROM[1767] <= 32'b00000100000000011010001110000011;
ROM[1768] <= 32'b11111111110000010000000100010011;
ROM[1769] <= 32'b00000000000000010010010000000011;
ROM[1770] <= 32'b00000000011101000000001110110011;
ROM[1771] <= 32'b00000000011100010010000000100011;
ROM[1772] <= 32'b00000000010000010000000100010011;
ROM[1773] <= 32'b00000000101100000000001110010011;
ROM[1774] <= 32'b00000000011101100010000000100011;
ROM[1775] <= 32'b11111111110000010000000100010011;
ROM[1776] <= 32'b00000000000000010010001110000011;
ROM[1777] <= 32'b00000000000000111000001100010011;
ROM[1778] <= 32'b00000000000001100010001110000011;
ROM[1779] <= 32'b00000000110100110000010000110011;
ROM[1780] <= 32'b00000000011101000010000000100011;
ROM[1781] <= 32'b00000000100000000000001110010011;
ROM[1782] <= 32'b00000000011100010010000000100011;
ROM[1783] <= 32'b00000000010000010000000100010011;
ROM[1784] <= 32'b00000100000000011010001110000011;
ROM[1785] <= 32'b11111111110000010000000100010011;
ROM[1786] <= 32'b00000000000000010010010000000011;
ROM[1787] <= 32'b00000000011101000000001110110011;
ROM[1788] <= 32'b00000000011100010010000000100011;
ROM[1789] <= 32'b00000000010000010000000100010011;
ROM[1790] <= 32'b00000000100000000000001110010011;
ROM[1791] <= 32'b00000000011101100010000000100011;
ROM[1792] <= 32'b11111111110000010000000100010011;
ROM[1793] <= 32'b00000000000000010010001110000011;
ROM[1794] <= 32'b00000000000000111000001100010011;
ROM[1795] <= 32'b00000000000001100010001110000011;
ROM[1796] <= 32'b00000000110100110000010000110011;
ROM[1797] <= 32'b00000000011101000010000000100011;
ROM[1798] <= 32'b00000000110000000000001110010011;
ROM[1799] <= 32'b00000000011100010010000000100011;
ROM[1800] <= 32'b00000000010000010000000100010011;
ROM[1801] <= 32'b00000100000000011010001110000011;
ROM[1802] <= 32'b11111111110000010000000100010011;
ROM[1803] <= 32'b00000000000000010010010000000011;
ROM[1804] <= 32'b00000000011101000000001110110011;
ROM[1805] <= 32'b00000000011100010010000000100011;
ROM[1806] <= 32'b00000000010000010000000100010011;
ROM[1807] <= 32'b00000000100000000000001110010011;
ROM[1808] <= 32'b00000000011101100010000000100011;
ROM[1809] <= 32'b11111111110000010000000100010011;
ROM[1810] <= 32'b00000000000000010010001110000011;
ROM[1811] <= 32'b00000000000000111000001100010011;
ROM[1812] <= 32'b00000000000001100010001110000011;
ROM[1813] <= 32'b00000000110100110000010000110011;
ROM[1814] <= 32'b00000000011101000010000000100011;
ROM[1815] <= 32'b00000001000000000000001110010011;
ROM[1816] <= 32'b00000000011100010010000000100011;
ROM[1817] <= 32'b00000000010000010000000100010011;
ROM[1818] <= 32'b00000100000000011010001110000011;
ROM[1819] <= 32'b11111111110000010000000100010011;
ROM[1820] <= 32'b00000000000000010010010000000011;
ROM[1821] <= 32'b00000000011101000000001110110011;
ROM[1822] <= 32'b00000000011100010010000000100011;
ROM[1823] <= 32'b00000000010000010000000100010011;
ROM[1824] <= 32'b00000000011100000000001110010011;
ROM[1825] <= 32'b00000000011101100010000000100011;
ROM[1826] <= 32'b11111111110000010000000100010011;
ROM[1827] <= 32'b00000000000000010010001110000011;
ROM[1828] <= 32'b00000000000000111000001100010011;
ROM[1829] <= 32'b00000000000001100010001110000011;
ROM[1830] <= 32'b00000000110100110000010000110011;
ROM[1831] <= 32'b00000000011101000010000000100011;
ROM[1832] <= 32'b00000000000000000000001110010011;
ROM[1833] <= 32'b00000000011100011010010000100011;
ROM[1834] <= 32'b00000101111100000000001110010011;
ROM[1835] <= 32'b00000010011100011010100000100011;
ROM[1836] <= 32'b00000000011000000000001110010011;
ROM[1837] <= 32'b00000000011100010010000000100011;
ROM[1838] <= 32'b00000000010000010000000100010011;
ROM[1839] <= 32'b00000000000000000010001110110111;
ROM[1840] <= 32'b11010000100000111000001110010011;
ROM[1841] <= 32'b00000000111000111000001110110011;
ROM[1842] <= 32'b00000000011100010010000000100011;
ROM[1843] <= 32'b00000000010000010000000100010011;
ROM[1844] <= 32'b00000000001100010010000000100011;
ROM[1845] <= 32'b00000000010000010000000100010011;
ROM[1846] <= 32'b00000000010000010010000000100011;
ROM[1847] <= 32'b00000000010000010000000100010011;
ROM[1848] <= 32'b00000000010100010010000000100011;
ROM[1849] <= 32'b00000000010000010000000100010011;
ROM[1850] <= 32'b00000000011000010010000000100011;
ROM[1851] <= 32'b00000000010000010000000100010011;
ROM[1852] <= 32'b00000001010000000000001110010011;
ROM[1853] <= 32'b00000000010000111000001110010011;
ROM[1854] <= 32'b01000000011100010000001110110011;
ROM[1855] <= 32'b00000000011100000000001000110011;
ROM[1856] <= 32'b00000000001000000000000110110011;
ROM[1857] <= 32'b00111111110100001111000011101111;
ROM[1858] <= 32'b11111111110000010000000100010011;
ROM[1859] <= 32'b00000000000000010010001110000011;
ROM[1860] <= 32'b00000110011100011010001000100011;
ROM[1861] <= 32'b00000110010000011010001110000011;
ROM[1862] <= 32'b00000000011100010010000000100011;
ROM[1863] <= 32'b00000000010000010000000100010011;
ROM[1864] <= 32'b00000111011100000000001110010011;
ROM[1865] <= 32'b00000000011100010010000000100011;
ROM[1866] <= 32'b00000000010000010000000100010011;
ROM[1867] <= 32'b00000000000000000010001110110111;
ROM[1868] <= 32'b11010111100000111000001110010011;
ROM[1869] <= 32'b00000000111000111000001110110011;
ROM[1870] <= 32'b00000000011100010010000000100011;
ROM[1871] <= 32'b00000000010000010000000100010011;
ROM[1872] <= 32'b00000000001100010010000000100011;
ROM[1873] <= 32'b00000000010000010000000100010011;
ROM[1874] <= 32'b00000000010000010010000000100011;
ROM[1875] <= 32'b00000000010000010000000100010011;
ROM[1876] <= 32'b00000000010100010010000000100011;
ROM[1877] <= 32'b00000000010000010000000100010011;
ROM[1878] <= 32'b00000000011000010010000000100011;
ROM[1879] <= 32'b00000000010000010000000100010011;
ROM[1880] <= 32'b00000001010000000000001110010011;
ROM[1881] <= 32'b00000000100000111000001110010011;
ROM[1882] <= 32'b01000000011100010000001110110011;
ROM[1883] <= 32'b00000000011100000000001000110011;
ROM[1884] <= 32'b00000000001000000000000110110011;
ROM[1885] <= 32'b01110100100100001111000011101111;
ROM[1886] <= 32'b11111111110000010000000100010011;
ROM[1887] <= 32'b00000000000000010010001110000011;
ROM[1888] <= 32'b00000000011101100010000000100011;
ROM[1889] <= 32'b00000110010000011010001110000011;
ROM[1890] <= 32'b00000000011100010010000000100011;
ROM[1891] <= 32'b00000000010000010000000100010011;
ROM[1892] <= 32'b00000110111100000000001110010011;
ROM[1893] <= 32'b00000000011100010010000000100011;
ROM[1894] <= 32'b00000000010000010000000100010011;
ROM[1895] <= 32'b00000000000000000010001110110111;
ROM[1896] <= 32'b11011110100000111000001110010011;
ROM[1897] <= 32'b00000000111000111000001110110011;
ROM[1898] <= 32'b00000000011100010010000000100011;
ROM[1899] <= 32'b00000000010000010000000100010011;
ROM[1900] <= 32'b00000000001100010010000000100011;
ROM[1901] <= 32'b00000000010000010000000100010011;
ROM[1902] <= 32'b00000000010000010010000000100011;
ROM[1903] <= 32'b00000000010000010000000100010011;
ROM[1904] <= 32'b00000000010100010010000000100011;
ROM[1905] <= 32'b00000000010000010000000100010011;
ROM[1906] <= 32'b00000000011000010010000000100011;
ROM[1907] <= 32'b00000000010000010000000100010011;
ROM[1908] <= 32'b00000001010000000000001110010011;
ROM[1909] <= 32'b00000000100000111000001110010011;
ROM[1910] <= 32'b01000000011100010000001110110011;
ROM[1911] <= 32'b00000000011100000000001000110011;
ROM[1912] <= 32'b00000000001000000000000110110011;
ROM[1913] <= 32'b01101101100100001111000011101111;
ROM[1914] <= 32'b11111111110000010000000100010011;
ROM[1915] <= 32'b00000000000000010010001110000011;
ROM[1916] <= 32'b00000000011101100010000000100011;
ROM[1917] <= 32'b00000110010000011010001110000011;
ROM[1918] <= 32'b00000000011100010010000000100011;
ROM[1919] <= 32'b00000000010000010000000100010011;
ROM[1920] <= 32'b00000111001000000000001110010011;
ROM[1921] <= 32'b00000000011100010010000000100011;
ROM[1922] <= 32'b00000000010000010000000100010011;
ROM[1923] <= 32'b00000000000000000010001110110111;
ROM[1924] <= 32'b11100101100000111000001110010011;
ROM[1925] <= 32'b00000000111000111000001110110011;
ROM[1926] <= 32'b00000000011100010010000000100011;
ROM[1927] <= 32'b00000000010000010000000100010011;
ROM[1928] <= 32'b00000000001100010010000000100011;
ROM[1929] <= 32'b00000000010000010000000100010011;
ROM[1930] <= 32'b00000000010000010010000000100011;
ROM[1931] <= 32'b00000000010000010000000100010011;
ROM[1932] <= 32'b00000000010100010010000000100011;
ROM[1933] <= 32'b00000000010000010000000100010011;
ROM[1934] <= 32'b00000000011000010010000000100011;
ROM[1935] <= 32'b00000000010000010000000100010011;
ROM[1936] <= 32'b00000001010000000000001110010011;
ROM[1937] <= 32'b00000000100000111000001110010011;
ROM[1938] <= 32'b01000000011100010000001110110011;
ROM[1939] <= 32'b00000000011100000000001000110011;
ROM[1940] <= 32'b00000000001000000000000110110011;
ROM[1941] <= 32'b01100110100100001111000011101111;
ROM[1942] <= 32'b11111111110000010000000100010011;
ROM[1943] <= 32'b00000000000000010010001110000011;
ROM[1944] <= 32'b00000000011101100010000000100011;
ROM[1945] <= 32'b00000110010000011010001110000011;
ROM[1946] <= 32'b00000000011100010010000000100011;
ROM[1947] <= 32'b00000000010000010000000100010011;
ROM[1948] <= 32'b00000110010000000000001110010011;
ROM[1949] <= 32'b00000000011100010010000000100011;
ROM[1950] <= 32'b00000000010000010000000100010011;
ROM[1951] <= 32'b00000000000000000010001110110111;
ROM[1952] <= 32'b11101100100000111000001110010011;
ROM[1953] <= 32'b00000000111000111000001110110011;
ROM[1954] <= 32'b00000000011100010010000000100011;
ROM[1955] <= 32'b00000000010000010000000100010011;
ROM[1956] <= 32'b00000000001100010010000000100011;
ROM[1957] <= 32'b00000000010000010000000100010011;
ROM[1958] <= 32'b00000000010000010010000000100011;
ROM[1959] <= 32'b00000000010000010000000100010011;
ROM[1960] <= 32'b00000000010100010010000000100011;
ROM[1961] <= 32'b00000000010000010000000100010011;
ROM[1962] <= 32'b00000000011000010010000000100011;
ROM[1963] <= 32'b00000000010000010000000100010011;
ROM[1964] <= 32'b00000001010000000000001110010011;
ROM[1965] <= 32'b00000000100000111000001110010011;
ROM[1966] <= 32'b01000000011100010000001110110011;
ROM[1967] <= 32'b00000000011100000000001000110011;
ROM[1968] <= 32'b00000000001000000000000110110011;
ROM[1969] <= 32'b01011111100100001111000011101111;
ROM[1970] <= 32'b11111111110000010000000100010011;
ROM[1971] <= 32'b00000000000000010010001110000011;
ROM[1972] <= 32'b00000000011101100010000000100011;
ROM[1973] <= 32'b00000110010000011010001110000011;
ROM[1974] <= 32'b00000000011100010010000000100011;
ROM[1975] <= 32'b00000000010000010000000100010011;
ROM[1976] <= 32'b00000011101000000000001110010011;
ROM[1977] <= 32'b00000000011100010010000000100011;
ROM[1978] <= 32'b00000000010000010000000100010011;
ROM[1979] <= 32'b00000000000000000010001110110111;
ROM[1980] <= 32'b11110011100000111000001110010011;
ROM[1981] <= 32'b00000000111000111000001110110011;
ROM[1982] <= 32'b00000000011100010010000000100011;
ROM[1983] <= 32'b00000000010000010000000100010011;
ROM[1984] <= 32'b00000000001100010010000000100011;
ROM[1985] <= 32'b00000000010000010000000100010011;
ROM[1986] <= 32'b00000000010000010010000000100011;
ROM[1987] <= 32'b00000000010000010000000100010011;
ROM[1988] <= 32'b00000000010100010010000000100011;
ROM[1989] <= 32'b00000000010000010000000100010011;
ROM[1990] <= 32'b00000000011000010010000000100011;
ROM[1991] <= 32'b00000000010000010000000100010011;
ROM[1992] <= 32'b00000001010000000000001110010011;
ROM[1993] <= 32'b00000000100000111000001110010011;
ROM[1994] <= 32'b01000000011100010000001110110011;
ROM[1995] <= 32'b00000000011100000000001000110011;
ROM[1996] <= 32'b00000000001000000000000110110011;
ROM[1997] <= 32'b01011000100100001111000011101111;
ROM[1998] <= 32'b11111111110000010000000100010011;
ROM[1999] <= 32'b00000000000000010010001110000011;
ROM[2000] <= 32'b00000000011101100010000000100011;
ROM[2001] <= 32'b00000110010000011010001110000011;
ROM[2002] <= 32'b00000000011100010010000000100011;
ROM[2003] <= 32'b00000000010000010000000100010011;
ROM[2004] <= 32'b00000010000000000000001110010011;
ROM[2005] <= 32'b00000000011100010010000000100011;
ROM[2006] <= 32'b00000000010000010000000100010011;
ROM[2007] <= 32'b00000000000000000010001110110111;
ROM[2008] <= 32'b11111010100000111000001110010011;
ROM[2009] <= 32'b00000000111000111000001110110011;
ROM[2010] <= 32'b00000000011100010010000000100011;
ROM[2011] <= 32'b00000000010000010000000100010011;
ROM[2012] <= 32'b00000000001100010010000000100011;
ROM[2013] <= 32'b00000000010000010000000100010011;
ROM[2014] <= 32'b00000000010000010010000000100011;
ROM[2015] <= 32'b00000000010000010000000100010011;
ROM[2016] <= 32'b00000000010100010010000000100011;
ROM[2017] <= 32'b00000000010000010000000100010011;
ROM[2018] <= 32'b00000000011000010010000000100011;
ROM[2019] <= 32'b00000000010000010000000100010011;
ROM[2020] <= 32'b00000001010000000000001110010011;
ROM[2021] <= 32'b00000000100000111000001110010011;
ROM[2022] <= 32'b01000000011100010000001110110011;
ROM[2023] <= 32'b00000000011100000000001000110011;
ROM[2024] <= 32'b00000000001000000000000110110011;
ROM[2025] <= 32'b01010001100100001111000011101111;
ROM[2026] <= 32'b11111111110000010000000100010011;
ROM[2027] <= 32'b00000000000000010010001110000011;
ROM[2028] <= 32'b00000000011101100010000000100011;
ROM[2029] <= 32'b00000110010000011010001110000011;
ROM[2030] <= 32'b00000110011100011010001000100011;
ROM[2031] <= 32'b00000000011100000000001110010011;
ROM[2032] <= 32'b00000000011100010010000000100011;
ROM[2033] <= 32'b00000000010000010000000100010011;
ROM[2034] <= 32'b00000000000000000010001110110111;
ROM[2035] <= 32'b00000001010000111000001110010011;
ROM[2036] <= 32'b00000000111000111000001110110011;
ROM[2037] <= 32'b00000000011100010010000000100011;
ROM[2038] <= 32'b00000000010000010000000100010011;
ROM[2039] <= 32'b00000000001100010010000000100011;
ROM[2040] <= 32'b00000000010000010000000100010011;
ROM[2041] <= 32'b00000000010000010010000000100011;
ROM[2042] <= 32'b00000000010000010000000100010011;
ROM[2043] <= 32'b00000000010100010010000000100011;
ROM[2044] <= 32'b00000000010000010000000100010011;
ROM[2045] <= 32'b00000000011000010010000000100011;
ROM[2046] <= 32'b00000000010000010000000100010011;
ROM[2047] <= 32'b00000001010000000000001110010011;
ROM[2048] <= 32'b00000000010000111000001110010011;
ROM[2049] <= 32'b01000000011100010000001110110011;
ROM[2050] <= 32'b00000000011100000000001000110011;
ROM[2051] <= 32'b00000000001000000000000110110011;
ROM[2052] <= 32'b00001111000100001111000011101111;
ROM[2053] <= 32'b11111111110000010000000100010011;
ROM[2054] <= 32'b00000000000000010010001110000011;
ROM[2055] <= 32'b00000110011100011010010000100011;
ROM[2056] <= 32'b00000110100000011010001110000011;
ROM[2057] <= 32'b00000000011100010010000000100011;
ROM[2058] <= 32'b00000000010000010000000100010011;
ROM[2059] <= 32'b00000100010100000000001110010011;
ROM[2060] <= 32'b00000000011100010010000000100011;
ROM[2061] <= 32'b00000000010000010000000100010011;
ROM[2062] <= 32'b00000000000000000010001110110111;
ROM[2063] <= 32'b00001000010000111000001110010011;
ROM[2064] <= 32'b00000000111000111000001110110011;
ROM[2065] <= 32'b00000000011100010010000000100011;
ROM[2066] <= 32'b00000000010000010000000100010011;
ROM[2067] <= 32'b00000000001100010010000000100011;
ROM[2068] <= 32'b00000000010000010000000100010011;
ROM[2069] <= 32'b00000000010000010010000000100011;
ROM[2070] <= 32'b00000000010000010000000100010011;
ROM[2071] <= 32'b00000000010100010010000000100011;
ROM[2072] <= 32'b00000000010000010000000100010011;
ROM[2073] <= 32'b00000000011000010010000000100011;
ROM[2074] <= 32'b00000000010000010000000100010011;
ROM[2075] <= 32'b00000001010000000000001110010011;
ROM[2076] <= 32'b00000000100000111000001110010011;
ROM[2077] <= 32'b01000000011100010000001110110011;
ROM[2078] <= 32'b00000000011100000000001000110011;
ROM[2079] <= 32'b00000000001000000000000110110011;
ROM[2080] <= 32'b01000011110100001111000011101111;
ROM[2081] <= 32'b11111111110000010000000100010011;
ROM[2082] <= 32'b00000000000000010010001110000011;
ROM[2083] <= 32'b00000000011101100010000000100011;
ROM[2084] <= 32'b00000110100000011010001110000011;
ROM[2085] <= 32'b00000000011100010010000000100011;
ROM[2086] <= 32'b00000000010000010000000100010011;
ROM[2087] <= 32'b00000110111000000000001110010011;
ROM[2088] <= 32'b00000000011100010010000000100011;
ROM[2089] <= 32'b00000000010000010000000100010011;
ROM[2090] <= 32'b00000000000000000010001110110111;
ROM[2091] <= 32'b00001111010000111000001110010011;
ROM[2092] <= 32'b00000000111000111000001110110011;
ROM[2093] <= 32'b00000000011100010010000000100011;
ROM[2094] <= 32'b00000000010000010000000100010011;
ROM[2095] <= 32'b00000000001100010010000000100011;
ROM[2096] <= 32'b00000000010000010000000100010011;
ROM[2097] <= 32'b00000000010000010010000000100011;
ROM[2098] <= 32'b00000000010000010000000100010011;
ROM[2099] <= 32'b00000000010100010010000000100011;
ROM[2100] <= 32'b00000000010000010000000100010011;
ROM[2101] <= 32'b00000000011000010010000000100011;
ROM[2102] <= 32'b00000000010000010000000100010011;
ROM[2103] <= 32'b00000001010000000000001110010011;
ROM[2104] <= 32'b00000000100000111000001110010011;
ROM[2105] <= 32'b01000000011100010000001110110011;
ROM[2106] <= 32'b00000000011100000000001000110011;
ROM[2107] <= 32'b00000000001000000000000110110011;
ROM[2108] <= 32'b00111100110100001111000011101111;
ROM[2109] <= 32'b11111111110000010000000100010011;
ROM[2110] <= 32'b00000000000000010010001110000011;
ROM[2111] <= 32'b00000000011101100010000000100011;
ROM[2112] <= 32'b00000110100000011010001110000011;
ROM[2113] <= 32'b00000000011100010010000000100011;
ROM[2114] <= 32'b00000000010000010000000100010011;
ROM[2115] <= 32'b00000111010000000000001110010011;
ROM[2116] <= 32'b00000000011100010010000000100011;
ROM[2117] <= 32'b00000000010000010000000100010011;
ROM[2118] <= 32'b00000000000000000010001110110111;
ROM[2119] <= 32'b00010110010000111000001110010011;
ROM[2120] <= 32'b00000000111000111000001110110011;
ROM[2121] <= 32'b00000000011100010010000000100011;
ROM[2122] <= 32'b00000000010000010000000100010011;
ROM[2123] <= 32'b00000000001100010010000000100011;
ROM[2124] <= 32'b00000000010000010000000100010011;
ROM[2125] <= 32'b00000000010000010010000000100011;
ROM[2126] <= 32'b00000000010000010000000100010011;
ROM[2127] <= 32'b00000000010100010010000000100011;
ROM[2128] <= 32'b00000000010000010000000100010011;
ROM[2129] <= 32'b00000000011000010010000000100011;
ROM[2130] <= 32'b00000000010000010000000100010011;
ROM[2131] <= 32'b00000001010000000000001110010011;
ROM[2132] <= 32'b00000000100000111000001110010011;
ROM[2133] <= 32'b01000000011100010000001110110011;
ROM[2134] <= 32'b00000000011100000000001000110011;
ROM[2135] <= 32'b00000000001000000000000110110011;
ROM[2136] <= 32'b00110101110100001111000011101111;
ROM[2137] <= 32'b11111111110000010000000100010011;
ROM[2138] <= 32'b00000000000000010010001110000011;
ROM[2139] <= 32'b00000000011101100010000000100011;
ROM[2140] <= 32'b00000110100000011010001110000011;
ROM[2141] <= 32'b00000000011100010010000000100011;
ROM[2142] <= 32'b00000000010000010000000100010011;
ROM[2143] <= 32'b00000110010100000000001110010011;
ROM[2144] <= 32'b00000000011100010010000000100011;
ROM[2145] <= 32'b00000000010000010000000100010011;
ROM[2146] <= 32'b00000000000000000010001110110111;
ROM[2147] <= 32'b00011101010000111000001110010011;
ROM[2148] <= 32'b00000000111000111000001110110011;
ROM[2149] <= 32'b00000000011100010010000000100011;
ROM[2150] <= 32'b00000000010000010000000100010011;
ROM[2151] <= 32'b00000000001100010010000000100011;
ROM[2152] <= 32'b00000000010000010000000100010011;
ROM[2153] <= 32'b00000000010000010010000000100011;
ROM[2154] <= 32'b00000000010000010000000100010011;
ROM[2155] <= 32'b00000000010100010010000000100011;
ROM[2156] <= 32'b00000000010000010000000100010011;
ROM[2157] <= 32'b00000000011000010010000000100011;
ROM[2158] <= 32'b00000000010000010000000100010011;
ROM[2159] <= 32'b00000001010000000000001110010011;
ROM[2160] <= 32'b00000000100000111000001110010011;
ROM[2161] <= 32'b01000000011100010000001110110011;
ROM[2162] <= 32'b00000000011100000000001000110011;
ROM[2163] <= 32'b00000000001000000000000110110011;
ROM[2164] <= 32'b00101110110100001111000011101111;
ROM[2165] <= 32'b11111111110000010000000100010011;
ROM[2166] <= 32'b00000000000000010010001110000011;
ROM[2167] <= 32'b00000000011101100010000000100011;
ROM[2168] <= 32'b00000110100000011010001110000011;
ROM[2169] <= 32'b00000000011100010010000000100011;
ROM[2170] <= 32'b00000000010000010000000100010011;
ROM[2171] <= 32'b00000111001000000000001110010011;
ROM[2172] <= 32'b00000000011100010010000000100011;
ROM[2173] <= 32'b00000000010000010000000100010011;
ROM[2174] <= 32'b00000000000000000010001110110111;
ROM[2175] <= 32'b00100100010000111000001110010011;
ROM[2176] <= 32'b00000000111000111000001110110011;
ROM[2177] <= 32'b00000000011100010010000000100011;
ROM[2178] <= 32'b00000000010000010000000100010011;
ROM[2179] <= 32'b00000000001100010010000000100011;
ROM[2180] <= 32'b00000000010000010000000100010011;
ROM[2181] <= 32'b00000000010000010010000000100011;
ROM[2182] <= 32'b00000000010000010000000100010011;
ROM[2183] <= 32'b00000000010100010010000000100011;
ROM[2184] <= 32'b00000000010000010000000100010011;
ROM[2185] <= 32'b00000000011000010010000000100011;
ROM[2186] <= 32'b00000000010000010000000100010011;
ROM[2187] <= 32'b00000001010000000000001110010011;
ROM[2188] <= 32'b00000000100000111000001110010011;
ROM[2189] <= 32'b01000000011100010000001110110011;
ROM[2190] <= 32'b00000000011100000000001000110011;
ROM[2191] <= 32'b00000000001000000000000110110011;
ROM[2192] <= 32'b00100111110100001111000011101111;
ROM[2193] <= 32'b11111111110000010000000100010011;
ROM[2194] <= 32'b00000000000000010010001110000011;
ROM[2195] <= 32'b00000000011101100010000000100011;
ROM[2196] <= 32'b00000110100000011010001110000011;
ROM[2197] <= 32'b00000000011100010010000000100011;
ROM[2198] <= 32'b00000000010000010000000100010011;
ROM[2199] <= 32'b00000011101000000000001110010011;
ROM[2200] <= 32'b00000000011100010010000000100011;
ROM[2201] <= 32'b00000000010000010000000100010011;
ROM[2202] <= 32'b00000000000000000010001110110111;
ROM[2203] <= 32'b00101011010000111000001110010011;
ROM[2204] <= 32'b00000000111000111000001110110011;
ROM[2205] <= 32'b00000000011100010010000000100011;
ROM[2206] <= 32'b00000000010000010000000100010011;
ROM[2207] <= 32'b00000000001100010010000000100011;
ROM[2208] <= 32'b00000000010000010000000100010011;
ROM[2209] <= 32'b00000000010000010010000000100011;
ROM[2210] <= 32'b00000000010000010000000100010011;
ROM[2211] <= 32'b00000000010100010010000000100011;
ROM[2212] <= 32'b00000000010000010000000100010011;
ROM[2213] <= 32'b00000000011000010010000000100011;
ROM[2214] <= 32'b00000000010000010000000100010011;
ROM[2215] <= 32'b00000001010000000000001110010011;
ROM[2216] <= 32'b00000000100000111000001110010011;
ROM[2217] <= 32'b01000000011100010000001110110011;
ROM[2218] <= 32'b00000000011100000000001000110011;
ROM[2219] <= 32'b00000000001000000000000110110011;
ROM[2220] <= 32'b00100000110100001111000011101111;
ROM[2221] <= 32'b11111111110000010000000100010011;
ROM[2222] <= 32'b00000000000000010010001110000011;
ROM[2223] <= 32'b00000000011101100010000000100011;
ROM[2224] <= 32'b00000110100000011010001110000011;
ROM[2225] <= 32'b00000000011100010010000000100011;
ROM[2226] <= 32'b00000000010000010000000100010011;
ROM[2227] <= 32'b00000010000000000000001110010011;
ROM[2228] <= 32'b00000000011100010010000000100011;
ROM[2229] <= 32'b00000000010000010000000100010011;
ROM[2230] <= 32'b00000000000000000010001110110111;
ROM[2231] <= 32'b00110010010000111000001110010011;
ROM[2232] <= 32'b00000000111000111000001110110011;
ROM[2233] <= 32'b00000000011100010010000000100011;
ROM[2234] <= 32'b00000000010000010000000100010011;
ROM[2235] <= 32'b00000000001100010010000000100011;
ROM[2236] <= 32'b00000000010000010000000100010011;
ROM[2237] <= 32'b00000000010000010010000000100011;
ROM[2238] <= 32'b00000000010000010000000100010011;
ROM[2239] <= 32'b00000000010100010010000000100011;
ROM[2240] <= 32'b00000000010000010000000100010011;
ROM[2241] <= 32'b00000000011000010010000000100011;
ROM[2242] <= 32'b00000000010000010000000100010011;
ROM[2243] <= 32'b00000001010000000000001110010011;
ROM[2244] <= 32'b00000000100000111000001110010011;
ROM[2245] <= 32'b01000000011100010000001110110011;
ROM[2246] <= 32'b00000000011100000000001000110011;
ROM[2247] <= 32'b00000000001000000000000110110011;
ROM[2248] <= 32'b00011001110100001111000011101111;
ROM[2249] <= 32'b11111111110000010000000100010011;
ROM[2250] <= 32'b00000000000000010010001110000011;
ROM[2251] <= 32'b00000000011101100010000000100011;
ROM[2252] <= 32'b00000110100000011010001110000011;
ROM[2253] <= 32'b00000110011100011010010000100011;
ROM[2254] <= 32'b00000000010100000000001110010011;
ROM[2255] <= 32'b00000000011100010010000000100011;
ROM[2256] <= 32'b00000000010000010000000100010011;
ROM[2257] <= 32'b00000000000000000010001110110111;
ROM[2258] <= 32'b00111001000000111000001110010011;
ROM[2259] <= 32'b00000000111000111000001110110011;
ROM[2260] <= 32'b00000000011100010010000000100011;
ROM[2261] <= 32'b00000000010000010000000100010011;
ROM[2262] <= 32'b00000000001100010010000000100011;
ROM[2263] <= 32'b00000000010000010000000100010011;
ROM[2264] <= 32'b00000000010000010010000000100011;
ROM[2265] <= 32'b00000000010000010000000100010011;
ROM[2266] <= 32'b00000000010100010010000000100011;
ROM[2267] <= 32'b00000000010000010000000100010011;
ROM[2268] <= 32'b00000000011000010010000000100011;
ROM[2269] <= 32'b00000000010000010000000100010011;
ROM[2270] <= 32'b00000001010000000000001110010011;
ROM[2271] <= 32'b00000000010000111000001110010011;
ROM[2272] <= 32'b01000000011100010000001110110011;
ROM[2273] <= 32'b00000000011100000000001000110011;
ROM[2274] <= 32'b00000000001000000000000110110011;
ROM[2275] <= 32'b01010111010000001111000011101111;
ROM[2276] <= 32'b11111111110000010000000100010011;
ROM[2277] <= 32'b00000000000000010010001110000011;
ROM[2278] <= 32'b00000110011100011010011000100011;
ROM[2279] <= 32'b00000110110000011010001110000011;
ROM[2280] <= 32'b00000000011100010010000000100011;
ROM[2281] <= 32'b00000000010000010000000100010011;
ROM[2282] <= 32'b00000110111100000000001110010011;
ROM[2283] <= 32'b00000000011100010010000000100011;
ROM[2284] <= 32'b00000000010000010000000100010011;
ROM[2285] <= 32'b00000000000000000010001110110111;
ROM[2286] <= 32'b01000000000000111000001110010011;
ROM[2287] <= 32'b00000000111000111000001110110011;
ROM[2288] <= 32'b00000000011100010010000000100011;
ROM[2289] <= 32'b00000000010000010000000100010011;
ROM[2290] <= 32'b00000000001100010010000000100011;
ROM[2291] <= 32'b00000000010000010000000100010011;
ROM[2292] <= 32'b00000000010000010010000000100011;
ROM[2293] <= 32'b00000000010000010000000100010011;
ROM[2294] <= 32'b00000000010100010010000000100011;
ROM[2295] <= 32'b00000000010000010000000100010011;
ROM[2296] <= 32'b00000000011000010010000000100011;
ROM[2297] <= 32'b00000000010000010000000100010011;
ROM[2298] <= 32'b00000001010000000000001110010011;
ROM[2299] <= 32'b00000000100000111000001110010011;
ROM[2300] <= 32'b01000000011100010000001110110011;
ROM[2301] <= 32'b00000000011100000000001000110011;
ROM[2302] <= 32'b00000000001000000000000110110011;
ROM[2303] <= 32'b00001100000100001111000011101111;
ROM[2304] <= 32'b11111111110000010000000100010011;
ROM[2305] <= 32'b00000000000000010010001110000011;
ROM[2306] <= 32'b00000000011101100010000000100011;
ROM[2307] <= 32'b00000110110000011010001110000011;
ROM[2308] <= 32'b00000000011100010010000000100011;
ROM[2309] <= 32'b00000000010000010000000100010011;
ROM[2310] <= 32'b00000111011000000000001110010011;
ROM[2311] <= 32'b00000000011100010010000000100011;
ROM[2312] <= 32'b00000000010000010000000100010011;
ROM[2313] <= 32'b00000000000000000010001110110111;
ROM[2314] <= 32'b01000111000000111000001110010011;
ROM[2315] <= 32'b00000000111000111000001110110011;
ROM[2316] <= 32'b00000000011100010010000000100011;
ROM[2317] <= 32'b00000000010000010000000100010011;
ROM[2318] <= 32'b00000000001100010010000000100011;
ROM[2319] <= 32'b00000000010000010000000100010011;
ROM[2320] <= 32'b00000000010000010010000000100011;
ROM[2321] <= 32'b00000000010000010000000100010011;
ROM[2322] <= 32'b00000000010100010010000000100011;
ROM[2323] <= 32'b00000000010000010000000100010011;
ROM[2324] <= 32'b00000000011000010010000000100011;
ROM[2325] <= 32'b00000000010000010000000100010011;
ROM[2326] <= 32'b00000001010000000000001110010011;
ROM[2327] <= 32'b00000000100000111000001110010011;
ROM[2328] <= 32'b01000000011100010000001110110011;
ROM[2329] <= 32'b00000000011100000000001000110011;
ROM[2330] <= 32'b00000000001000000000000110110011;
ROM[2331] <= 32'b00000101000100001111000011101111;
ROM[2332] <= 32'b11111111110000010000000100010011;
ROM[2333] <= 32'b00000000000000010010001110000011;
ROM[2334] <= 32'b00000000011101100010000000100011;
ROM[2335] <= 32'b00000110110000011010001110000011;
ROM[2336] <= 32'b00000000011100010010000000100011;
ROM[2337] <= 32'b00000000010000010000000100010011;
ROM[2338] <= 32'b00000110010100000000001110010011;
ROM[2339] <= 32'b00000000011100010010000000100011;
ROM[2340] <= 32'b00000000010000010000000100010011;
ROM[2341] <= 32'b00000000000000000010001110110111;
ROM[2342] <= 32'b01001110000000111000001110010011;
ROM[2343] <= 32'b00000000111000111000001110110011;
ROM[2344] <= 32'b00000000011100010010000000100011;
ROM[2345] <= 32'b00000000010000010000000100010011;
ROM[2346] <= 32'b00000000001100010010000000100011;
ROM[2347] <= 32'b00000000010000010000000100010011;
ROM[2348] <= 32'b00000000010000010010000000100011;
ROM[2349] <= 32'b00000000010000010000000100010011;
ROM[2350] <= 32'b00000000010100010010000000100011;
ROM[2351] <= 32'b00000000010000010000000100010011;
ROM[2352] <= 32'b00000000011000010010000000100011;
ROM[2353] <= 32'b00000000010000010000000100010011;
ROM[2354] <= 32'b00000001010000000000001110010011;
ROM[2355] <= 32'b00000000100000111000001110010011;
ROM[2356] <= 32'b01000000011100010000001110110011;
ROM[2357] <= 32'b00000000011100000000001000110011;
ROM[2358] <= 32'b00000000001000000000000110110011;
ROM[2359] <= 32'b01111110000000001111000011101111;
ROM[2360] <= 32'b11111111110000010000000100010011;
ROM[2361] <= 32'b00000000000000010010001110000011;
ROM[2362] <= 32'b00000000011101100010000000100011;
ROM[2363] <= 32'b00000110110000011010001110000011;
ROM[2364] <= 32'b00000000011100010010000000100011;
ROM[2365] <= 32'b00000000010000010000000100010011;
ROM[2366] <= 32'b00000111001000000000001110010011;
ROM[2367] <= 32'b00000000011100010010000000100011;
ROM[2368] <= 32'b00000000010000010000000100010011;
ROM[2369] <= 32'b00000000000000000010001110110111;
ROM[2370] <= 32'b01010101000000111000001110010011;
ROM[2371] <= 32'b00000000111000111000001110110011;
ROM[2372] <= 32'b00000000011100010010000000100011;
ROM[2373] <= 32'b00000000010000010000000100010011;
ROM[2374] <= 32'b00000000001100010010000000100011;
ROM[2375] <= 32'b00000000010000010000000100010011;
ROM[2376] <= 32'b00000000010000010010000000100011;
ROM[2377] <= 32'b00000000010000010000000100010011;
ROM[2378] <= 32'b00000000010100010010000000100011;
ROM[2379] <= 32'b00000000010000010000000100010011;
ROM[2380] <= 32'b00000000011000010010000000100011;
ROM[2381] <= 32'b00000000010000010000000100010011;
ROM[2382] <= 32'b00000001010000000000001110010011;
ROM[2383] <= 32'b00000000100000111000001110010011;
ROM[2384] <= 32'b01000000011100010000001110110011;
ROM[2385] <= 32'b00000000011100000000001000110011;
ROM[2386] <= 32'b00000000001000000000000110110011;
ROM[2387] <= 32'b01110111000000001111000011101111;
ROM[2388] <= 32'b11111111110000010000000100010011;
ROM[2389] <= 32'b00000000000000010010001110000011;
ROM[2390] <= 32'b00000000011101100010000000100011;
ROM[2391] <= 32'b00000110110000011010001110000011;
ROM[2392] <= 32'b00000000011100010010000000100011;
ROM[2393] <= 32'b00000000010000010000000100010011;
ROM[2394] <= 32'b00000010000100000000001110010011;
ROM[2395] <= 32'b00000000011100010010000000100011;
ROM[2396] <= 32'b00000000010000010000000100010011;
ROM[2397] <= 32'b00000000000000000010001110110111;
ROM[2398] <= 32'b01011100000000111000001110010011;
ROM[2399] <= 32'b00000000111000111000001110110011;
ROM[2400] <= 32'b00000000011100010010000000100011;
ROM[2401] <= 32'b00000000010000010000000100010011;
ROM[2402] <= 32'b00000000001100010010000000100011;
ROM[2403] <= 32'b00000000010000010000000100010011;
ROM[2404] <= 32'b00000000010000010010000000100011;
ROM[2405] <= 32'b00000000010000010000000100010011;
ROM[2406] <= 32'b00000000010100010010000000100011;
ROM[2407] <= 32'b00000000010000010000000100010011;
ROM[2408] <= 32'b00000000011000010010000000100011;
ROM[2409] <= 32'b00000000010000010000000100010011;
ROM[2410] <= 32'b00000001010000000000001110010011;
ROM[2411] <= 32'b00000000100000111000001110010011;
ROM[2412] <= 32'b01000000011100010000001110110011;
ROM[2413] <= 32'b00000000011100000000001000110011;
ROM[2414] <= 32'b00000000001000000000000110110011;
ROM[2415] <= 32'b01110000000000001111000011101111;
ROM[2416] <= 32'b11111111110000010000000100010011;
ROM[2417] <= 32'b00000000000000010010001110000011;
ROM[2418] <= 32'b00000000011101100010000000100011;
ROM[2419] <= 32'b00000110110000011010001110000011;
ROM[2420] <= 32'b00000110011100011010011000100011;
ROM[2421] <= 32'b00000000010100000000001110010011;
ROM[2422] <= 32'b00000000011100010010000000100011;
ROM[2423] <= 32'b00000000010000010000000100010011;
ROM[2424] <= 32'b00000000000000000010001110110111;
ROM[2425] <= 32'b01100010110000111000001110010011;
ROM[2426] <= 32'b00000000111000111000001110110011;
ROM[2427] <= 32'b00000000011100010010000000100011;
ROM[2428] <= 32'b00000000010000010000000100010011;
ROM[2429] <= 32'b00000000001100010010000000100011;
ROM[2430] <= 32'b00000000010000010000000100010011;
ROM[2431] <= 32'b00000000010000010010000000100011;
ROM[2432] <= 32'b00000000010000010000000100010011;
ROM[2433] <= 32'b00000000010100010010000000100011;
ROM[2434] <= 32'b00000000010000010000000100010011;
ROM[2435] <= 32'b00000000011000010010000000100011;
ROM[2436] <= 32'b00000000010000010000000100010011;
ROM[2437] <= 32'b00000001010000000000001110010011;
ROM[2438] <= 32'b00000000010000111000001110010011;
ROM[2439] <= 32'b01000000011100010000001110110011;
ROM[2440] <= 32'b00000000011100000000001000110011;
ROM[2441] <= 32'b00000000001000000000000110110011;
ROM[2442] <= 32'b00101101100000001111000011101111;
ROM[2443] <= 32'b11111111110000010000000100010011;
ROM[2444] <= 32'b00000000000000010010001110000011;
ROM[2445] <= 32'b00000110011100011010100000100011;
ROM[2446] <= 32'b00000111000000011010001110000011;
ROM[2447] <= 32'b00000000011100010010000000100011;
ROM[2448] <= 32'b00000000010000010000000100010011;
ROM[2449] <= 32'b00000101011100000000001110010011;
ROM[2450] <= 32'b00000000011100010010000000100011;
ROM[2451] <= 32'b00000000010000010000000100010011;
ROM[2452] <= 32'b00000000000000000010001110110111;
ROM[2453] <= 32'b01101001110000111000001110010011;
ROM[2454] <= 32'b00000000111000111000001110110011;
ROM[2455] <= 32'b00000000011100010010000000100011;
ROM[2456] <= 32'b00000000010000010000000100010011;
ROM[2457] <= 32'b00000000001100010010000000100011;
ROM[2458] <= 32'b00000000010000010000000100010011;
ROM[2459] <= 32'b00000000010000010010000000100011;
ROM[2460] <= 32'b00000000010000010000000100010011;
ROM[2461] <= 32'b00000000010100010010000000100011;
ROM[2462] <= 32'b00000000010000010000000100010011;
ROM[2463] <= 32'b00000000011000010010000000100011;
ROM[2464] <= 32'b00000000010000010000000100010011;
ROM[2465] <= 32'b00000001010000000000001110010011;
ROM[2466] <= 32'b00000000100000111000001110010011;
ROM[2467] <= 32'b01000000011100010000001110110011;
ROM[2468] <= 32'b00000000011100000000001000110011;
ROM[2469] <= 32'b00000000001000000000000110110011;
ROM[2470] <= 32'b01100010010000001111000011101111;
ROM[2471] <= 32'b11111111110000010000000100010011;
ROM[2472] <= 32'b00000000000000010010001110000011;
ROM[2473] <= 32'b00000000011101100010000000100011;
ROM[2474] <= 32'b00000111000000011010001110000011;
ROM[2475] <= 32'b00000000011100010010000000100011;
ROM[2476] <= 32'b00000000010000010000000100010011;
ROM[2477] <= 32'b00000110111100000000001110010011;
ROM[2478] <= 32'b00000000011100010010000000100011;
ROM[2479] <= 32'b00000000010000010000000100010011;
ROM[2480] <= 32'b00000000000000000010001110110111;
ROM[2481] <= 32'b01110000110000111000001110010011;
ROM[2482] <= 32'b00000000111000111000001110110011;
ROM[2483] <= 32'b00000000011100010010000000100011;
ROM[2484] <= 32'b00000000010000010000000100010011;
ROM[2485] <= 32'b00000000001100010010000000100011;
ROM[2486] <= 32'b00000000010000010000000100010011;
ROM[2487] <= 32'b00000000010000010010000000100011;
ROM[2488] <= 32'b00000000010000010000000100010011;
ROM[2489] <= 32'b00000000010100010010000000100011;
ROM[2490] <= 32'b00000000010000010000000100010011;
ROM[2491] <= 32'b00000000011000010010000000100011;
ROM[2492] <= 32'b00000000010000010000000100010011;
ROM[2493] <= 32'b00000001010000000000001110010011;
ROM[2494] <= 32'b00000000100000111000001110010011;
ROM[2495] <= 32'b01000000011100010000001110110011;
ROM[2496] <= 32'b00000000011100000000001000110011;
ROM[2497] <= 32'b00000000001000000000000110110011;
ROM[2498] <= 32'b01011011010000001111000011101111;
ROM[2499] <= 32'b11111111110000010000000100010011;
ROM[2500] <= 32'b00000000000000010010001110000011;
ROM[2501] <= 32'b00000000011101100010000000100011;
ROM[2502] <= 32'b00000111000000011010001110000011;
ROM[2503] <= 32'b00000000011100010010000000100011;
ROM[2504] <= 32'b00000000010000010000000100010011;
ROM[2505] <= 32'b00000111001000000000001110010011;
ROM[2506] <= 32'b00000000011100010010000000100011;
ROM[2507] <= 32'b00000000010000010000000100010011;
ROM[2508] <= 32'b00000000000000000010001110110111;
ROM[2509] <= 32'b01110111110000111000001110010011;
ROM[2510] <= 32'b00000000111000111000001110110011;
ROM[2511] <= 32'b00000000011100010010000000100011;
ROM[2512] <= 32'b00000000010000010000000100010011;
ROM[2513] <= 32'b00000000001100010010000000100011;
ROM[2514] <= 32'b00000000010000010000000100010011;
ROM[2515] <= 32'b00000000010000010010000000100011;
ROM[2516] <= 32'b00000000010000010000000100010011;
ROM[2517] <= 32'b00000000010100010010000000100011;
ROM[2518] <= 32'b00000000010000010000000100010011;
ROM[2519] <= 32'b00000000011000010010000000100011;
ROM[2520] <= 32'b00000000010000010000000100010011;
ROM[2521] <= 32'b00000001010000000000001110010011;
ROM[2522] <= 32'b00000000100000111000001110010011;
ROM[2523] <= 32'b01000000011100010000001110110011;
ROM[2524] <= 32'b00000000011100000000001000110011;
ROM[2525] <= 32'b00000000001000000000000110110011;
ROM[2526] <= 32'b01010100010000001111000011101111;
ROM[2527] <= 32'b11111111110000010000000100010011;
ROM[2528] <= 32'b00000000000000010010001110000011;
ROM[2529] <= 32'b00000000011101100010000000100011;
ROM[2530] <= 32'b00000111000000011010001110000011;
ROM[2531] <= 32'b00000000011100010010000000100011;
ROM[2532] <= 32'b00000000010000010000000100010011;
ROM[2533] <= 32'b00000110010000000000001110010011;
ROM[2534] <= 32'b00000000011100010010000000100011;
ROM[2535] <= 32'b00000000010000010000000100010011;
ROM[2536] <= 32'b00000000000000000010001110110111;
ROM[2537] <= 32'b01111110110000111000001110010011;
ROM[2538] <= 32'b00000000111000111000001110110011;
ROM[2539] <= 32'b00000000011100010010000000100011;
ROM[2540] <= 32'b00000000010000010000000100010011;
ROM[2541] <= 32'b00000000001100010010000000100011;
ROM[2542] <= 32'b00000000010000010000000100010011;
ROM[2543] <= 32'b00000000010000010010000000100011;
ROM[2544] <= 32'b00000000010000010000000100010011;
ROM[2545] <= 32'b00000000010100010010000000100011;
ROM[2546] <= 32'b00000000010000010000000100010011;
ROM[2547] <= 32'b00000000011000010010000000100011;
ROM[2548] <= 32'b00000000010000010000000100010011;
ROM[2549] <= 32'b00000001010000000000001110010011;
ROM[2550] <= 32'b00000000100000111000001110010011;
ROM[2551] <= 32'b01000000011100010000001110110011;
ROM[2552] <= 32'b00000000011100000000001000110011;
ROM[2553] <= 32'b00000000001000000000000110110011;
ROM[2554] <= 32'b01001101010000001111000011101111;
ROM[2555] <= 32'b11111111110000010000000100010011;
ROM[2556] <= 32'b00000000000000010010001110000011;
ROM[2557] <= 32'b00000000011101100010000000100011;
ROM[2558] <= 32'b00000111000000011010001110000011;
ROM[2559] <= 32'b00000000011100010010000000100011;
ROM[2560] <= 32'b00000000010000010000000100010011;
ROM[2561] <= 32'b00000011101000000000001110010011;
ROM[2562] <= 32'b00000000011100010010000000100011;
ROM[2563] <= 32'b00000000010000010000000100010011;
ROM[2564] <= 32'b00000000000000000011001110110111;
ROM[2565] <= 32'b10000101110000111000001110010011;
ROM[2566] <= 32'b00000000111000111000001110110011;
ROM[2567] <= 32'b00000000011100010010000000100011;
ROM[2568] <= 32'b00000000010000010000000100010011;
ROM[2569] <= 32'b00000000001100010010000000100011;
ROM[2570] <= 32'b00000000010000010000000100010011;
ROM[2571] <= 32'b00000000010000010010000000100011;
ROM[2572] <= 32'b00000000010000010000000100010011;
ROM[2573] <= 32'b00000000010100010010000000100011;
ROM[2574] <= 32'b00000000010000010000000100010011;
ROM[2575] <= 32'b00000000011000010010000000100011;
ROM[2576] <= 32'b00000000010000010000000100010011;
ROM[2577] <= 32'b00000001010000000000001110010011;
ROM[2578] <= 32'b00000000100000111000001110010011;
ROM[2579] <= 32'b01000000011100010000001110110011;
ROM[2580] <= 32'b00000000011100000000001000110011;
ROM[2581] <= 32'b00000000001000000000000110110011;
ROM[2582] <= 32'b01000110010000001111000011101111;
ROM[2583] <= 32'b11111111110000010000000100010011;
ROM[2584] <= 32'b00000000000000010010001110000011;
ROM[2585] <= 32'b00000000011101100010000000100011;
ROM[2586] <= 32'b00000111000000011010001110000011;
ROM[2587] <= 32'b00000110011100011010100000100011;
ROM[2588] <= 32'b00000000001100000000001110010011;
ROM[2589] <= 32'b00000000011100010010000000100011;
ROM[2590] <= 32'b00000000010000010000000100010011;
ROM[2591] <= 32'b00000000000000000011001110110111;
ROM[2592] <= 32'b10001100100000111000001110010011;
ROM[2593] <= 32'b00000000111000111000001110110011;
ROM[2594] <= 32'b00000000011100010010000000100011;
ROM[2595] <= 32'b00000000010000010000000100010011;
ROM[2596] <= 32'b00000000001100010010000000100011;
ROM[2597] <= 32'b00000000010000010000000100010011;
ROM[2598] <= 32'b00000000010000010010000000100011;
ROM[2599] <= 32'b00000000010000010000000100010011;
ROM[2600] <= 32'b00000000010100010010000000100011;
ROM[2601] <= 32'b00000000010000010000000100010011;
ROM[2602] <= 32'b00000000011000010010000000100011;
ROM[2603] <= 32'b00000000010000010000000100010011;
ROM[2604] <= 32'b00000001010000000000001110010011;
ROM[2605] <= 32'b00000000010000111000001110010011;
ROM[2606] <= 32'b01000000011100010000001110110011;
ROM[2607] <= 32'b00000000011100000000001000110011;
ROM[2608] <= 32'b00000000001000000000000110110011;
ROM[2609] <= 32'b00000011110000001111000011101111;
ROM[2610] <= 32'b11111111110000010000000100010011;
ROM[2611] <= 32'b00000000000000010010001110000011;
ROM[2612] <= 32'b00000110011100011010101000100011;
ROM[2613] <= 32'b00000111010000011010001110000011;
ROM[2614] <= 32'b00000000011100010010000000100011;
ROM[2615] <= 32'b00000000010000010000000100010011;
ROM[2616] <= 32'b00000111011100000000001110010011;
ROM[2617] <= 32'b00000000011100010010000000100011;
ROM[2618] <= 32'b00000000010000010000000100010011;
ROM[2619] <= 32'b00000000000000000011001110110111;
ROM[2620] <= 32'b10010011100000111000001110010011;
ROM[2621] <= 32'b00000000111000111000001110110011;
ROM[2622] <= 32'b00000000011100010010000000100011;
ROM[2623] <= 32'b00000000010000010000000100010011;
ROM[2624] <= 32'b00000000001100010010000000100011;
ROM[2625] <= 32'b00000000010000010000000100010011;
ROM[2626] <= 32'b00000000010000010010000000100011;
ROM[2627] <= 32'b00000000010000010000000100010011;
ROM[2628] <= 32'b00000000010100010010000000100011;
ROM[2629] <= 32'b00000000010000010000000100010011;
ROM[2630] <= 32'b00000000011000010010000000100011;
ROM[2631] <= 32'b00000000010000010000000100010011;
ROM[2632] <= 32'b00000001010000000000001110010011;
ROM[2633] <= 32'b00000000100000111000001110010011;
ROM[2634] <= 32'b01000000011100010000001110110011;
ROM[2635] <= 32'b00000000011100000000001000110011;
ROM[2636] <= 32'b00000000001000000000000110110011;
ROM[2637] <= 32'b00111000100000001111000011101111;
ROM[2638] <= 32'b11111111110000010000000100010011;
ROM[2639] <= 32'b00000000000000010010001110000011;
ROM[2640] <= 32'b00000000011101100010000000100011;
ROM[2641] <= 32'b00000111010000011010001110000011;
ROM[2642] <= 32'b00000000011100010010000000100011;
ROM[2643] <= 32'b00000000010000010000000100010011;
ROM[2644] <= 32'b00000110100100000000001110010011;
ROM[2645] <= 32'b00000000011100010010000000100011;
ROM[2646] <= 32'b00000000010000010000000100010011;
ROM[2647] <= 32'b00000000000000000011001110110111;
ROM[2648] <= 32'b10011010100000111000001110010011;
ROM[2649] <= 32'b00000000111000111000001110110011;
ROM[2650] <= 32'b00000000011100010010000000100011;
ROM[2651] <= 32'b00000000010000010000000100010011;
ROM[2652] <= 32'b00000000001100010010000000100011;
ROM[2653] <= 32'b00000000010000010000000100010011;
ROM[2654] <= 32'b00000000010000010010000000100011;
ROM[2655] <= 32'b00000000010000010000000100010011;
ROM[2656] <= 32'b00000000010100010010000000100011;
ROM[2657] <= 32'b00000000010000010000000100010011;
ROM[2658] <= 32'b00000000011000010010000000100011;
ROM[2659] <= 32'b00000000010000010000000100010011;
ROM[2660] <= 32'b00000001010000000000001110010011;
ROM[2661] <= 32'b00000000100000111000001110010011;
ROM[2662] <= 32'b01000000011100010000001110110011;
ROM[2663] <= 32'b00000000011100000000001000110011;
ROM[2664] <= 32'b00000000001000000000000110110011;
ROM[2665] <= 32'b00110001100000001111000011101111;
ROM[2666] <= 32'b11111111110000010000000100010011;
ROM[2667] <= 32'b00000000000000010010001110000011;
ROM[2668] <= 32'b00000000011101100010000000100011;
ROM[2669] <= 32'b00000111010000011010001110000011;
ROM[2670] <= 32'b00000000011100010010000000100011;
ROM[2671] <= 32'b00000000010000010000000100010011;
ROM[2672] <= 32'b00000110111000000000001110010011;
ROM[2673] <= 32'b00000000011100010010000000100011;
ROM[2674] <= 32'b00000000010000010000000100010011;
ROM[2675] <= 32'b00000000000000000011001110110111;
ROM[2676] <= 32'b10100001100000111000001110010011;
ROM[2677] <= 32'b00000000111000111000001110110011;
ROM[2678] <= 32'b00000000011100010010000000100011;
ROM[2679] <= 32'b00000000010000010000000100010011;
ROM[2680] <= 32'b00000000001100010010000000100011;
ROM[2681] <= 32'b00000000010000010000000100010011;
ROM[2682] <= 32'b00000000010000010010000000100011;
ROM[2683] <= 32'b00000000010000010000000100010011;
ROM[2684] <= 32'b00000000010100010010000000100011;
ROM[2685] <= 32'b00000000010000010000000100010011;
ROM[2686] <= 32'b00000000011000010010000000100011;
ROM[2687] <= 32'b00000000010000010000000100010011;
ROM[2688] <= 32'b00000001010000000000001110010011;
ROM[2689] <= 32'b00000000100000111000001110010011;
ROM[2690] <= 32'b01000000011100010000001110110011;
ROM[2691] <= 32'b00000000011100000000001000110011;
ROM[2692] <= 32'b00000000001000000000000110110011;
ROM[2693] <= 32'b00101010100000001111000011101111;
ROM[2694] <= 32'b11111111110000010000000100010011;
ROM[2695] <= 32'b00000000000000010010001110000011;
ROM[2696] <= 32'b00000000011101100010000000100011;
ROM[2697] <= 32'b00000111010000011010001110000011;
ROM[2698] <= 32'b00000110011100011010101000100011;
ROM[2699] <= 32'b00000000011000000000001110010011;
ROM[2700] <= 32'b00000000011100010010000000100011;
ROM[2701] <= 32'b00000000010000010000000100010011;
ROM[2702] <= 32'b00000000000000000011001110110111;
ROM[2703] <= 32'b10101000010000111000001110010011;
ROM[2704] <= 32'b00000000111000111000001110110011;
ROM[2705] <= 32'b00000000011100010010000000100011;
ROM[2706] <= 32'b00000000010000010000000100010011;
ROM[2707] <= 32'b00000000001100010010000000100011;
ROM[2708] <= 32'b00000000010000010000000100010011;
ROM[2709] <= 32'b00000000010000010010000000100011;
ROM[2710] <= 32'b00000000010000010000000100010011;
ROM[2711] <= 32'b00000000010100010010000000100011;
ROM[2712] <= 32'b00000000010000010000000100010011;
ROM[2713] <= 32'b00000000011000010010000000100011;
ROM[2714] <= 32'b00000000010000010000000100010011;
ROM[2715] <= 32'b00000001010000000000001110010011;
ROM[2716] <= 32'b00000000010000111000001110010011;
ROM[2717] <= 32'b01000000011100010000001110110011;
ROM[2718] <= 32'b00000000011100000000001000110011;
ROM[2719] <= 32'b00000000001000000000000110110011;
ROM[2720] <= 32'b01101000000100001110000011101111;
ROM[2721] <= 32'b11111111110000010000000100010011;
ROM[2722] <= 32'b00000000000000010010001110000011;
ROM[2723] <= 32'b00000110011100011010110000100011;
ROM[2724] <= 32'b00000111100000011010001110000011;
ROM[2725] <= 32'b00000000011100010010000000100011;
ROM[2726] <= 32'b00000000010000010000000100010011;
ROM[2727] <= 32'b00000101011100000000001110010011;
ROM[2728] <= 32'b00000000011100010010000000100011;
ROM[2729] <= 32'b00000000010000010000000100010011;
ROM[2730] <= 32'b00000000000000000011001110110111;
ROM[2731] <= 32'b10101111010000111000001110010011;
ROM[2732] <= 32'b00000000111000111000001110110011;
ROM[2733] <= 32'b00000000011100010010000000100011;
ROM[2734] <= 32'b00000000010000010000000100010011;
ROM[2735] <= 32'b00000000001100010010000000100011;
ROM[2736] <= 32'b00000000010000010000000100010011;
ROM[2737] <= 32'b00000000010000010010000000100011;
ROM[2738] <= 32'b00000000010000010000000100010011;
ROM[2739] <= 32'b00000000010100010010000000100011;
ROM[2740] <= 32'b00000000010000010000000100010011;
ROM[2741] <= 32'b00000000011000010010000000100011;
ROM[2742] <= 32'b00000000010000010000000100010011;
ROM[2743] <= 32'b00000001010000000000001110010011;
ROM[2744] <= 32'b00000000100000111000001110010011;
ROM[2745] <= 32'b01000000011100010000001110110011;
ROM[2746] <= 32'b00000000011100000000001000110011;
ROM[2747] <= 32'b00000000001000000000000110110011;
ROM[2748] <= 32'b00011100110000001111000011101111;
ROM[2749] <= 32'b11111111110000010000000100010011;
ROM[2750] <= 32'b00000000000000010010001110000011;
ROM[2751] <= 32'b00000000011101100010000000100011;
ROM[2752] <= 32'b00000111100000011010001110000011;
ROM[2753] <= 32'b00000000011100010010000000100011;
ROM[2754] <= 32'b00000000010000010000000100010011;
ROM[2755] <= 32'b00000110111100000000001110010011;
ROM[2756] <= 32'b00000000011100010010000000100011;
ROM[2757] <= 32'b00000000010000010000000100010011;
ROM[2758] <= 32'b00000000000000000011001110110111;
ROM[2759] <= 32'b10110110010000111000001110010011;
ROM[2760] <= 32'b00000000111000111000001110110011;
ROM[2761] <= 32'b00000000011100010010000000100011;
ROM[2762] <= 32'b00000000010000010000000100010011;
ROM[2763] <= 32'b00000000001100010010000000100011;
ROM[2764] <= 32'b00000000010000010000000100010011;
ROM[2765] <= 32'b00000000010000010010000000100011;
ROM[2766] <= 32'b00000000010000010000000100010011;
ROM[2767] <= 32'b00000000010100010010000000100011;
ROM[2768] <= 32'b00000000010000010000000100010011;
ROM[2769] <= 32'b00000000011000010010000000100011;
ROM[2770] <= 32'b00000000010000010000000100010011;
ROM[2771] <= 32'b00000001010000000000001110010011;
ROM[2772] <= 32'b00000000100000111000001110010011;
ROM[2773] <= 32'b01000000011100010000001110110011;
ROM[2774] <= 32'b00000000011100000000001000110011;
ROM[2775] <= 32'b00000000001000000000000110110011;
ROM[2776] <= 32'b00010101110000001111000011101111;
ROM[2777] <= 32'b11111111110000010000000100010011;
ROM[2778] <= 32'b00000000000000010010001110000011;
ROM[2779] <= 32'b00000000011101100010000000100011;
ROM[2780] <= 32'b00000111100000011010001110000011;
ROM[2781] <= 32'b00000000011100010010000000100011;
ROM[2782] <= 32'b00000000010000010000000100010011;
ROM[2783] <= 32'b00000111001000000000001110010011;
ROM[2784] <= 32'b00000000011100010010000000100011;
ROM[2785] <= 32'b00000000010000010000000100010011;
ROM[2786] <= 32'b00000000000000000011001110110111;
ROM[2787] <= 32'b10111101010000111000001110010011;
ROM[2788] <= 32'b00000000111000111000001110110011;
ROM[2789] <= 32'b00000000011100010010000000100011;
ROM[2790] <= 32'b00000000010000010000000100010011;
ROM[2791] <= 32'b00000000001100010010000000100011;
ROM[2792] <= 32'b00000000010000010000000100010011;
ROM[2793] <= 32'b00000000010000010010000000100011;
ROM[2794] <= 32'b00000000010000010000000100010011;
ROM[2795] <= 32'b00000000010100010010000000100011;
ROM[2796] <= 32'b00000000010000010000000100010011;
ROM[2797] <= 32'b00000000011000010010000000100011;
ROM[2798] <= 32'b00000000010000010000000100010011;
ROM[2799] <= 32'b00000001010000000000001110010011;
ROM[2800] <= 32'b00000000100000111000001110010011;
ROM[2801] <= 32'b01000000011100010000001110110011;
ROM[2802] <= 32'b00000000011100000000001000110011;
ROM[2803] <= 32'b00000000001000000000000110110011;
ROM[2804] <= 32'b00001110110000001111000011101111;
ROM[2805] <= 32'b11111111110000010000000100010011;
ROM[2806] <= 32'b00000000000000010010001110000011;
ROM[2807] <= 32'b00000000011101100010000000100011;
ROM[2808] <= 32'b00000111100000011010001110000011;
ROM[2809] <= 32'b00000000011100010010000000100011;
ROM[2810] <= 32'b00000000010000010000000100010011;
ROM[2811] <= 32'b00000110010000000000001110010011;
ROM[2812] <= 32'b00000000011100010010000000100011;
ROM[2813] <= 32'b00000000010000010000000100010011;
ROM[2814] <= 32'b00000000000000000011001110110111;
ROM[2815] <= 32'b11000100010000111000001110010011;
ROM[2816] <= 32'b00000000111000111000001110110011;
ROM[2817] <= 32'b00000000011100010010000000100011;
ROM[2818] <= 32'b00000000010000010000000100010011;
ROM[2819] <= 32'b00000000001100010010000000100011;
ROM[2820] <= 32'b00000000010000010000000100010011;
ROM[2821] <= 32'b00000000010000010010000000100011;
ROM[2822] <= 32'b00000000010000010000000100010011;
ROM[2823] <= 32'b00000000010100010010000000100011;
ROM[2824] <= 32'b00000000010000010000000100010011;
ROM[2825] <= 32'b00000000011000010010000000100011;
ROM[2826] <= 32'b00000000010000010000000100010011;
ROM[2827] <= 32'b00000001010000000000001110010011;
ROM[2828] <= 32'b00000000100000111000001110010011;
ROM[2829] <= 32'b01000000011100010000001110110011;
ROM[2830] <= 32'b00000000011100000000001000110011;
ROM[2831] <= 32'b00000000001000000000000110110011;
ROM[2832] <= 32'b00000111110000001111000011101111;
ROM[2833] <= 32'b11111111110000010000000100010011;
ROM[2834] <= 32'b00000000000000010010001110000011;
ROM[2835] <= 32'b00000000011101100010000000100011;
ROM[2836] <= 32'b00000111100000011010001110000011;
ROM[2837] <= 32'b00000000011100010010000000100011;
ROM[2838] <= 32'b00000000010000010000000100010011;
ROM[2839] <= 32'b00000011101000000000001110010011;
ROM[2840] <= 32'b00000000011100010010000000100011;
ROM[2841] <= 32'b00000000010000010000000100010011;
ROM[2842] <= 32'b00000000000000000011001110110111;
ROM[2843] <= 32'b11001011010000111000001110010011;
ROM[2844] <= 32'b00000000111000111000001110110011;
ROM[2845] <= 32'b00000000011100010010000000100011;
ROM[2846] <= 32'b00000000010000010000000100010011;
ROM[2847] <= 32'b00000000001100010010000000100011;
ROM[2848] <= 32'b00000000010000010000000100010011;
ROM[2849] <= 32'b00000000010000010010000000100011;
ROM[2850] <= 32'b00000000010000010000000100010011;
ROM[2851] <= 32'b00000000010100010010000000100011;
ROM[2852] <= 32'b00000000010000010000000100010011;
ROM[2853] <= 32'b00000000011000010010000000100011;
ROM[2854] <= 32'b00000000010000010000000100010011;
ROM[2855] <= 32'b00000001010000000000001110010011;
ROM[2856] <= 32'b00000000100000111000001110010011;
ROM[2857] <= 32'b01000000011100010000001110110011;
ROM[2858] <= 32'b00000000011100000000001000110011;
ROM[2859] <= 32'b00000000001000000000000110110011;
ROM[2860] <= 32'b00000000110000001111000011101111;
ROM[2861] <= 32'b11111111110000010000000100010011;
ROM[2862] <= 32'b00000000000000010010001110000011;
ROM[2863] <= 32'b00000000011101100010000000100011;
ROM[2864] <= 32'b00000111100000011010001110000011;
ROM[2865] <= 32'b00000000011100010010000000100011;
ROM[2866] <= 32'b00000000010000010000000100010011;
ROM[2867] <= 32'b00000010000000000000001110010011;
ROM[2868] <= 32'b00000000011100010010000000100011;
ROM[2869] <= 32'b00000000010000010000000100010011;
ROM[2870] <= 32'b00000000000000000011001110110111;
ROM[2871] <= 32'b11010010010000111000001110010011;
ROM[2872] <= 32'b00000000111000111000001110110011;
ROM[2873] <= 32'b00000000011100010010000000100011;
ROM[2874] <= 32'b00000000010000010000000100010011;
ROM[2875] <= 32'b00000000001100010010000000100011;
ROM[2876] <= 32'b00000000010000010000000100010011;
ROM[2877] <= 32'b00000000010000010010000000100011;
ROM[2878] <= 32'b00000000010000010000000100010011;
ROM[2879] <= 32'b00000000010100010010000000100011;
ROM[2880] <= 32'b00000000010000010000000100010011;
ROM[2881] <= 32'b00000000011000010010000000100011;
ROM[2882] <= 32'b00000000010000010000000100010011;
ROM[2883] <= 32'b00000001010000000000001110010011;
ROM[2884] <= 32'b00000000100000111000001110010011;
ROM[2885] <= 32'b01000000011100010000001110110011;
ROM[2886] <= 32'b00000000011100000000001000110011;
ROM[2887] <= 32'b00000000001000000000000110110011;
ROM[2888] <= 32'b01111001110100001110000011101111;
ROM[2889] <= 32'b11111111110000010000000100010011;
ROM[2890] <= 32'b00000000000000010010001110000011;
ROM[2891] <= 32'b00000000011101100010000000100011;
ROM[2892] <= 32'b00000111100000011010001110000011;
ROM[2893] <= 32'b00000110011100011010110000100011;
ROM[2894] <= 32'b00000000100000011010001110000011;
ROM[2895] <= 32'b00000000011100010010000000100011;
ROM[2896] <= 32'b00000000010000010000000100010011;
ROM[2897] <= 32'b00000000010100000000001110010011;
ROM[2898] <= 32'b11111111110000010000000100010011;
ROM[2899] <= 32'b00000000000000010010010000000011;
ROM[2900] <= 32'b00000000011101000010001110110011;
ROM[2901] <= 32'b01000000011100000000001110110011;
ROM[2902] <= 32'b00000000000100111000001110010011;
ROM[2903] <= 32'b00000000000000111000101001100011;
ROM[2904] <= 32'b00000000000000000101001110110111;
ROM[2905] <= 32'b00101001000000111000001110010011;
ROM[2906] <= 32'b00000000111000111000001110110011;
ROM[2907] <= 32'b00000000000000111000000011100111;
ROM[2908] <= 32'b00000000011000000000001110010011;
ROM[2909] <= 32'b00000000011100011010110000100011;
ROM[2910] <= 32'b00000001101000000000001110010011;
ROM[2911] <= 32'b00000000011100010010000000100011;
ROM[2912] <= 32'b00000000010000010000000100010011;
ROM[2913] <= 32'b00000000000000000011001110110111;
ROM[2914] <= 32'b11011101000000111000001110010011;
ROM[2915] <= 32'b00000000111000111000001110110011;
ROM[2916] <= 32'b00000000011100010010000000100011;
ROM[2917] <= 32'b00000000010000010000000100010011;
ROM[2918] <= 32'b00000000001100010010000000100011;
ROM[2919] <= 32'b00000000010000010000000100010011;
ROM[2920] <= 32'b00000000010000010010000000100011;
ROM[2921] <= 32'b00000000010000010000000100010011;
ROM[2922] <= 32'b00000000010100010010000000100011;
ROM[2923] <= 32'b00000000010000010000000100010011;
ROM[2924] <= 32'b00000000011000010010000000100011;
ROM[2925] <= 32'b00000000010000010000000100010011;
ROM[2926] <= 32'b00000001010000000000001110010011;
ROM[2927] <= 32'b00000000010000111000001110010011;
ROM[2928] <= 32'b01000000011100010000001110110011;
ROM[2929] <= 32'b00000000011100000000001000110011;
ROM[2930] <= 32'b00000000001000000000000110110011;
ROM[2931] <= 32'b11100111010011111101000011101111;
ROM[2932] <= 32'b11111111110000010000000100010011;
ROM[2933] <= 32'b00000000000000010010001110000011;
ROM[2934] <= 32'b00000000011100011010001000100011;
ROM[2935] <= 32'b00000000000000000000001110010011;
ROM[2936] <= 32'b00000000011100011010011000100011;
ROM[2937] <= 32'b00000000110000011010001110000011;
ROM[2938] <= 32'b00000000011100010010000000100011;
ROM[2939] <= 32'b00000000010000010000000100010011;
ROM[2940] <= 32'b00000001101000000000001110010011;
ROM[2941] <= 32'b11111111110000010000000100010011;
ROM[2942] <= 32'b00000000000000010010010000000011;
ROM[2943] <= 32'b00000000011101000010001110110011;
ROM[2944] <= 32'b01000000011100000000001110110011;
ROM[2945] <= 32'b00000000000100111000001110010011;
ROM[2946] <= 32'b00000000000000111000101001100011;
ROM[2947] <= 32'b00000000000000000011001110110111;
ROM[2948] <= 32'b11101111010000111000001110010011;
ROM[2949] <= 32'b00000000111000111000001110110011;
ROM[2950] <= 32'b00000000000000111000000011100111;
ROM[2951] <= 32'b00000000110000011010001110000011;
ROM[2952] <= 32'b00000000011100010010000000100011;
ROM[2953] <= 32'b00000000010000010000000100010011;
ROM[2954] <= 32'b00000000010000000000001110010011;
ROM[2955] <= 32'b00000000011100010010000000100011;
ROM[2956] <= 32'b00000000010000010000000100010011;
ROM[2957] <= 32'b00000000000000000011001110110111;
ROM[2958] <= 32'b11101000000000111000001110010011;
ROM[2959] <= 32'b00000000111000111000001110110011;
ROM[2960] <= 32'b00000000011100010010000000100011;
ROM[2961] <= 32'b00000000010000010000000100010011;
ROM[2962] <= 32'b00000000001100010010000000100011;
ROM[2963] <= 32'b00000000010000010000000100010011;
ROM[2964] <= 32'b00000000010000010010000000100011;
ROM[2965] <= 32'b00000000010000010000000100010011;
ROM[2966] <= 32'b00000000010100010010000000100011;
ROM[2967] <= 32'b00000000010000010000000100010011;
ROM[2968] <= 32'b00000000011000010010000000100011;
ROM[2969] <= 32'b00000000010000010000000100010011;
ROM[2970] <= 32'b00000001010000000000001110010011;
ROM[2971] <= 32'b00000000100000111000001110010011;
ROM[2972] <= 32'b01000000011100010000001110110011;
ROM[2973] <= 32'b00000000011100000000001000110011;
ROM[2974] <= 32'b00000000001000000000000110110011;
ROM[2975] <= 32'b00100101100000000110000011101111;
ROM[2976] <= 32'b11111111110000010000000100010011;
ROM[2977] <= 32'b00000000000000010010001110000011;
ROM[2978] <= 32'b00000100011100011010001000100011;
ROM[2979] <= 32'b00000100010000011010001110000011;
ROM[2980] <= 32'b00000000011100010010000000100011;
ROM[2981] <= 32'b00000000010000010000000100010011;
ROM[2982] <= 32'b00000000010000011010001110000011;
ROM[2983] <= 32'b11111111110000010000000100010011;
ROM[2984] <= 32'b00000000000000010010010000000011;
ROM[2985] <= 32'b00000000011101000000001110110011;
ROM[2986] <= 32'b00000000011100010010000000100011;
ROM[2987] <= 32'b00000000010000010000000100010011;
ROM[2988] <= 32'b00000000000000000000001110010011;
ROM[2989] <= 32'b00000000011101100010000000100011;
ROM[2990] <= 32'b11111111110000010000000100010011;
ROM[2991] <= 32'b00000000000000010010001110000011;
ROM[2992] <= 32'b00000000000000111000001100010011;
ROM[2993] <= 32'b00000000000001100010001110000011;
ROM[2994] <= 32'b00000000110100110000010000110011;
ROM[2995] <= 32'b00000000011101000010000000100011;
ROM[2996] <= 32'b00000000110000011010001110000011;
ROM[2997] <= 32'b00000000011100010010000000100011;
ROM[2998] <= 32'b00000000010000010000000100010011;
ROM[2999] <= 32'b00000000000100000000001110010011;
ROM[3000] <= 32'b11111111110000010000000100010011;
ROM[3001] <= 32'b00000000000000010010010000000011;
ROM[3002] <= 32'b00000000011101000000001110110011;
ROM[3003] <= 32'b00000000011100011010011000100011;
ROM[3004] <= 32'b11101111010111111111000011101111;
ROM[3005] <= 32'b00000000100000011010001110000011;
ROM[3006] <= 32'b00000000011100010010000000100011;
ROM[3007] <= 32'b00000000010000010000000100010011;
ROM[3008] <= 32'b00000000010000000000001110010011;
ROM[3009] <= 32'b00000000011100010010000000100011;
ROM[3010] <= 32'b00000000010000010000000100010011;
ROM[3011] <= 32'b00000000000000000011001110110111;
ROM[3012] <= 32'b11110101100000111000001110010011;
ROM[3013] <= 32'b00000000111000111000001110110011;
ROM[3014] <= 32'b00000000011100010010000000100011;
ROM[3015] <= 32'b00000000010000010000000100010011;
ROM[3016] <= 32'b00000000001100010010000000100011;
ROM[3017] <= 32'b00000000010000010000000100010011;
ROM[3018] <= 32'b00000000010000010010000000100011;
ROM[3019] <= 32'b00000000010000010000000100010011;
ROM[3020] <= 32'b00000000010100010010000000100011;
ROM[3021] <= 32'b00000000010000010000000100010011;
ROM[3022] <= 32'b00000000011000010010000000100011;
ROM[3023] <= 32'b00000000010000010000000100010011;
ROM[3024] <= 32'b00000001010000000000001110010011;
ROM[3025] <= 32'b00000000100000111000001110010011;
ROM[3026] <= 32'b01000000011100010000001110110011;
ROM[3027] <= 32'b00000000011100000000001000110011;
ROM[3028] <= 32'b00000000001000000000000110110011;
ROM[3029] <= 32'b00011000000000000110000011101111;
ROM[3030] <= 32'b11111111110000010000000100010011;
ROM[3031] <= 32'b00000000000000010010001110000011;
ROM[3032] <= 32'b00000100011100011010010000100011;
ROM[3033] <= 32'b00000100100000011010001110000011;
ROM[3034] <= 32'b00000000011100010010000000100011;
ROM[3035] <= 32'b00000000010000010000000100010011;
ROM[3036] <= 32'b00000100000000011010001110000011;
ROM[3037] <= 32'b11111111110000010000000100010011;
ROM[3038] <= 32'b00000000000000010010010000000011;
ROM[3039] <= 32'b00000000011101000000001110110011;
ROM[3040] <= 32'b00000000000000111000001100010011;
ROM[3041] <= 32'b00000000110100110000010000110011;
ROM[3042] <= 32'b00000000000001000010001110000011;
ROM[3043] <= 32'b00000000011100011010100000100011;
ROM[3044] <= 32'b00000000100000011010001110000011;
ROM[3045] <= 32'b00000000011100010010000000100011;
ROM[3046] <= 32'b00000000010000010000000100010011;
ROM[3047] <= 32'b00000000000000000000001110010011;
ROM[3048] <= 32'b11111111110000010000000100010011;
ROM[3049] <= 32'b00000000000000010010010000000011;
ROM[3050] <= 32'b00000000011101000010010010110011;
ROM[3051] <= 32'b00000000100000111010010100110011;
ROM[3052] <= 32'b00000000101001001000001110110011;
ROM[3053] <= 32'b00000000000100111000001110010011;
ROM[3054] <= 32'b00000000000100111111001110010011;
ROM[3055] <= 32'b00000000000000111000101001100011;
ROM[3056] <= 32'b00000000000000000011001110110111;
ROM[3057] <= 32'b11111101010000111000001110010011;
ROM[3058] <= 32'b00000000111000111000001110110011;
ROM[3059] <= 32'b00000000000000111000000011100111;
ROM[3060] <= 32'b00100011010000000000000011101111;
ROM[3061] <= 32'b00000000010000000000001110010011;
ROM[3062] <= 32'b00000000011100010010000000100011;
ROM[3063] <= 32'b00000000010000010000000100010011;
ROM[3064] <= 32'b00000000000000000011001110110111;
ROM[3065] <= 32'b00000010110000111000001110010011;
ROM[3066] <= 32'b00000000111000111000001110110011;
ROM[3067] <= 32'b00000000011100010010000000100011;
ROM[3068] <= 32'b00000000010000010000000100010011;
ROM[3069] <= 32'b00000000001100010010000000100011;
ROM[3070] <= 32'b00000000010000010000000100010011;
ROM[3071] <= 32'b00000000010000010010000000100011;
ROM[3072] <= 32'b00000000010000010000000100010011;
ROM[3073] <= 32'b00000000010100010010000000100011;
ROM[3074] <= 32'b00000000010000010000000100010011;
ROM[3075] <= 32'b00000000011000010010000000100011;
ROM[3076] <= 32'b00000000010000010000000100010011;
ROM[3077] <= 32'b00000001010000000000001110010011;
ROM[3078] <= 32'b00000000010000111000001110010011;
ROM[3079] <= 32'b01000000011100010000001110110011;
ROM[3080] <= 32'b00000000011100000000001000110011;
ROM[3081] <= 32'b00000000001000000000000110110011;
ROM[3082] <= 32'b00001101100100001110000011101111;
ROM[3083] <= 32'b11111111110000010000000100010011;
ROM[3084] <= 32'b00000000000000010010001110000011;
ROM[3085] <= 32'b00000000011100011010111000100011;
ROM[3086] <= 32'b00000001110000011010001110000011;
ROM[3087] <= 32'b00000000011100010010000000100011;
ROM[3088] <= 32'b00000000010000010000000100010011;
ROM[3089] <= 32'b00000101111100000000001110010011;
ROM[3090] <= 32'b00000000011100010010000000100011;
ROM[3091] <= 32'b00000000010000010000000100010011;
ROM[3092] <= 32'b00000000000000000011001110110111;
ROM[3093] <= 32'b00001001110000111000001110010011;
ROM[3094] <= 32'b00000000111000111000001110110011;
ROM[3095] <= 32'b00000000011100010010000000100011;
ROM[3096] <= 32'b00000000010000010000000100010011;
ROM[3097] <= 32'b00000000001100010010000000100011;
ROM[3098] <= 32'b00000000010000010000000100010011;
ROM[3099] <= 32'b00000000010000010010000000100011;
ROM[3100] <= 32'b00000000010000010000000100010011;
ROM[3101] <= 32'b00000000010100010010000000100011;
ROM[3102] <= 32'b00000000010000010000000100010011;
ROM[3103] <= 32'b00000000011000010010000000100011;
ROM[3104] <= 32'b00000000010000010000000100010011;
ROM[3105] <= 32'b00000001010000000000001110010011;
ROM[3106] <= 32'b00000000100000111000001110010011;
ROM[3107] <= 32'b01000000011100010000001110110011;
ROM[3108] <= 32'b00000000011100000000001000110011;
ROM[3109] <= 32'b00000000001000000000000110110011;
ROM[3110] <= 32'b01000010010100001110000011101111;
ROM[3111] <= 32'b11111111110000010000000100010011;
ROM[3112] <= 32'b00000000000000010010001110000011;
ROM[3113] <= 32'b00000000011101100010000000100011;
ROM[3114] <= 32'b00000001110000011010001110000011;
ROM[3115] <= 32'b00000000011100010010000000100011;
ROM[3116] <= 32'b00000000010000010000000100010011;
ROM[3117] <= 32'b00000101111100000000001110010011;
ROM[3118] <= 32'b00000000011100010010000000100011;
ROM[3119] <= 32'b00000000010000010000000100010011;
ROM[3120] <= 32'b00000000000000000011001110110111;
ROM[3121] <= 32'b00010000110000111000001110010011;
ROM[3122] <= 32'b00000000111000111000001110110011;
ROM[3123] <= 32'b00000000011100010010000000100011;
ROM[3124] <= 32'b00000000010000010000000100010011;
ROM[3125] <= 32'b00000000001100010010000000100011;
ROM[3126] <= 32'b00000000010000010000000100010011;
ROM[3127] <= 32'b00000000010000010010000000100011;
ROM[3128] <= 32'b00000000010000010000000100010011;
ROM[3129] <= 32'b00000000010100010010000000100011;
ROM[3130] <= 32'b00000000010000010000000100010011;
ROM[3131] <= 32'b00000000011000010010000000100011;
ROM[3132] <= 32'b00000000010000010000000100010011;
ROM[3133] <= 32'b00000001010000000000001110010011;
ROM[3134] <= 32'b00000000100000111000001110010011;
ROM[3135] <= 32'b01000000011100010000001110110011;
ROM[3136] <= 32'b00000000011100000000001000110011;
ROM[3137] <= 32'b00000000001000000000000110110011;
ROM[3138] <= 32'b00111011010100001110000011101111;
ROM[3139] <= 32'b11111111110000010000000100010011;
ROM[3140] <= 32'b00000000000000010010001110000011;
ROM[3141] <= 32'b00000000011101100010000000100011;
ROM[3142] <= 32'b00000001110000011010001110000011;
ROM[3143] <= 32'b00000000011100010010000000100011;
ROM[3144] <= 32'b00000000010000010000000100010011;
ROM[3145] <= 32'b00000101111100000000001110010011;
ROM[3146] <= 32'b00000000011100010010000000100011;
ROM[3147] <= 32'b00000000010000010000000100010011;
ROM[3148] <= 32'b00000000000000000011001110110111;
ROM[3149] <= 32'b00010111110000111000001110010011;
ROM[3150] <= 32'b00000000111000111000001110110011;
ROM[3151] <= 32'b00000000011100010010000000100011;
ROM[3152] <= 32'b00000000010000010000000100010011;
ROM[3153] <= 32'b00000000001100010010000000100011;
ROM[3154] <= 32'b00000000010000010000000100010011;
ROM[3155] <= 32'b00000000010000010010000000100011;
ROM[3156] <= 32'b00000000010000010000000100010011;
ROM[3157] <= 32'b00000000010100010010000000100011;
ROM[3158] <= 32'b00000000010000010000000100010011;
ROM[3159] <= 32'b00000000011000010010000000100011;
ROM[3160] <= 32'b00000000010000010000000100010011;
ROM[3161] <= 32'b00000001010000000000001110010011;
ROM[3162] <= 32'b00000000100000111000001110010011;
ROM[3163] <= 32'b01000000011100010000001110110011;
ROM[3164] <= 32'b00000000011100000000001000110011;
ROM[3165] <= 32'b00000000001000000000000110110011;
ROM[3166] <= 32'b00110100010100001110000011101111;
ROM[3167] <= 32'b11111111110000010000000100010011;
ROM[3168] <= 32'b00000000000000010010001110000011;
ROM[3169] <= 32'b00000000011101100010000000100011;
ROM[3170] <= 32'b00000001110000011010001110000011;
ROM[3171] <= 32'b00000000011100010010000000100011;
ROM[3172] <= 32'b00000000010000010000000100010011;
ROM[3173] <= 32'b00000101111100000000001110010011;
ROM[3174] <= 32'b00000000011100010010000000100011;
ROM[3175] <= 32'b00000000010000010000000100010011;
ROM[3176] <= 32'b00000000000000000011001110110111;
ROM[3177] <= 32'b00011110110000111000001110010011;
ROM[3178] <= 32'b00000000111000111000001110110011;
ROM[3179] <= 32'b00000000011100010010000000100011;
ROM[3180] <= 32'b00000000010000010000000100010011;
ROM[3181] <= 32'b00000000001100010010000000100011;
ROM[3182] <= 32'b00000000010000010000000100010011;
ROM[3183] <= 32'b00000000010000010010000000100011;
ROM[3184] <= 32'b00000000010000010000000100010011;
ROM[3185] <= 32'b00000000010100010010000000100011;
ROM[3186] <= 32'b00000000010000010000000100010011;
ROM[3187] <= 32'b00000000011000010010000000100011;
ROM[3188] <= 32'b00000000010000010000000100010011;
ROM[3189] <= 32'b00000001010000000000001110010011;
ROM[3190] <= 32'b00000000100000111000001110010011;
ROM[3191] <= 32'b01000000011100010000001110110011;
ROM[3192] <= 32'b00000000011100000000001000110011;
ROM[3193] <= 32'b00000000001000000000000110110011;
ROM[3194] <= 32'b00101101010100001110000011101111;
ROM[3195] <= 32'b11111111110000010000000100010011;
ROM[3196] <= 32'b00000000000000010010001110000011;
ROM[3197] <= 32'b00000000011101100010000000100011;
ROM[3198] <= 32'b00000001110000011010001110000011;
ROM[3199] <= 32'b00000000011100011010111000100011;
ROM[3200] <= 32'b00010110110000000001000011101111;
ROM[3201] <= 32'b00000000100000011010001110000011;
ROM[3202] <= 32'b00000000011100010010000000100011;
ROM[3203] <= 32'b00000000010000010000000100010011;
ROM[3204] <= 32'b00000000000100000000001110010011;
ROM[3205] <= 32'b11111111110000010000000100010011;
ROM[3206] <= 32'b00000000000000010010010000000011;
ROM[3207] <= 32'b00000000011101000010010010110011;
ROM[3208] <= 32'b00000000100000111010010100110011;
ROM[3209] <= 32'b00000000101001001000001110110011;
ROM[3210] <= 32'b00000000000100111000001110010011;
ROM[3211] <= 32'b00000000000100111111001110010011;
ROM[3212] <= 32'b00000000000000111000101001100011;
ROM[3213] <= 32'b00000000000000000011001110110111;
ROM[3214] <= 32'b00100100100000111000001110010011;
ROM[3215] <= 32'b00000000111000111000001110110011;
ROM[3216] <= 32'b00000000000000111000000011100111;
ROM[3217] <= 32'b01010100010000000000000011101111;
ROM[3218] <= 32'b00000000101100000000001110010011;
ROM[3219] <= 32'b00000000011100010010000000100011;
ROM[3220] <= 32'b00000000010000010000000100010011;
ROM[3221] <= 32'b00000000000000000011001110110111;
ROM[3222] <= 32'b00101010000000111000001110010011;
ROM[3223] <= 32'b00000000111000111000001110110011;
ROM[3224] <= 32'b00000000011100010010000000100011;
ROM[3225] <= 32'b00000000010000010000000100010011;
ROM[3226] <= 32'b00000000001100010010000000100011;
ROM[3227] <= 32'b00000000010000010000000100010011;
ROM[3228] <= 32'b00000000010000010010000000100011;
ROM[3229] <= 32'b00000000010000010000000100010011;
ROM[3230] <= 32'b00000000010100010010000000100011;
ROM[3231] <= 32'b00000000010000010000000100010011;
ROM[3232] <= 32'b00000000011000010010000000100011;
ROM[3233] <= 32'b00000000010000010000000100010011;
ROM[3234] <= 32'b00000001010000000000001110010011;
ROM[3235] <= 32'b00000000010000111000001110010011;
ROM[3236] <= 32'b01000000011100010000001110110011;
ROM[3237] <= 32'b00000000011100000000001000110011;
ROM[3238] <= 32'b00000000001000000000000110110011;
ROM[3239] <= 32'b01100110010000001110000011101111;
ROM[3240] <= 32'b11111111110000010000000100010011;
ROM[3241] <= 32'b00000000000000010010001110000011;
ROM[3242] <= 32'b00000000011100011010111000100011;
ROM[3243] <= 32'b00000001110000011010001110000011;
ROM[3244] <= 32'b00000000011100010010000000100011;
ROM[3245] <= 32'b00000000010000010000000100010011;
ROM[3246] <= 32'b00000101111100000000001110010011;
ROM[3247] <= 32'b00000000011100010010000000100011;
ROM[3248] <= 32'b00000000010000010000000100010011;
ROM[3249] <= 32'b00000000000000000011001110110111;
ROM[3250] <= 32'b00110001000000111000001110010011;
ROM[3251] <= 32'b00000000111000111000001110110011;
ROM[3252] <= 32'b00000000011100010010000000100011;
ROM[3253] <= 32'b00000000010000010000000100010011;
ROM[3254] <= 32'b00000000001100010010000000100011;
ROM[3255] <= 32'b00000000010000010000000100010011;
ROM[3256] <= 32'b00000000010000010010000000100011;
ROM[3257] <= 32'b00000000010000010000000100010011;
ROM[3258] <= 32'b00000000010100010010000000100011;
ROM[3259] <= 32'b00000000010000010000000100010011;
ROM[3260] <= 32'b00000000011000010010000000100011;
ROM[3261] <= 32'b00000000010000010000000100010011;
ROM[3262] <= 32'b00000001010000000000001110010011;
ROM[3263] <= 32'b00000000100000111000001110010011;
ROM[3264] <= 32'b01000000011100010000001110110011;
ROM[3265] <= 32'b00000000011100000000001000110011;
ROM[3266] <= 32'b00000000001000000000000110110011;
ROM[3267] <= 32'b00011011000100001110000011101111;
ROM[3268] <= 32'b11111111110000010000000100010011;
ROM[3269] <= 32'b00000000000000010010001110000011;
ROM[3270] <= 32'b00000000011101100010000000100011;
ROM[3271] <= 32'b00000001110000011010001110000011;
ROM[3272] <= 32'b00000000011100010010000000100011;
ROM[3273] <= 32'b00000000010000010000000100010011;
ROM[3274] <= 32'b00000101111100000000001110010011;
ROM[3275] <= 32'b00000000011100010010000000100011;
ROM[3276] <= 32'b00000000010000010000000100010011;
ROM[3277] <= 32'b00000000000000000011001110110111;
ROM[3278] <= 32'b00111000000000111000001110010011;
ROM[3279] <= 32'b00000000111000111000001110110011;
ROM[3280] <= 32'b00000000011100010010000000100011;
ROM[3281] <= 32'b00000000010000010000000100010011;
ROM[3282] <= 32'b00000000001100010010000000100011;
ROM[3283] <= 32'b00000000010000010000000100010011;
ROM[3284] <= 32'b00000000010000010010000000100011;
ROM[3285] <= 32'b00000000010000010000000100010011;
ROM[3286] <= 32'b00000000010100010010000000100011;
ROM[3287] <= 32'b00000000010000010000000100010011;
ROM[3288] <= 32'b00000000011000010010000000100011;
ROM[3289] <= 32'b00000000010000010000000100010011;
ROM[3290] <= 32'b00000001010000000000001110010011;
ROM[3291] <= 32'b00000000100000111000001110010011;
ROM[3292] <= 32'b01000000011100010000001110110011;
ROM[3293] <= 32'b00000000011100000000001000110011;
ROM[3294] <= 32'b00000000001000000000000110110011;
ROM[3295] <= 32'b00010100000100001110000011101111;
ROM[3296] <= 32'b11111111110000010000000100010011;
ROM[3297] <= 32'b00000000000000010010001110000011;
ROM[3298] <= 32'b00000000011101100010000000100011;
ROM[3299] <= 32'b00000001110000011010001110000011;
ROM[3300] <= 32'b00000000011100010010000000100011;
ROM[3301] <= 32'b00000000010000010000000100010011;
ROM[3302] <= 32'b00000101111100000000001110010011;
ROM[3303] <= 32'b00000000011100010010000000100011;
ROM[3304] <= 32'b00000000010000010000000100010011;
ROM[3305] <= 32'b00000000000000000011001110110111;
ROM[3306] <= 32'b00111111000000111000001110010011;
ROM[3307] <= 32'b00000000111000111000001110110011;
ROM[3308] <= 32'b00000000011100010010000000100011;
ROM[3309] <= 32'b00000000010000010000000100010011;
ROM[3310] <= 32'b00000000001100010010000000100011;
ROM[3311] <= 32'b00000000010000010000000100010011;
ROM[3312] <= 32'b00000000010000010010000000100011;
ROM[3313] <= 32'b00000000010000010000000100010011;
ROM[3314] <= 32'b00000000010100010010000000100011;
ROM[3315] <= 32'b00000000010000010000000100010011;
ROM[3316] <= 32'b00000000011000010010000000100011;
ROM[3317] <= 32'b00000000010000010000000100010011;
ROM[3318] <= 32'b00000001010000000000001110010011;
ROM[3319] <= 32'b00000000100000111000001110010011;
ROM[3320] <= 32'b01000000011100010000001110110011;
ROM[3321] <= 32'b00000000011100000000001000110011;
ROM[3322] <= 32'b00000000001000000000000110110011;
ROM[3323] <= 32'b00001101000100001110000011101111;
ROM[3324] <= 32'b11111111110000010000000100010011;
ROM[3325] <= 32'b00000000000000010010001110000011;
ROM[3326] <= 32'b00000000011101100010000000100011;
ROM[3327] <= 32'b00000001110000011010001110000011;
ROM[3328] <= 32'b00000000011100010010000000100011;
ROM[3329] <= 32'b00000000010000010000000100010011;
ROM[3330] <= 32'b00000101111100000000001110010011;
ROM[3331] <= 32'b00000000011100010010000000100011;
ROM[3332] <= 32'b00000000010000010000000100010011;
ROM[3333] <= 32'b00000000000000000011001110110111;
ROM[3334] <= 32'b01000110000000111000001110010011;
ROM[3335] <= 32'b00000000111000111000001110110011;
ROM[3336] <= 32'b00000000011100010010000000100011;
ROM[3337] <= 32'b00000000010000010000000100010011;
ROM[3338] <= 32'b00000000001100010010000000100011;
ROM[3339] <= 32'b00000000010000010000000100010011;
ROM[3340] <= 32'b00000000010000010010000000100011;
ROM[3341] <= 32'b00000000010000010000000100010011;
ROM[3342] <= 32'b00000000010100010010000000100011;
ROM[3343] <= 32'b00000000010000010000000100010011;
ROM[3344] <= 32'b00000000011000010010000000100011;
ROM[3345] <= 32'b00000000010000010000000100010011;
ROM[3346] <= 32'b00000001010000000000001110010011;
ROM[3347] <= 32'b00000000100000111000001110010011;
ROM[3348] <= 32'b01000000011100010000001110110011;
ROM[3349] <= 32'b00000000011100000000001000110011;
ROM[3350] <= 32'b00000000001000000000000110110011;
ROM[3351] <= 32'b00000110000100001110000011101111;
ROM[3352] <= 32'b11111111110000010000000100010011;
ROM[3353] <= 32'b00000000000000010010001110000011;
ROM[3354] <= 32'b00000000011101100010000000100011;
ROM[3355] <= 32'b00000001110000011010001110000011;
ROM[3356] <= 32'b00000000011100010010000000100011;
ROM[3357] <= 32'b00000000010000010000000100010011;
ROM[3358] <= 32'b00000101111100000000001110010011;
ROM[3359] <= 32'b00000000011100010010000000100011;
ROM[3360] <= 32'b00000000010000010000000100010011;
ROM[3361] <= 32'b00000000000000000011001110110111;
ROM[3362] <= 32'b01001101000000111000001110010011;
ROM[3363] <= 32'b00000000111000111000001110110011;
ROM[3364] <= 32'b00000000011100010010000000100011;
ROM[3365] <= 32'b00000000010000010000000100010011;
ROM[3366] <= 32'b00000000001100010010000000100011;
ROM[3367] <= 32'b00000000010000010000000100010011;
ROM[3368] <= 32'b00000000010000010010000000100011;
ROM[3369] <= 32'b00000000010000010000000100010011;
ROM[3370] <= 32'b00000000010100010010000000100011;
ROM[3371] <= 32'b00000000010000010000000100010011;
ROM[3372] <= 32'b00000000011000010010000000100011;
ROM[3373] <= 32'b00000000010000010000000100010011;
ROM[3374] <= 32'b00000001010000000000001110010011;
ROM[3375] <= 32'b00000000100000111000001110010011;
ROM[3376] <= 32'b01000000011100010000001110110011;
ROM[3377] <= 32'b00000000011100000000001000110011;
ROM[3378] <= 32'b00000000001000000000000110110011;
ROM[3379] <= 32'b01111111000000001110000011101111;
ROM[3380] <= 32'b11111111110000010000000100010011;
ROM[3381] <= 32'b00000000000000010010001110000011;
ROM[3382] <= 32'b00000000011101100010000000100011;
ROM[3383] <= 32'b00000001110000011010001110000011;
ROM[3384] <= 32'b00000000011100010010000000100011;
ROM[3385] <= 32'b00000000010000010000000100010011;
ROM[3386] <= 32'b00000101111100000000001110010011;
ROM[3387] <= 32'b00000000011100010010000000100011;
ROM[3388] <= 32'b00000000010000010000000100010011;
ROM[3389] <= 32'b00000000000000000011001110110111;
ROM[3390] <= 32'b01010100000000111000001110010011;
ROM[3391] <= 32'b00000000111000111000001110110011;
ROM[3392] <= 32'b00000000011100010010000000100011;
ROM[3393] <= 32'b00000000010000010000000100010011;
ROM[3394] <= 32'b00000000001100010010000000100011;
ROM[3395] <= 32'b00000000010000010000000100010011;
ROM[3396] <= 32'b00000000010000010010000000100011;
ROM[3397] <= 32'b00000000010000010000000100010011;
ROM[3398] <= 32'b00000000010100010010000000100011;
ROM[3399] <= 32'b00000000010000010000000100010011;
ROM[3400] <= 32'b00000000011000010010000000100011;
ROM[3401] <= 32'b00000000010000010000000100010011;
ROM[3402] <= 32'b00000001010000000000001110010011;
ROM[3403] <= 32'b00000000100000111000001110010011;
ROM[3404] <= 32'b01000000011100010000001110110011;
ROM[3405] <= 32'b00000000011100000000001000110011;
ROM[3406] <= 32'b00000000001000000000000110110011;
ROM[3407] <= 32'b01111000000000001110000011101111;
ROM[3408] <= 32'b11111111110000010000000100010011;
ROM[3409] <= 32'b00000000000000010010001110000011;
ROM[3410] <= 32'b00000000011101100010000000100011;
ROM[3411] <= 32'b00000001110000011010001110000011;
ROM[3412] <= 32'b00000000011100010010000000100011;
ROM[3413] <= 32'b00000000010000010000000100010011;
ROM[3414] <= 32'b00000101111100000000001110010011;
ROM[3415] <= 32'b00000000011100010010000000100011;
ROM[3416] <= 32'b00000000010000010000000100010011;
ROM[3417] <= 32'b00000000000000000011001110110111;
ROM[3418] <= 32'b01011011000000111000001110010011;
ROM[3419] <= 32'b00000000111000111000001110110011;
ROM[3420] <= 32'b00000000011100010010000000100011;
ROM[3421] <= 32'b00000000010000010000000100010011;
ROM[3422] <= 32'b00000000001100010010000000100011;
ROM[3423] <= 32'b00000000010000010000000100010011;
ROM[3424] <= 32'b00000000010000010010000000100011;
ROM[3425] <= 32'b00000000010000010000000100010011;
ROM[3426] <= 32'b00000000010100010010000000100011;
ROM[3427] <= 32'b00000000010000010000000100010011;
ROM[3428] <= 32'b00000000011000010010000000100011;
ROM[3429] <= 32'b00000000010000010000000100010011;
ROM[3430] <= 32'b00000001010000000000001110010011;
ROM[3431] <= 32'b00000000100000111000001110010011;
ROM[3432] <= 32'b01000000011100010000001110110011;
ROM[3433] <= 32'b00000000011100000000001000110011;
ROM[3434] <= 32'b00000000001000000000000110110011;
ROM[3435] <= 32'b01110001000000001110000011101111;
ROM[3436] <= 32'b11111111110000010000000100010011;
ROM[3437] <= 32'b00000000000000010010001110000011;
ROM[3438] <= 32'b00000000011101100010000000100011;
ROM[3439] <= 32'b00000001110000011010001110000011;
ROM[3440] <= 32'b00000000011100010010000000100011;
ROM[3441] <= 32'b00000000010000010000000100010011;
ROM[3442] <= 32'b00000101111100000000001110010011;
ROM[3443] <= 32'b00000000011100010010000000100011;
ROM[3444] <= 32'b00000000010000010000000100010011;
ROM[3445] <= 32'b00000000000000000011001110110111;
ROM[3446] <= 32'b01100010000000111000001110010011;
ROM[3447] <= 32'b00000000111000111000001110110011;
ROM[3448] <= 32'b00000000011100010010000000100011;
ROM[3449] <= 32'b00000000010000010000000100010011;
ROM[3450] <= 32'b00000000001100010010000000100011;
ROM[3451] <= 32'b00000000010000010000000100010011;
ROM[3452] <= 32'b00000000010000010010000000100011;
ROM[3453] <= 32'b00000000010000010000000100010011;
ROM[3454] <= 32'b00000000010100010010000000100011;
ROM[3455] <= 32'b00000000010000010000000100010011;
ROM[3456] <= 32'b00000000011000010010000000100011;
ROM[3457] <= 32'b00000000010000010000000100010011;
ROM[3458] <= 32'b00000001010000000000001110010011;
ROM[3459] <= 32'b00000000100000111000001110010011;
ROM[3460] <= 32'b01000000011100010000001110110011;
ROM[3461] <= 32'b00000000011100000000001000110011;
ROM[3462] <= 32'b00000000001000000000000110110011;
ROM[3463] <= 32'b01101010000000001110000011101111;
ROM[3464] <= 32'b11111111110000010000000100010011;
ROM[3465] <= 32'b00000000000000010010001110000011;
ROM[3466] <= 32'b00000000011101100010000000100011;
ROM[3467] <= 32'b00000001110000011010001110000011;
ROM[3468] <= 32'b00000000011100010010000000100011;
ROM[3469] <= 32'b00000000010000010000000100010011;
ROM[3470] <= 32'b00000101111100000000001110010011;
ROM[3471] <= 32'b00000000011100010010000000100011;
ROM[3472] <= 32'b00000000010000010000000100010011;
ROM[3473] <= 32'b00000000000000000011001110110111;
ROM[3474] <= 32'b01101001000000111000001110010011;
ROM[3475] <= 32'b00000000111000111000001110110011;
ROM[3476] <= 32'b00000000011100010010000000100011;
ROM[3477] <= 32'b00000000010000010000000100010011;
ROM[3478] <= 32'b00000000001100010010000000100011;
ROM[3479] <= 32'b00000000010000010000000100010011;
ROM[3480] <= 32'b00000000010000010010000000100011;
ROM[3481] <= 32'b00000000010000010000000100010011;
ROM[3482] <= 32'b00000000010100010010000000100011;
ROM[3483] <= 32'b00000000010000010000000100010011;
ROM[3484] <= 32'b00000000011000010010000000100011;
ROM[3485] <= 32'b00000000010000010000000100010011;
ROM[3486] <= 32'b00000001010000000000001110010011;
ROM[3487] <= 32'b00000000100000111000001110010011;
ROM[3488] <= 32'b01000000011100010000001110110011;
ROM[3489] <= 32'b00000000011100000000001000110011;
ROM[3490] <= 32'b00000000001000000000000110110011;
ROM[3491] <= 32'b01100011000000001110000011101111;
ROM[3492] <= 32'b11111111110000010000000100010011;
ROM[3493] <= 32'b00000000000000010010001110000011;
ROM[3494] <= 32'b00000000011101100010000000100011;
ROM[3495] <= 32'b00000001110000011010001110000011;
ROM[3496] <= 32'b00000000011100010010000000100011;
ROM[3497] <= 32'b00000000010000010000000100010011;
ROM[3498] <= 32'b00000101111100000000001110010011;
ROM[3499] <= 32'b00000000011100010010000000100011;
ROM[3500] <= 32'b00000000010000010000000100010011;
ROM[3501] <= 32'b00000000000000000011001110110111;
ROM[3502] <= 32'b01110000000000111000001110010011;
ROM[3503] <= 32'b00000000111000111000001110110011;
ROM[3504] <= 32'b00000000011100010010000000100011;
ROM[3505] <= 32'b00000000010000010000000100010011;
ROM[3506] <= 32'b00000000001100010010000000100011;
ROM[3507] <= 32'b00000000010000010000000100010011;
ROM[3508] <= 32'b00000000010000010010000000100011;
ROM[3509] <= 32'b00000000010000010000000100010011;
ROM[3510] <= 32'b00000000010100010010000000100011;
ROM[3511] <= 32'b00000000010000010000000100010011;
ROM[3512] <= 32'b00000000011000010010000000100011;
ROM[3513] <= 32'b00000000010000010000000100010011;
ROM[3514] <= 32'b00000001010000000000001110010011;
ROM[3515] <= 32'b00000000100000111000001110010011;
ROM[3516] <= 32'b01000000011100010000001110110011;
ROM[3517] <= 32'b00000000011100000000001000110011;
ROM[3518] <= 32'b00000000001000000000000110110011;
ROM[3519] <= 32'b01011100000000001110000011101111;
ROM[3520] <= 32'b11111111110000010000000100010011;
ROM[3521] <= 32'b00000000000000010010001110000011;
ROM[3522] <= 32'b00000000011101100010000000100011;
ROM[3523] <= 32'b00000001110000011010001110000011;
ROM[3524] <= 32'b00000000011100010010000000100011;
ROM[3525] <= 32'b00000000010000010000000100010011;
ROM[3526] <= 32'b00000101111100000000001110010011;
ROM[3527] <= 32'b00000000011100010010000000100011;
ROM[3528] <= 32'b00000000010000010000000100010011;
ROM[3529] <= 32'b00000000000000000011001110110111;
ROM[3530] <= 32'b01110111000000111000001110010011;
ROM[3531] <= 32'b00000000111000111000001110110011;
ROM[3532] <= 32'b00000000011100010010000000100011;
ROM[3533] <= 32'b00000000010000010000000100010011;
ROM[3534] <= 32'b00000000001100010010000000100011;
ROM[3535] <= 32'b00000000010000010000000100010011;
ROM[3536] <= 32'b00000000010000010010000000100011;
ROM[3537] <= 32'b00000000010000010000000100010011;
ROM[3538] <= 32'b00000000010100010010000000100011;
ROM[3539] <= 32'b00000000010000010000000100010011;
ROM[3540] <= 32'b00000000011000010010000000100011;
ROM[3541] <= 32'b00000000010000010000000100010011;
ROM[3542] <= 32'b00000001010000000000001110010011;
ROM[3543] <= 32'b00000000100000111000001110010011;
ROM[3544] <= 32'b01000000011100010000001110110011;
ROM[3545] <= 32'b00000000011100000000001000110011;
ROM[3546] <= 32'b00000000001000000000000110110011;
ROM[3547] <= 32'b01010101000000001110000011101111;
ROM[3548] <= 32'b11111111110000010000000100010011;
ROM[3549] <= 32'b00000000000000010010001110000011;
ROM[3550] <= 32'b00000000011101100010000000100011;
ROM[3551] <= 32'b00000001110000011010001110000011;
ROM[3552] <= 32'b00000000011100011010111000100011;
ROM[3553] <= 32'b00111110100100000000000011101111;
ROM[3554] <= 32'b00000000100000011010001110000011;
ROM[3555] <= 32'b00000000011100010010000000100011;
ROM[3556] <= 32'b00000000010000010000000100010011;
ROM[3557] <= 32'b00000000001000000000001110010011;
ROM[3558] <= 32'b11111111110000010000000100010011;
ROM[3559] <= 32'b00000000000000010010010000000011;
ROM[3560] <= 32'b00000000011101000010010010110011;
ROM[3561] <= 32'b00000000100000111010010100110011;
ROM[3562] <= 32'b00000000101001001000001110110011;
ROM[3563] <= 32'b00000000000100111000001110010011;
ROM[3564] <= 32'b00000000000100111111001110010011;
ROM[3565] <= 32'b00000000000000111000101001100011;
ROM[3566] <= 32'b00000000000000000011001110110111;
ROM[3567] <= 32'b01111100110000111000001110010011;
ROM[3568] <= 32'b00000000111000111000001110110011;
ROM[3569] <= 32'b00000000000000111000000011100111;
ROM[3570] <= 32'b00111111010000000000000011101111;
ROM[3571] <= 32'b00000000100000000000001110010011;
ROM[3572] <= 32'b00000000011100010010000000100011;
ROM[3573] <= 32'b00000000010000010000000100010011;
ROM[3574] <= 32'b00000000000000000100001110110111;
ROM[3575] <= 32'b10000010010000111000001110010011;
ROM[3576] <= 32'b00000000111000111000001110110011;
ROM[3577] <= 32'b00000000011100010010000000100011;
ROM[3578] <= 32'b00000000010000010000000100010011;
ROM[3579] <= 32'b00000000001100010010000000100011;
ROM[3580] <= 32'b00000000010000010000000100010011;
ROM[3581] <= 32'b00000000010000010010000000100011;
ROM[3582] <= 32'b00000000010000010000000100010011;
ROM[3583] <= 32'b00000000010100010010000000100011;
ROM[3584] <= 32'b00000000010000010000000100010011;
ROM[3585] <= 32'b00000000011000010010000000100011;
ROM[3586] <= 32'b00000000010000010000000100010011;
ROM[3587] <= 32'b00000001010000000000001110010011;
ROM[3588] <= 32'b00000000010000111000001110010011;
ROM[3589] <= 32'b01000000011100010000001110110011;
ROM[3590] <= 32'b00000000011100000000001000110011;
ROM[3591] <= 32'b00000000001000000000000110110011;
ROM[3592] <= 32'b00001110000000001110000011101111;
ROM[3593] <= 32'b11111111110000010000000100010011;
ROM[3594] <= 32'b00000000000000010010001110000011;
ROM[3595] <= 32'b00000000011100011010111000100011;
ROM[3596] <= 32'b00000001110000011010001110000011;
ROM[3597] <= 32'b00000000011100010010000000100011;
ROM[3598] <= 32'b00000000010000010000000100010011;
ROM[3599] <= 32'b00000101111100000000001110010011;
ROM[3600] <= 32'b00000000011100010010000000100011;
ROM[3601] <= 32'b00000000010000010000000100010011;
ROM[3602] <= 32'b00000000000000000100001110110111;
ROM[3603] <= 32'b10001001010000111000001110010011;
ROM[3604] <= 32'b00000000111000111000001110110011;
ROM[3605] <= 32'b00000000011100010010000000100011;
ROM[3606] <= 32'b00000000010000010000000100010011;
ROM[3607] <= 32'b00000000001100010010000000100011;
ROM[3608] <= 32'b00000000010000010000000100010011;
ROM[3609] <= 32'b00000000010000010010000000100011;
ROM[3610] <= 32'b00000000010000010000000100010011;
ROM[3611] <= 32'b00000000010100010010000000100011;
ROM[3612] <= 32'b00000000010000010000000100010011;
ROM[3613] <= 32'b00000000011000010010000000100011;
ROM[3614] <= 32'b00000000010000010000000100010011;
ROM[3615] <= 32'b00000001010000000000001110010011;
ROM[3616] <= 32'b00000000100000111000001110010011;
ROM[3617] <= 32'b01000000011100010000001110110011;
ROM[3618] <= 32'b00000000011100000000001000110011;
ROM[3619] <= 32'b00000000001000000000000110110011;
ROM[3620] <= 32'b01000010110000001110000011101111;
ROM[3621] <= 32'b11111111110000010000000100010011;
ROM[3622] <= 32'b00000000000000010010001110000011;
ROM[3623] <= 32'b00000000011101100010000000100011;
ROM[3624] <= 32'b00000001110000011010001110000011;
ROM[3625] <= 32'b00000000011100010010000000100011;
ROM[3626] <= 32'b00000000010000010000000100010011;
ROM[3627] <= 32'b00000101111100000000001110010011;
ROM[3628] <= 32'b00000000011100010010000000100011;
ROM[3629] <= 32'b00000000010000010000000100010011;
ROM[3630] <= 32'b00000000000000000100001110110111;
ROM[3631] <= 32'b10010000010000111000001110010011;
ROM[3632] <= 32'b00000000111000111000001110110011;
ROM[3633] <= 32'b00000000011100010010000000100011;
ROM[3634] <= 32'b00000000010000010000000100010011;
ROM[3635] <= 32'b00000000001100010010000000100011;
ROM[3636] <= 32'b00000000010000010000000100010011;
ROM[3637] <= 32'b00000000010000010010000000100011;
ROM[3638] <= 32'b00000000010000010000000100010011;
ROM[3639] <= 32'b00000000010100010010000000100011;
ROM[3640] <= 32'b00000000010000010000000100010011;
ROM[3641] <= 32'b00000000011000010010000000100011;
ROM[3642] <= 32'b00000000010000010000000100010011;
ROM[3643] <= 32'b00000001010000000000001110010011;
ROM[3644] <= 32'b00000000100000111000001110010011;
ROM[3645] <= 32'b01000000011100010000001110110011;
ROM[3646] <= 32'b00000000011100000000001000110011;
ROM[3647] <= 32'b00000000001000000000000110110011;
ROM[3648] <= 32'b00111011110000001110000011101111;
ROM[3649] <= 32'b11111111110000010000000100010011;
ROM[3650] <= 32'b00000000000000010010001110000011;
ROM[3651] <= 32'b00000000011101100010000000100011;
ROM[3652] <= 32'b00000001110000011010001110000011;
ROM[3653] <= 32'b00000000011100010010000000100011;
ROM[3654] <= 32'b00000000010000010000000100010011;
ROM[3655] <= 32'b00000101111100000000001110010011;
ROM[3656] <= 32'b00000000011100010010000000100011;
ROM[3657] <= 32'b00000000010000010000000100010011;
ROM[3658] <= 32'b00000000000000000100001110110111;
ROM[3659] <= 32'b10010111010000111000001110010011;
ROM[3660] <= 32'b00000000111000111000001110110011;
ROM[3661] <= 32'b00000000011100010010000000100011;
ROM[3662] <= 32'b00000000010000010000000100010011;
ROM[3663] <= 32'b00000000001100010010000000100011;
ROM[3664] <= 32'b00000000010000010000000100010011;
ROM[3665] <= 32'b00000000010000010010000000100011;
ROM[3666] <= 32'b00000000010000010000000100010011;
ROM[3667] <= 32'b00000000010100010010000000100011;
ROM[3668] <= 32'b00000000010000010000000100010011;
ROM[3669] <= 32'b00000000011000010010000000100011;
ROM[3670] <= 32'b00000000010000010000000100010011;
ROM[3671] <= 32'b00000001010000000000001110010011;
ROM[3672] <= 32'b00000000100000111000001110010011;
ROM[3673] <= 32'b01000000011100010000001110110011;
ROM[3674] <= 32'b00000000011100000000001000110011;
ROM[3675] <= 32'b00000000001000000000000110110011;
ROM[3676] <= 32'b00110100110000001110000011101111;
ROM[3677] <= 32'b11111111110000010000000100010011;
ROM[3678] <= 32'b00000000000000010010001110000011;
ROM[3679] <= 32'b00000000011101100010000000100011;
ROM[3680] <= 32'b00000001110000011010001110000011;
ROM[3681] <= 32'b00000000011100010010000000100011;
ROM[3682] <= 32'b00000000010000010000000100010011;
ROM[3683] <= 32'b00000101111100000000001110010011;
ROM[3684] <= 32'b00000000011100010010000000100011;
ROM[3685] <= 32'b00000000010000010000000100010011;
ROM[3686] <= 32'b00000000000000000100001110110111;
ROM[3687] <= 32'b10011110010000111000001110010011;
ROM[3688] <= 32'b00000000111000111000001110110011;
ROM[3689] <= 32'b00000000011100010010000000100011;
ROM[3690] <= 32'b00000000010000010000000100010011;
ROM[3691] <= 32'b00000000001100010010000000100011;
ROM[3692] <= 32'b00000000010000010000000100010011;
ROM[3693] <= 32'b00000000010000010010000000100011;
ROM[3694] <= 32'b00000000010000010000000100010011;
ROM[3695] <= 32'b00000000010100010010000000100011;
ROM[3696] <= 32'b00000000010000010000000100010011;
ROM[3697] <= 32'b00000000011000010010000000100011;
ROM[3698] <= 32'b00000000010000010000000100010011;
ROM[3699] <= 32'b00000001010000000000001110010011;
ROM[3700] <= 32'b00000000100000111000001110010011;
ROM[3701] <= 32'b01000000011100010000001110110011;
ROM[3702] <= 32'b00000000011100000000001000110011;
ROM[3703] <= 32'b00000000001000000000000110110011;
ROM[3704] <= 32'b00101101110000001110000011101111;
ROM[3705] <= 32'b11111111110000010000000100010011;
ROM[3706] <= 32'b00000000000000010010001110000011;
ROM[3707] <= 32'b00000000011101100010000000100011;
ROM[3708] <= 32'b00000001110000011010001110000011;
ROM[3709] <= 32'b00000000011100010010000000100011;
ROM[3710] <= 32'b00000000010000010000000100010011;
ROM[3711] <= 32'b00000101111100000000001110010011;
ROM[3712] <= 32'b00000000011100010010000000100011;
ROM[3713] <= 32'b00000000010000010000000100010011;
ROM[3714] <= 32'b00000000000000000100001110110111;
ROM[3715] <= 32'b10100101010000111000001110010011;
ROM[3716] <= 32'b00000000111000111000001110110011;
ROM[3717] <= 32'b00000000011100010010000000100011;
ROM[3718] <= 32'b00000000010000010000000100010011;
ROM[3719] <= 32'b00000000001100010010000000100011;
ROM[3720] <= 32'b00000000010000010000000100010011;
ROM[3721] <= 32'b00000000010000010010000000100011;
ROM[3722] <= 32'b00000000010000010000000100010011;
ROM[3723] <= 32'b00000000010100010010000000100011;
ROM[3724] <= 32'b00000000010000010000000100010011;
ROM[3725] <= 32'b00000000011000010010000000100011;
ROM[3726] <= 32'b00000000010000010000000100010011;
ROM[3727] <= 32'b00000001010000000000001110010011;
ROM[3728] <= 32'b00000000100000111000001110010011;
ROM[3729] <= 32'b01000000011100010000001110110011;
ROM[3730] <= 32'b00000000011100000000001000110011;
ROM[3731] <= 32'b00000000001000000000000110110011;
ROM[3732] <= 32'b00100110110000001110000011101111;
ROM[3733] <= 32'b11111111110000010000000100010011;
ROM[3734] <= 32'b00000000000000010010001110000011;
ROM[3735] <= 32'b00000000011101100010000000100011;
ROM[3736] <= 32'b00000001110000011010001110000011;
ROM[3737] <= 32'b00000000011100010010000000100011;
ROM[3738] <= 32'b00000000010000010000000100010011;
ROM[3739] <= 32'b00000101111100000000001110010011;
ROM[3740] <= 32'b00000000011100010010000000100011;
ROM[3741] <= 32'b00000000010000010000000100010011;
ROM[3742] <= 32'b00000000000000000100001110110111;
ROM[3743] <= 32'b10101100010000111000001110010011;
ROM[3744] <= 32'b00000000111000111000001110110011;
ROM[3745] <= 32'b00000000011100010010000000100011;
ROM[3746] <= 32'b00000000010000010000000100010011;
ROM[3747] <= 32'b00000000001100010010000000100011;
ROM[3748] <= 32'b00000000010000010000000100010011;
ROM[3749] <= 32'b00000000010000010010000000100011;
ROM[3750] <= 32'b00000000010000010000000100010011;
ROM[3751] <= 32'b00000000010100010010000000100011;
ROM[3752] <= 32'b00000000010000010000000100010011;
ROM[3753] <= 32'b00000000011000010010000000100011;
ROM[3754] <= 32'b00000000010000010000000100010011;
ROM[3755] <= 32'b00000001010000000000001110010011;
ROM[3756] <= 32'b00000000100000111000001110010011;
ROM[3757] <= 32'b01000000011100010000001110110011;
ROM[3758] <= 32'b00000000011100000000001000110011;
ROM[3759] <= 32'b00000000001000000000000110110011;
ROM[3760] <= 32'b00011111110000001110000011101111;
ROM[3761] <= 32'b11111111110000010000000100010011;
ROM[3762] <= 32'b00000000000000010010001110000011;
ROM[3763] <= 32'b00000000011101100010000000100011;
ROM[3764] <= 32'b00000001110000011010001110000011;
ROM[3765] <= 32'b00000000011100010010000000100011;
ROM[3766] <= 32'b00000000010000010000000100010011;
ROM[3767] <= 32'b00000101111100000000001110010011;
ROM[3768] <= 32'b00000000011100010010000000100011;
ROM[3769] <= 32'b00000000010000010000000100010011;
ROM[3770] <= 32'b00000000000000000100001110110111;
ROM[3771] <= 32'b10110011010000111000001110010011;
ROM[3772] <= 32'b00000000111000111000001110110011;
ROM[3773] <= 32'b00000000011100010010000000100011;
ROM[3774] <= 32'b00000000010000010000000100010011;
ROM[3775] <= 32'b00000000001100010010000000100011;
ROM[3776] <= 32'b00000000010000010000000100010011;
ROM[3777] <= 32'b00000000010000010010000000100011;
ROM[3778] <= 32'b00000000010000010000000100010011;
ROM[3779] <= 32'b00000000010100010010000000100011;
ROM[3780] <= 32'b00000000010000010000000100010011;
ROM[3781] <= 32'b00000000011000010010000000100011;
ROM[3782] <= 32'b00000000010000010000000100010011;
ROM[3783] <= 32'b00000001010000000000001110010011;
ROM[3784] <= 32'b00000000100000111000001110010011;
ROM[3785] <= 32'b01000000011100010000001110110011;
ROM[3786] <= 32'b00000000011100000000001000110011;
ROM[3787] <= 32'b00000000001000000000000110110011;
ROM[3788] <= 32'b00011000110000001110000011101111;
ROM[3789] <= 32'b11111111110000010000000100010011;
ROM[3790] <= 32'b00000000000000010010001110000011;
ROM[3791] <= 32'b00000000011101100010000000100011;
ROM[3792] <= 32'b00000001110000011010001110000011;
ROM[3793] <= 32'b00000000011100010010000000100011;
ROM[3794] <= 32'b00000000010000010000000100010011;
ROM[3795] <= 32'b00000101111100000000001110010011;
ROM[3796] <= 32'b00000000011100010010000000100011;
ROM[3797] <= 32'b00000000010000010000000100010011;
ROM[3798] <= 32'b00000000000000000100001110110111;
ROM[3799] <= 32'b10111010010000111000001110010011;
ROM[3800] <= 32'b00000000111000111000001110110011;
ROM[3801] <= 32'b00000000011100010010000000100011;
ROM[3802] <= 32'b00000000010000010000000100010011;
ROM[3803] <= 32'b00000000001100010010000000100011;
ROM[3804] <= 32'b00000000010000010000000100010011;
ROM[3805] <= 32'b00000000010000010010000000100011;
ROM[3806] <= 32'b00000000010000010000000100010011;
ROM[3807] <= 32'b00000000010100010010000000100011;
ROM[3808] <= 32'b00000000010000010000000100010011;
ROM[3809] <= 32'b00000000011000010010000000100011;
ROM[3810] <= 32'b00000000010000010000000100010011;
ROM[3811] <= 32'b00000001010000000000001110010011;
ROM[3812] <= 32'b00000000100000111000001110010011;
ROM[3813] <= 32'b01000000011100010000001110110011;
ROM[3814] <= 32'b00000000011100000000001000110011;
ROM[3815] <= 32'b00000000001000000000000110110011;
ROM[3816] <= 32'b00010001110000001110000011101111;
ROM[3817] <= 32'b11111111110000010000000100010011;
ROM[3818] <= 32'b00000000000000010010001110000011;
ROM[3819] <= 32'b00000000011101100010000000100011;
ROM[3820] <= 32'b00000001110000011010001110000011;
ROM[3821] <= 32'b00000000011100011010111000100011;
ROM[3822] <= 32'b01111011010000000000000011101111;
ROM[3823] <= 32'b00000000100000011010001110000011;
ROM[3824] <= 32'b00000000011100010010000000100011;
ROM[3825] <= 32'b00000000010000010000000100010011;
ROM[3826] <= 32'b00000000001100000000001110010011;
ROM[3827] <= 32'b11111111110000010000000100010011;
ROM[3828] <= 32'b00000000000000010010010000000011;
ROM[3829] <= 32'b00000000011101000010010010110011;
ROM[3830] <= 32'b00000000100000111010010100110011;
ROM[3831] <= 32'b00000000101001001000001110110011;
ROM[3832] <= 32'b00000000000100111000001110010011;
ROM[3833] <= 32'b00000000000100111111001110010011;
ROM[3834] <= 32'b00000000000000111000101001100011;
ROM[3835] <= 32'b00000000000000000100001110110111;
ROM[3836] <= 32'b11000000000000111000001110010011;
ROM[3837] <= 32'b00000000111000111000001110110011;
ROM[3838] <= 32'b00000000000000111000000011100111;
ROM[3839] <= 32'b00111111010000000000000011101111;
ROM[3840] <= 32'b00000000100000000000001110010011;
ROM[3841] <= 32'b00000000011100010010000000100011;
ROM[3842] <= 32'b00000000010000010000000100010011;
ROM[3843] <= 32'b00000000000000000100001110110111;
ROM[3844] <= 32'b11000101100000111000001110010011;
ROM[3845] <= 32'b00000000111000111000001110110011;
ROM[3846] <= 32'b00000000011100010010000000100011;
ROM[3847] <= 32'b00000000010000010000000100010011;
ROM[3848] <= 32'b00000000001100010010000000100011;
ROM[3849] <= 32'b00000000010000010000000100010011;
ROM[3850] <= 32'b00000000010000010010000000100011;
ROM[3851] <= 32'b00000000010000010000000100010011;
ROM[3852] <= 32'b00000000010100010010000000100011;
ROM[3853] <= 32'b00000000010000010000000100010011;
ROM[3854] <= 32'b00000000011000010010000000100011;
ROM[3855] <= 32'b00000000010000010000000100010011;
ROM[3856] <= 32'b00000001010000000000001110010011;
ROM[3857] <= 32'b00000000010000111000001110010011;
ROM[3858] <= 32'b01000000011100010000001110110011;
ROM[3859] <= 32'b00000000011100000000001000110011;
ROM[3860] <= 32'b00000000001000000000000110110011;
ROM[3861] <= 32'b01001010110100001101000011101111;
ROM[3862] <= 32'b11111111110000010000000100010011;
ROM[3863] <= 32'b00000000000000010010001110000011;
ROM[3864] <= 32'b00000000011100011010111000100011;
ROM[3865] <= 32'b00000001110000011010001110000011;
ROM[3866] <= 32'b00000000011100010010000000100011;
ROM[3867] <= 32'b00000000010000010000000100010011;
ROM[3868] <= 32'b00000101111100000000001110010011;
ROM[3869] <= 32'b00000000011100010010000000100011;
ROM[3870] <= 32'b00000000010000010000000100010011;
ROM[3871] <= 32'b00000000000000000100001110110111;
ROM[3872] <= 32'b11001100100000111000001110010011;
ROM[3873] <= 32'b00000000111000111000001110110011;
ROM[3874] <= 32'b00000000011100010010000000100011;
ROM[3875] <= 32'b00000000010000010000000100010011;
ROM[3876] <= 32'b00000000001100010010000000100011;
ROM[3877] <= 32'b00000000010000010000000100010011;
ROM[3878] <= 32'b00000000010000010010000000100011;
ROM[3879] <= 32'b00000000010000010000000100010011;
ROM[3880] <= 32'b00000000010100010010000000100011;
ROM[3881] <= 32'b00000000010000010000000100010011;
ROM[3882] <= 32'b00000000011000010010000000100011;
ROM[3883] <= 32'b00000000010000010000000100010011;
ROM[3884] <= 32'b00000001010000000000001110010011;
ROM[3885] <= 32'b00000000100000111000001110010011;
ROM[3886] <= 32'b01000000011100010000001110110011;
ROM[3887] <= 32'b00000000011100000000001000110011;
ROM[3888] <= 32'b00000000001000000000000110110011;
ROM[3889] <= 32'b01111111100100001101000011101111;
ROM[3890] <= 32'b11111111110000010000000100010011;
ROM[3891] <= 32'b00000000000000010010001110000011;
ROM[3892] <= 32'b00000000011101100010000000100011;
ROM[3893] <= 32'b00000001110000011010001110000011;
ROM[3894] <= 32'b00000000011100010010000000100011;
ROM[3895] <= 32'b00000000010000010000000100010011;
ROM[3896] <= 32'b00000101111100000000001110010011;
ROM[3897] <= 32'b00000000011100010010000000100011;
ROM[3898] <= 32'b00000000010000010000000100010011;
ROM[3899] <= 32'b00000000000000000100001110110111;
ROM[3900] <= 32'b11010011100000111000001110010011;
ROM[3901] <= 32'b00000000111000111000001110110011;
ROM[3902] <= 32'b00000000011100010010000000100011;
ROM[3903] <= 32'b00000000010000010000000100010011;
ROM[3904] <= 32'b00000000001100010010000000100011;
ROM[3905] <= 32'b00000000010000010000000100010011;
ROM[3906] <= 32'b00000000010000010010000000100011;
ROM[3907] <= 32'b00000000010000010000000100010011;
ROM[3908] <= 32'b00000000010100010010000000100011;
ROM[3909] <= 32'b00000000010000010000000100010011;
ROM[3910] <= 32'b00000000011000010010000000100011;
ROM[3911] <= 32'b00000000010000010000000100010011;
ROM[3912] <= 32'b00000001010000000000001110010011;
ROM[3913] <= 32'b00000000100000111000001110010011;
ROM[3914] <= 32'b01000000011100010000001110110011;
ROM[3915] <= 32'b00000000011100000000001000110011;
ROM[3916] <= 32'b00000000001000000000000110110011;
ROM[3917] <= 32'b01111000100100001101000011101111;
ROM[3918] <= 32'b11111111110000010000000100010011;
ROM[3919] <= 32'b00000000000000010010001110000011;
ROM[3920] <= 32'b00000000011101100010000000100011;
ROM[3921] <= 32'b00000001110000011010001110000011;
ROM[3922] <= 32'b00000000011100010010000000100011;
ROM[3923] <= 32'b00000000010000010000000100010011;
ROM[3924] <= 32'b00000101111100000000001110010011;
ROM[3925] <= 32'b00000000011100010010000000100011;
ROM[3926] <= 32'b00000000010000010000000100010011;
ROM[3927] <= 32'b00000000000000000100001110110111;
ROM[3928] <= 32'b11011010100000111000001110010011;
ROM[3929] <= 32'b00000000111000111000001110110011;
ROM[3930] <= 32'b00000000011100010010000000100011;
ROM[3931] <= 32'b00000000010000010000000100010011;
ROM[3932] <= 32'b00000000001100010010000000100011;
ROM[3933] <= 32'b00000000010000010000000100010011;
ROM[3934] <= 32'b00000000010000010010000000100011;
ROM[3935] <= 32'b00000000010000010000000100010011;
ROM[3936] <= 32'b00000000010100010010000000100011;
ROM[3937] <= 32'b00000000010000010000000100010011;
ROM[3938] <= 32'b00000000011000010010000000100011;
ROM[3939] <= 32'b00000000010000010000000100010011;
ROM[3940] <= 32'b00000001010000000000001110010011;
ROM[3941] <= 32'b00000000100000111000001110010011;
ROM[3942] <= 32'b01000000011100010000001110110011;
ROM[3943] <= 32'b00000000011100000000001000110011;
ROM[3944] <= 32'b00000000001000000000000110110011;
ROM[3945] <= 32'b01110001100100001101000011101111;
ROM[3946] <= 32'b11111111110000010000000100010011;
ROM[3947] <= 32'b00000000000000010010001110000011;
ROM[3948] <= 32'b00000000011101100010000000100011;
ROM[3949] <= 32'b00000001110000011010001110000011;
ROM[3950] <= 32'b00000000011100010010000000100011;
ROM[3951] <= 32'b00000000010000010000000100010011;
ROM[3952] <= 32'b00000101111100000000001110010011;
ROM[3953] <= 32'b00000000011100010010000000100011;
ROM[3954] <= 32'b00000000010000010000000100010011;
ROM[3955] <= 32'b00000000000000000100001110110111;
ROM[3956] <= 32'b11100001100000111000001110010011;
ROM[3957] <= 32'b00000000111000111000001110110011;
ROM[3958] <= 32'b00000000011100010010000000100011;
ROM[3959] <= 32'b00000000010000010000000100010011;
ROM[3960] <= 32'b00000000001100010010000000100011;
ROM[3961] <= 32'b00000000010000010000000100010011;
ROM[3962] <= 32'b00000000010000010010000000100011;
ROM[3963] <= 32'b00000000010000010000000100010011;
ROM[3964] <= 32'b00000000010100010010000000100011;
ROM[3965] <= 32'b00000000010000010000000100010011;
ROM[3966] <= 32'b00000000011000010010000000100011;
ROM[3967] <= 32'b00000000010000010000000100010011;
ROM[3968] <= 32'b00000001010000000000001110010011;
ROM[3969] <= 32'b00000000100000111000001110010011;
ROM[3970] <= 32'b01000000011100010000001110110011;
ROM[3971] <= 32'b00000000011100000000001000110011;
ROM[3972] <= 32'b00000000001000000000000110110011;
ROM[3973] <= 32'b01101010100100001101000011101111;
ROM[3974] <= 32'b11111111110000010000000100010011;
ROM[3975] <= 32'b00000000000000010010001110000011;
ROM[3976] <= 32'b00000000011101100010000000100011;
ROM[3977] <= 32'b00000001110000011010001110000011;
ROM[3978] <= 32'b00000000011100010010000000100011;
ROM[3979] <= 32'b00000000010000010000000100010011;
ROM[3980] <= 32'b00000101111100000000001110010011;
ROM[3981] <= 32'b00000000011100010010000000100011;
ROM[3982] <= 32'b00000000010000010000000100010011;
ROM[3983] <= 32'b00000000000000000100001110110111;
ROM[3984] <= 32'b11101000100000111000001110010011;
ROM[3985] <= 32'b00000000111000111000001110110011;
ROM[3986] <= 32'b00000000011100010010000000100011;
ROM[3987] <= 32'b00000000010000010000000100010011;
ROM[3988] <= 32'b00000000001100010010000000100011;
ROM[3989] <= 32'b00000000010000010000000100010011;
ROM[3990] <= 32'b00000000010000010010000000100011;
ROM[3991] <= 32'b00000000010000010000000100010011;
ROM[3992] <= 32'b00000000010100010010000000100011;
ROM[3993] <= 32'b00000000010000010000000100010011;
ROM[3994] <= 32'b00000000011000010010000000100011;
ROM[3995] <= 32'b00000000010000010000000100010011;
ROM[3996] <= 32'b00000001010000000000001110010011;
ROM[3997] <= 32'b00000000100000111000001110010011;
ROM[3998] <= 32'b01000000011100010000001110110011;
ROM[3999] <= 32'b00000000011100000000001000110011;
ROM[4000] <= 32'b00000000001000000000000110110011;
ROM[4001] <= 32'b01100011100100001101000011101111;
ROM[4002] <= 32'b11111111110000010000000100010011;
ROM[4003] <= 32'b00000000000000010010001110000011;
ROM[4004] <= 32'b00000000011101100010000000100011;
ROM[4005] <= 32'b00000001110000011010001110000011;
ROM[4006] <= 32'b00000000011100010010000000100011;
ROM[4007] <= 32'b00000000010000010000000100010011;
ROM[4008] <= 32'b00000101111100000000001110010011;
ROM[4009] <= 32'b00000000011100010010000000100011;
ROM[4010] <= 32'b00000000010000010000000100010011;
ROM[4011] <= 32'b00000000000000000100001110110111;
ROM[4012] <= 32'b11101111100000111000001110010011;
ROM[4013] <= 32'b00000000111000111000001110110011;
ROM[4014] <= 32'b00000000011100010010000000100011;
ROM[4015] <= 32'b00000000010000010000000100010011;
ROM[4016] <= 32'b00000000001100010010000000100011;
ROM[4017] <= 32'b00000000010000010000000100010011;
ROM[4018] <= 32'b00000000010000010010000000100011;
ROM[4019] <= 32'b00000000010000010000000100010011;
ROM[4020] <= 32'b00000000010100010010000000100011;
ROM[4021] <= 32'b00000000010000010000000100010011;
ROM[4022] <= 32'b00000000011000010010000000100011;
ROM[4023] <= 32'b00000000010000010000000100010011;
ROM[4024] <= 32'b00000001010000000000001110010011;
ROM[4025] <= 32'b00000000100000111000001110010011;
ROM[4026] <= 32'b01000000011100010000001110110011;
ROM[4027] <= 32'b00000000011100000000001000110011;
ROM[4028] <= 32'b00000000001000000000000110110011;
ROM[4029] <= 32'b01011100100100001101000011101111;
ROM[4030] <= 32'b11111111110000010000000100010011;
ROM[4031] <= 32'b00000000000000010010001110000011;
ROM[4032] <= 32'b00000000011101100010000000100011;
ROM[4033] <= 32'b00000001110000011010001110000011;
ROM[4034] <= 32'b00000000011100010010000000100011;
ROM[4035] <= 32'b00000000010000010000000100010011;
ROM[4036] <= 32'b00000101111100000000001110010011;
ROM[4037] <= 32'b00000000011100010010000000100011;
ROM[4038] <= 32'b00000000010000010000000100010011;
ROM[4039] <= 32'b00000000000000000100001110110111;
ROM[4040] <= 32'b11110110100000111000001110010011;
ROM[4041] <= 32'b00000000111000111000001110110011;
ROM[4042] <= 32'b00000000011100010010000000100011;
ROM[4043] <= 32'b00000000010000010000000100010011;
ROM[4044] <= 32'b00000000001100010010000000100011;
ROM[4045] <= 32'b00000000010000010000000100010011;
ROM[4046] <= 32'b00000000010000010010000000100011;
ROM[4047] <= 32'b00000000010000010000000100010011;
ROM[4048] <= 32'b00000000010100010010000000100011;
ROM[4049] <= 32'b00000000010000010000000100010011;
ROM[4050] <= 32'b00000000011000010010000000100011;
ROM[4051] <= 32'b00000000010000010000000100010011;
ROM[4052] <= 32'b00000001010000000000001110010011;
ROM[4053] <= 32'b00000000100000111000001110010011;
ROM[4054] <= 32'b01000000011100010000001110110011;
ROM[4055] <= 32'b00000000011100000000001000110011;
ROM[4056] <= 32'b00000000001000000000000110110011;
ROM[4057] <= 32'b01010101100100001101000011101111;
ROM[4058] <= 32'b11111111110000010000000100010011;
ROM[4059] <= 32'b00000000000000010010001110000011;
ROM[4060] <= 32'b00000000011101100010000000100011;
ROM[4061] <= 32'b00000001110000011010001110000011;
ROM[4062] <= 32'b00000000011100010010000000100011;
ROM[4063] <= 32'b00000000010000010000000100010011;
ROM[4064] <= 32'b00000101111100000000001110010011;
ROM[4065] <= 32'b00000000011100010010000000100011;
ROM[4066] <= 32'b00000000010000010000000100010011;
ROM[4067] <= 32'b00000000000000000100001110110111;
ROM[4068] <= 32'b11111101100000111000001110010011;
ROM[4069] <= 32'b00000000111000111000001110110011;
ROM[4070] <= 32'b00000000011100010010000000100011;
ROM[4071] <= 32'b00000000010000010000000100010011;
ROM[4072] <= 32'b00000000001100010010000000100011;
ROM[4073] <= 32'b00000000010000010000000100010011;
ROM[4074] <= 32'b00000000010000010010000000100011;
ROM[4075] <= 32'b00000000010000010000000100010011;
ROM[4076] <= 32'b00000000010100010010000000100011;
ROM[4077] <= 32'b00000000010000010000000100010011;
ROM[4078] <= 32'b00000000011000010010000000100011;
ROM[4079] <= 32'b00000000010000010000000100010011;
ROM[4080] <= 32'b00000001010000000000001110010011;
ROM[4081] <= 32'b00000000100000111000001110010011;
ROM[4082] <= 32'b01000000011100010000001110110011;
ROM[4083] <= 32'b00000000011100000000001000110011;
ROM[4084] <= 32'b00000000001000000000000110110011;
ROM[4085] <= 32'b01001110100100001101000011101111;
ROM[4086] <= 32'b11111111110000010000000100010011;
ROM[4087] <= 32'b00000000000000010010001110000011;
ROM[4088] <= 32'b00000000011101100010000000100011;
ROM[4089] <= 32'b00000001110000011010001110000011;
ROM[4090] <= 32'b00000000011100011010111000100011;
ROM[4091] <= 32'b00111000000000000000000011101111;
ROM[4092] <= 32'b00000000011100000000001110010011;
ROM[4093] <= 32'b00000000011100010010000000100011;
ROM[4094] <= 32'b00000000010000010000000100010011;
ROM[4095] <= 32'b00000000000000000100001110110111;
ROM[4096] <= 32'b00000100100000111000001110010011;
ROM[4097] <= 32'b00000000111000111000001110110011;
ROM[4098] <= 32'b00000000011100010010000000100011;
ROM[4099] <= 32'b00000000010000010000000100010011;
ROM[4100] <= 32'b00000000001100010010000000100011;
ROM[4101] <= 32'b00000000010000010000000100010011;
ROM[4102] <= 32'b00000000010000010010000000100011;
ROM[4103] <= 32'b00000000010000010000000100010011;
ROM[4104] <= 32'b00000000010100010010000000100011;
ROM[4105] <= 32'b00000000010000010000000100010011;
ROM[4106] <= 32'b00000000011000010010000000100011;
ROM[4107] <= 32'b00000000010000010000000100010011;
ROM[4108] <= 32'b00000001010000000000001110010011;
ROM[4109] <= 32'b00000000010000111000001110010011;
ROM[4110] <= 32'b01000000011100010000001110110011;
ROM[4111] <= 32'b00000000011100000000001000110011;
ROM[4112] <= 32'b00000000001000000000000110110011;
ROM[4113] <= 32'b00001011110100001101000011101111;
ROM[4114] <= 32'b11111111110000010000000100010011;
ROM[4115] <= 32'b00000000000000010010001110000011;
ROM[4116] <= 32'b00000000011100011010111000100011;
ROM[4117] <= 32'b00000001110000011010001110000011;
ROM[4118] <= 32'b00000000011100010010000000100011;
ROM[4119] <= 32'b00000000010000010000000100010011;
ROM[4120] <= 32'b00000101111100000000001110010011;
ROM[4121] <= 32'b00000000011100010010000000100011;
ROM[4122] <= 32'b00000000010000010000000100010011;
ROM[4123] <= 32'b00000000000000000100001110110111;
ROM[4124] <= 32'b00001011100000111000001110010011;
ROM[4125] <= 32'b00000000111000111000001110110011;
ROM[4126] <= 32'b00000000011100010010000000100011;
ROM[4127] <= 32'b00000000010000010000000100010011;
ROM[4128] <= 32'b00000000001100010010000000100011;
ROM[4129] <= 32'b00000000010000010000000100010011;
ROM[4130] <= 32'b00000000010000010010000000100011;
ROM[4131] <= 32'b00000000010000010000000100010011;
ROM[4132] <= 32'b00000000010100010010000000100011;
ROM[4133] <= 32'b00000000010000010000000100010011;
ROM[4134] <= 32'b00000000011000010010000000100011;
ROM[4135] <= 32'b00000000010000010000000100010011;
ROM[4136] <= 32'b00000001010000000000001110010011;
ROM[4137] <= 32'b00000000100000111000001110010011;
ROM[4138] <= 32'b01000000011100010000001110110011;
ROM[4139] <= 32'b00000000011100000000001000110011;
ROM[4140] <= 32'b00000000001000000000000110110011;
ROM[4141] <= 32'b01000000100100001101000011101111;
ROM[4142] <= 32'b11111111110000010000000100010011;
ROM[4143] <= 32'b00000000000000010010001110000011;
ROM[4144] <= 32'b00000000011101100010000000100011;
ROM[4145] <= 32'b00000001110000011010001110000011;
ROM[4146] <= 32'b00000000011100010010000000100011;
ROM[4147] <= 32'b00000000010000010000000100010011;
ROM[4148] <= 32'b00000101111100000000001110010011;
ROM[4149] <= 32'b00000000011100010010000000100011;
ROM[4150] <= 32'b00000000010000010000000100010011;
ROM[4151] <= 32'b00000000000000000100001110110111;
ROM[4152] <= 32'b00010010100000111000001110010011;
ROM[4153] <= 32'b00000000111000111000001110110011;
ROM[4154] <= 32'b00000000011100010010000000100011;
ROM[4155] <= 32'b00000000010000010000000100010011;
ROM[4156] <= 32'b00000000001100010010000000100011;
ROM[4157] <= 32'b00000000010000010000000100010011;
ROM[4158] <= 32'b00000000010000010010000000100011;
ROM[4159] <= 32'b00000000010000010000000100010011;
ROM[4160] <= 32'b00000000010100010010000000100011;
ROM[4161] <= 32'b00000000010000010000000100010011;
ROM[4162] <= 32'b00000000011000010010000000100011;
ROM[4163] <= 32'b00000000010000010000000100010011;
ROM[4164] <= 32'b00000001010000000000001110010011;
ROM[4165] <= 32'b00000000100000111000001110010011;
ROM[4166] <= 32'b01000000011100010000001110110011;
ROM[4167] <= 32'b00000000011100000000001000110011;
ROM[4168] <= 32'b00000000001000000000000110110011;
ROM[4169] <= 32'b00111001100100001101000011101111;
ROM[4170] <= 32'b11111111110000010000000100010011;
ROM[4171] <= 32'b00000000000000010010001110000011;
ROM[4172] <= 32'b00000000011101100010000000100011;
ROM[4173] <= 32'b00000001110000011010001110000011;
ROM[4174] <= 32'b00000000011100010010000000100011;
ROM[4175] <= 32'b00000000010000010000000100010011;
ROM[4176] <= 32'b00000101111100000000001110010011;
ROM[4177] <= 32'b00000000011100010010000000100011;
ROM[4178] <= 32'b00000000010000010000000100010011;
ROM[4179] <= 32'b00000000000000000100001110110111;
ROM[4180] <= 32'b00011001100000111000001110010011;
ROM[4181] <= 32'b00000000111000111000001110110011;
ROM[4182] <= 32'b00000000011100010010000000100011;
ROM[4183] <= 32'b00000000010000010000000100010011;
ROM[4184] <= 32'b00000000001100010010000000100011;
ROM[4185] <= 32'b00000000010000010000000100010011;
ROM[4186] <= 32'b00000000010000010010000000100011;
ROM[4187] <= 32'b00000000010000010000000100010011;
ROM[4188] <= 32'b00000000010100010010000000100011;
ROM[4189] <= 32'b00000000010000010000000100010011;
ROM[4190] <= 32'b00000000011000010010000000100011;
ROM[4191] <= 32'b00000000010000010000000100010011;
ROM[4192] <= 32'b00000001010000000000001110010011;
ROM[4193] <= 32'b00000000100000111000001110010011;
ROM[4194] <= 32'b01000000011100010000001110110011;
ROM[4195] <= 32'b00000000011100000000001000110011;
ROM[4196] <= 32'b00000000001000000000000110110011;
ROM[4197] <= 32'b00110010100100001101000011101111;
ROM[4198] <= 32'b11111111110000010000000100010011;
ROM[4199] <= 32'b00000000000000010010001110000011;
ROM[4200] <= 32'b00000000011101100010000000100011;
ROM[4201] <= 32'b00000001110000011010001110000011;
ROM[4202] <= 32'b00000000011100010010000000100011;
ROM[4203] <= 32'b00000000010000010000000100010011;
ROM[4204] <= 32'b00000101111100000000001110010011;
ROM[4205] <= 32'b00000000011100010010000000100011;
ROM[4206] <= 32'b00000000010000010000000100010011;
ROM[4207] <= 32'b00000000000000000100001110110111;
ROM[4208] <= 32'b00100000100000111000001110010011;
ROM[4209] <= 32'b00000000111000111000001110110011;
ROM[4210] <= 32'b00000000011100010010000000100011;
ROM[4211] <= 32'b00000000010000010000000100010011;
ROM[4212] <= 32'b00000000001100010010000000100011;
ROM[4213] <= 32'b00000000010000010000000100010011;
ROM[4214] <= 32'b00000000010000010010000000100011;
ROM[4215] <= 32'b00000000010000010000000100010011;
ROM[4216] <= 32'b00000000010100010010000000100011;
ROM[4217] <= 32'b00000000010000010000000100010011;
ROM[4218] <= 32'b00000000011000010010000000100011;
ROM[4219] <= 32'b00000000010000010000000100010011;
ROM[4220] <= 32'b00000001010000000000001110010011;
ROM[4221] <= 32'b00000000100000111000001110010011;
ROM[4222] <= 32'b01000000011100010000001110110011;
ROM[4223] <= 32'b00000000011100000000001000110011;
ROM[4224] <= 32'b00000000001000000000000110110011;
ROM[4225] <= 32'b00101011100100001101000011101111;
ROM[4226] <= 32'b11111111110000010000000100010011;
ROM[4227] <= 32'b00000000000000010010001110000011;
ROM[4228] <= 32'b00000000011101100010000000100011;
ROM[4229] <= 32'b00000001110000011010001110000011;
ROM[4230] <= 32'b00000000011100010010000000100011;
ROM[4231] <= 32'b00000000010000010000000100010011;
ROM[4232] <= 32'b00000101111100000000001110010011;
ROM[4233] <= 32'b00000000011100010010000000100011;
ROM[4234] <= 32'b00000000010000010000000100010011;
ROM[4235] <= 32'b00000000000000000100001110110111;
ROM[4236] <= 32'b00100111100000111000001110010011;
ROM[4237] <= 32'b00000000111000111000001110110011;
ROM[4238] <= 32'b00000000011100010010000000100011;
ROM[4239] <= 32'b00000000010000010000000100010011;
ROM[4240] <= 32'b00000000001100010010000000100011;
ROM[4241] <= 32'b00000000010000010000000100010011;
ROM[4242] <= 32'b00000000010000010010000000100011;
ROM[4243] <= 32'b00000000010000010000000100010011;
ROM[4244] <= 32'b00000000010100010010000000100011;
ROM[4245] <= 32'b00000000010000010000000100010011;
ROM[4246] <= 32'b00000000011000010010000000100011;
ROM[4247] <= 32'b00000000010000010000000100010011;
ROM[4248] <= 32'b00000001010000000000001110010011;
ROM[4249] <= 32'b00000000100000111000001110010011;
ROM[4250] <= 32'b01000000011100010000001110110011;
ROM[4251] <= 32'b00000000011100000000001000110011;
ROM[4252] <= 32'b00000000001000000000000110110011;
ROM[4253] <= 32'b00100100100100001101000011101111;
ROM[4254] <= 32'b11111111110000010000000100010011;
ROM[4255] <= 32'b00000000000000010010001110000011;
ROM[4256] <= 32'b00000000011101100010000000100011;
ROM[4257] <= 32'b00000001110000011010001110000011;
ROM[4258] <= 32'b00000000011100010010000000100011;
ROM[4259] <= 32'b00000000010000010000000100010011;
ROM[4260] <= 32'b00000101111100000000001110010011;
ROM[4261] <= 32'b00000000011100010010000000100011;
ROM[4262] <= 32'b00000000010000010000000100010011;
ROM[4263] <= 32'b00000000000000000100001110110111;
ROM[4264] <= 32'b00101110100000111000001110010011;
ROM[4265] <= 32'b00000000111000111000001110110011;
ROM[4266] <= 32'b00000000011100010010000000100011;
ROM[4267] <= 32'b00000000010000010000000100010011;
ROM[4268] <= 32'b00000000001100010010000000100011;
ROM[4269] <= 32'b00000000010000010000000100010011;
ROM[4270] <= 32'b00000000010000010010000000100011;
ROM[4271] <= 32'b00000000010000010000000100010011;
ROM[4272] <= 32'b00000000010100010010000000100011;
ROM[4273] <= 32'b00000000010000010000000100010011;
ROM[4274] <= 32'b00000000011000010010000000100011;
ROM[4275] <= 32'b00000000010000010000000100010011;
ROM[4276] <= 32'b00000001010000000000001110010011;
ROM[4277] <= 32'b00000000100000111000001110010011;
ROM[4278] <= 32'b01000000011100010000001110110011;
ROM[4279] <= 32'b00000000011100000000001000110011;
ROM[4280] <= 32'b00000000001000000000000110110011;
ROM[4281] <= 32'b00011101100100001101000011101111;
ROM[4282] <= 32'b11111111110000010000000100010011;
ROM[4283] <= 32'b00000000000000010010001110000011;
ROM[4284] <= 32'b00000000011101100010000000100011;
ROM[4285] <= 32'b00000001110000011010001110000011;
ROM[4286] <= 32'b00000000011100010010000000100011;
ROM[4287] <= 32'b00000000010000010000000100010011;
ROM[4288] <= 32'b00000101111100000000001110010011;
ROM[4289] <= 32'b00000000011100010010000000100011;
ROM[4290] <= 32'b00000000010000010000000100010011;
ROM[4291] <= 32'b00000000000000000100001110110111;
ROM[4292] <= 32'b00110101100000111000001110010011;
ROM[4293] <= 32'b00000000111000111000001110110011;
ROM[4294] <= 32'b00000000011100010010000000100011;
ROM[4295] <= 32'b00000000010000010000000100010011;
ROM[4296] <= 32'b00000000001100010010000000100011;
ROM[4297] <= 32'b00000000010000010000000100010011;
ROM[4298] <= 32'b00000000010000010010000000100011;
ROM[4299] <= 32'b00000000010000010000000100010011;
ROM[4300] <= 32'b00000000010100010010000000100011;
ROM[4301] <= 32'b00000000010000010000000100010011;
ROM[4302] <= 32'b00000000011000010010000000100011;
ROM[4303] <= 32'b00000000010000010000000100010011;
ROM[4304] <= 32'b00000001010000000000001110010011;
ROM[4305] <= 32'b00000000100000111000001110010011;
ROM[4306] <= 32'b01000000011100010000001110110011;
ROM[4307] <= 32'b00000000011100000000001000110011;
ROM[4308] <= 32'b00000000001000000000000110110011;
ROM[4309] <= 32'b00010110100100001101000011101111;
ROM[4310] <= 32'b11111111110000010000000100010011;
ROM[4311] <= 32'b00000000000000010010001110000011;
ROM[4312] <= 32'b00000000011101100010000000100011;
ROM[4313] <= 32'b00000001110000011010001110000011;
ROM[4314] <= 32'b00000000011100011010111000100011;
ROM[4315] <= 32'b00000000000000000000001110010011;
ROM[4316] <= 32'b00000010011100011010001000100011;
ROM[4317] <= 32'b00000100010000000000001110010011;
ROM[4318] <= 32'b00000000011100010010000000100011;
ROM[4319] <= 32'b00000000010000010000000100010011;
ROM[4320] <= 32'b00000000000000000100001110110111;
ROM[4321] <= 32'b00111100110000111000001110010011;
ROM[4322] <= 32'b00000000111000111000001110110011;
ROM[4323] <= 32'b00000000011100010010000000100011;
ROM[4324] <= 32'b00000000010000010000000100010011;
ROM[4325] <= 32'b00000000001100010010000000100011;
ROM[4326] <= 32'b00000000010000010000000100010011;
ROM[4327] <= 32'b00000000010000010010000000100011;
ROM[4328] <= 32'b00000000010000010000000100010011;
ROM[4329] <= 32'b00000000010100010010000000100011;
ROM[4330] <= 32'b00000000010000010000000100010011;
ROM[4331] <= 32'b00000000011000010010000000100011;
ROM[4332] <= 32'b00000000010000010000000100010011;
ROM[4333] <= 32'b00000001010000000000001110010011;
ROM[4334] <= 32'b00000000010000111000001110010011;
ROM[4335] <= 32'b01000000011100010000001110110011;
ROM[4336] <= 32'b00000000011100000000001000110011;
ROM[4337] <= 32'b00000000001000000000000110110011;
ROM[4338] <= 32'b01010111100000001011000011101111;
ROM[4339] <= 32'b11111111110000010000000100010011;
ROM[4340] <= 32'b00000000000000010010001110000011;
ROM[4341] <= 32'b00000000011101100010000000100011;
ROM[4342] <= 32'b00000000000000000000001110010011;
ROM[4343] <= 32'b00000000011100011010101000100011;
ROM[4344] <= 32'b00000010010000011010001110000011;
ROM[4345] <= 32'b00000000011100010010000000100011;
ROM[4346] <= 32'b00000000010000010000000100010011;
ROM[4347] <= 32'b00000000000000000000001110010011;
ROM[4348] <= 32'b11111111110000010000000100010011;
ROM[4349] <= 32'b00000000000000010010010000000011;
ROM[4350] <= 32'b00000000011101000010010010110011;
ROM[4351] <= 32'b00000000100000111010010100110011;
ROM[4352] <= 32'b00000000101001001000001110110011;
ROM[4353] <= 32'b00000000000100111000001110010011;
ROM[4354] <= 32'b00000000000100111111001110010011;
ROM[4355] <= 32'b00000000000000111000101001100011;
ROM[4356] <= 32'b00000000000000000100001110110111;
ROM[4357] <= 32'b01000010010000111000001110010011;
ROM[4358] <= 32'b00000000111000111000001110110011;
ROM[4359] <= 32'b00000000000000111000000011100111;
ROM[4360] <= 32'b00000100100000000000000011101111;
ROM[4361] <= 32'b00000001100000011010001110000011;
ROM[4362] <= 32'b00000000011100010010000000100011;
ROM[4363] <= 32'b00000000010000010000000100010011;
ROM[4364] <= 32'b00000000000000000000001110010011;
ROM[4365] <= 32'b11111111110000010000000100010011;
ROM[4366] <= 32'b00000000000000010010010000000011;
ROM[4367] <= 32'b00000000100000111010001110110011;
ROM[4368] <= 32'b00000000000000111000101001100011;
ROM[4369] <= 32'b00000000000000000100001110110111;
ROM[4370] <= 32'b01000101100000111000001110010011;
ROM[4371] <= 32'b00000000111000111000001110110011;
ROM[4372] <= 32'b00000000000000111000000011100111;
ROM[4373] <= 32'b00000001000000000000000011101111;
ROM[4374] <= 32'b00000000000100000000001110010011;
ROM[4375] <= 32'b00000000011100011010101000100011;
ROM[4376] <= 32'b00000000010000000000000011101111;
ROM[4377] <= 32'b00000000010000000000000011101111;
ROM[4378] <= 32'b00000001010000011010001110000011;
ROM[4379] <= 32'b00000000011100010010000000100011;
ROM[4380] <= 32'b00000000010000010000000100010011;
ROM[4381] <= 32'b00000000000100000000001110010011;
ROM[4382] <= 32'b11111111110000010000000100010011;
ROM[4383] <= 32'b00000000000000010010010000000011;
ROM[4384] <= 32'b00000000011101000010010010110011;
ROM[4385] <= 32'b00000000100000111010010100110011;
ROM[4386] <= 32'b00000000101001001000001110110011;
ROM[4387] <= 32'b00000000000100111000001110010011;
ROM[4388] <= 32'b00000000000100111111001110010011;
ROM[4389] <= 32'b01000000011100000000001110110011;
ROM[4390] <= 32'b00000000000100111000001110010011;
ROM[4391] <= 32'b00000000000000111000101001100011;
ROM[4392] <= 32'b00000000000000000101001110110111;
ROM[4393] <= 32'b00100110110000111000001110010011;
ROM[4394] <= 32'b00000000111000111000001110110011;
ROM[4395] <= 32'b00000000000000111000000011100111;
ROM[4396] <= 32'b00000110010000011010001110000011;
ROM[4397] <= 32'b00000000011100010010000000100011;
ROM[4398] <= 32'b00000000010000010000000100010011;
ROM[4399] <= 32'b00000000000000000100001110110111;
ROM[4400] <= 32'b01010000100000111000001110010011;
ROM[4401] <= 32'b00000000111000111000001110110011;
ROM[4402] <= 32'b00000000011100010010000000100011;
ROM[4403] <= 32'b00000000010000010000000100010011;
ROM[4404] <= 32'b00000000001100010010000000100011;
ROM[4405] <= 32'b00000000010000010000000100010011;
ROM[4406] <= 32'b00000000010000010010000000100011;
ROM[4407] <= 32'b00000000010000010000000100010011;
ROM[4408] <= 32'b00000000010100010010000000100011;
ROM[4409] <= 32'b00000000010000010000000100010011;
ROM[4410] <= 32'b00000000011000010010000000100011;
ROM[4411] <= 32'b00000000010000010000000100010011;
ROM[4412] <= 32'b00000001010000000000001110010011;
ROM[4413] <= 32'b00000000010000111000001110010011;
ROM[4414] <= 32'b01000000011100010000001110110011;
ROM[4415] <= 32'b00000000011100000000001000110011;
ROM[4416] <= 32'b00000000001000000000000110110011;
ROM[4417] <= 32'b00011011000000001100000011101111;
ROM[4418] <= 32'b11111111110000010000000100010011;
ROM[4419] <= 32'b00000000000000010010001110000011;
ROM[4420] <= 32'b00000000011101100010000000100011;
ROM[4421] <= 32'b00000001110000011010001110000011;
ROM[4422] <= 32'b00000000011100010010000000100011;
ROM[4423] <= 32'b00000000010000010000000100010011;
ROM[4424] <= 32'b00000000000000000100001110110111;
ROM[4425] <= 32'b01010110110000111000001110010011;
ROM[4426] <= 32'b00000000111000111000001110110011;
ROM[4427] <= 32'b00000000011100010010000000100011;
ROM[4428] <= 32'b00000000010000010000000100010011;
ROM[4429] <= 32'b00000000001100010010000000100011;
ROM[4430] <= 32'b00000000010000010000000100010011;
ROM[4431] <= 32'b00000000010000010010000000100011;
ROM[4432] <= 32'b00000000010000010000000100010011;
ROM[4433] <= 32'b00000000010100010010000000100011;
ROM[4434] <= 32'b00000000010000010000000100010011;
ROM[4435] <= 32'b00000000011000010010000000100011;
ROM[4436] <= 32'b00000000010000010000000100010011;
ROM[4437] <= 32'b00000001010000000000001110010011;
ROM[4438] <= 32'b00000000010000111000001110010011;
ROM[4439] <= 32'b01000000011100010000001110110011;
ROM[4440] <= 32'b00000000011100000000001000110011;
ROM[4441] <= 32'b00000000001000000000000110110011;
ROM[4442] <= 32'b00010100110000001100000011101111;
ROM[4443] <= 32'b11111111110000010000000100010011;
ROM[4444] <= 32'b00000000000000010010001110000011;
ROM[4445] <= 32'b00000000011101100010000000100011;
ROM[4446] <= 32'b00000000000000000100001110110111;
ROM[4447] <= 32'b01011100010000111000001110010011;
ROM[4448] <= 32'b00000000111000111000001110110011;
ROM[4449] <= 32'b00000000011100010010000000100011;
ROM[4450] <= 32'b00000000010000010000000100010011;
ROM[4451] <= 32'b00000000001100010010000000100011;
ROM[4452] <= 32'b00000000010000010000000100010011;
ROM[4453] <= 32'b00000000010000010010000000100011;
ROM[4454] <= 32'b00000000010000010000000100010011;
ROM[4455] <= 32'b00000000010100010010000000100011;
ROM[4456] <= 32'b00000000010000010000000100010011;
ROM[4457] <= 32'b00000000011000010010000000100011;
ROM[4458] <= 32'b00000000010000010000000100010011;
ROM[4459] <= 32'b00000001010000000000001110010011;
ROM[4460] <= 32'b00000000000000111000001110010011;
ROM[4461] <= 32'b01000000011100010000001110110011;
ROM[4462] <= 32'b00000000011100000000001000110011;
ROM[4463] <= 32'b00000000001000000000000110110011;
ROM[4464] <= 32'b01001010010000001100000011101111;
ROM[4465] <= 32'b11111111110000010000000100010011;
ROM[4466] <= 32'b00000000000000010010001110000011;
ROM[4467] <= 32'b00000000011101100010000000100011;
ROM[4468] <= 32'b00000110100000011010001110000011;
ROM[4469] <= 32'b00000000011100010010000000100011;
ROM[4470] <= 32'b00000000010000010000000100010011;
ROM[4471] <= 32'b00000000000000000100001110110111;
ROM[4472] <= 32'b01100010100000111000001110010011;
ROM[4473] <= 32'b00000000111000111000001110110011;
ROM[4474] <= 32'b00000000011100010010000000100011;
ROM[4475] <= 32'b00000000010000010000000100010011;
ROM[4476] <= 32'b00000000001100010010000000100011;
ROM[4477] <= 32'b00000000010000010000000100010011;
ROM[4478] <= 32'b00000000010000010010000000100011;
ROM[4479] <= 32'b00000000010000010000000100010011;
ROM[4480] <= 32'b00000000010100010010000000100011;
ROM[4481] <= 32'b00000000010000010000000100010011;
ROM[4482] <= 32'b00000000011000010010000000100011;
ROM[4483] <= 32'b00000000010000010000000100010011;
ROM[4484] <= 32'b00000001010000000000001110010011;
ROM[4485] <= 32'b00000000010000111000001110010011;
ROM[4486] <= 32'b01000000011100010000001110110011;
ROM[4487] <= 32'b00000000011100000000001000110011;
ROM[4488] <= 32'b00000000001000000000000110110011;
ROM[4489] <= 32'b00001001000000001100000011101111;
ROM[4490] <= 32'b11111111110000010000000100010011;
ROM[4491] <= 32'b00000000000000010010001110000011;
ROM[4492] <= 32'b00000000011101100010000000100011;
ROM[4493] <= 32'b00000000000000000100001110110111;
ROM[4494] <= 32'b01101000000000111000001110010011;
ROM[4495] <= 32'b00000000111000111000001110110011;
ROM[4496] <= 32'b00000000011100010010000000100011;
ROM[4497] <= 32'b00000000010000010000000100010011;
ROM[4498] <= 32'b00000000001100010010000000100011;
ROM[4499] <= 32'b00000000010000010000000100010011;
ROM[4500] <= 32'b00000000010000010010000000100011;
ROM[4501] <= 32'b00000000010000010000000100010011;
ROM[4502] <= 32'b00000000010100010010000000100011;
ROM[4503] <= 32'b00000000010000010000000100010011;
ROM[4504] <= 32'b00000000011000010010000000100011;
ROM[4505] <= 32'b00000000010000010000000100010011;
ROM[4506] <= 32'b00000001010000000000001110010011;
ROM[4507] <= 32'b00000000000000111000001110010011;
ROM[4508] <= 32'b01000000011100010000001110110011;
ROM[4509] <= 32'b00000000011100000000001000110011;
ROM[4510] <= 32'b00000000001000000000000110110011;
ROM[4511] <= 32'b01011000100100000000000011101111;
ROM[4512] <= 32'b11111111110000010000000100010011;
ROM[4513] <= 32'b00000000000000010010001110000011;
ROM[4514] <= 32'b00000010011100011010000000100011;
ROM[4515] <= 32'b00000010100000011010001110000011;
ROM[4516] <= 32'b00000000011100010010000000100011;
ROM[4517] <= 32'b00000000010000010000000100010011;
ROM[4518] <= 32'b00000000010000000000001110010011;
ROM[4519] <= 32'b00000000011100010010000000100011;
ROM[4520] <= 32'b00000000010000010000000100010011;
ROM[4521] <= 32'b00000000000000000100001110110111;
ROM[4522] <= 32'b01101111000000111000001110010011;
ROM[4523] <= 32'b00000000111000111000001110110011;
ROM[4524] <= 32'b00000000011100010010000000100011;
ROM[4525] <= 32'b00000000010000010000000100010011;
ROM[4526] <= 32'b00000000001100010010000000100011;
ROM[4527] <= 32'b00000000010000010000000100010011;
ROM[4528] <= 32'b00000000010000010010000000100011;
ROM[4529] <= 32'b00000000010000010000000100010011;
ROM[4530] <= 32'b00000000010100010010000000100011;
ROM[4531] <= 32'b00000000010000010000000100010011;
ROM[4532] <= 32'b00000000011000010010000000100011;
ROM[4533] <= 32'b00000000010000010000000100010011;
ROM[4534] <= 32'b00000001010000000000001110010011;
ROM[4535] <= 32'b00000000100000111000001110010011;
ROM[4536] <= 32'b01000000011100010000001110110011;
ROM[4537] <= 32'b00000000011100000000001000110011;
ROM[4538] <= 32'b00000000001000000000000110110011;
ROM[4539] <= 32'b00011110100100000100000011101111;
ROM[4540] <= 32'b11111111110000010000000100010011;
ROM[4541] <= 32'b00000000000000010010001110000011;
ROM[4542] <= 32'b00000100011100011010011000100011;
ROM[4543] <= 32'b00000100110000011010001110000011;
ROM[4544] <= 32'b00000000011100010010000000100011;
ROM[4545] <= 32'b00000000010000010000000100010011;
ROM[4546] <= 32'b00000000010000011010001110000011;
ROM[4547] <= 32'b11111111110000010000000100010011;
ROM[4548] <= 32'b00000000000000010010010000000011;
ROM[4549] <= 32'b00000000011101000000001110110011;
ROM[4550] <= 32'b00000000011100010010000000100011;
ROM[4551] <= 32'b00000000010000010000000100010011;
ROM[4552] <= 32'b00000000000100000000001110010011;
ROM[4553] <= 32'b00000000011101100010000000100011;
ROM[4554] <= 32'b11111111110000010000000100010011;
ROM[4555] <= 32'b00000000000000010010001110000011;
ROM[4556] <= 32'b00000000000000111000001100010011;
ROM[4557] <= 32'b00000000000001100010001110000011;
ROM[4558] <= 32'b00000000110100110000010000110011;
ROM[4559] <= 32'b00000000011101000010000000100011;
ROM[4560] <= 32'b00000000000000000000001110010011;
ROM[4561] <= 32'b00000010011100011010101000100011;
ROM[4562] <= 32'b00000000000000000000001110010011;
ROM[4563] <= 32'b00000000011100011010011000100011;
ROM[4564] <= 32'b00000000110000011010001110000011;
ROM[4565] <= 32'b00000000011100010010000000100011;
ROM[4566] <= 32'b00000000010000010000000100010011;
ROM[4567] <= 32'b00000001000000011010001110000011;
ROM[4568] <= 32'b11111111110000010000000100010011;
ROM[4569] <= 32'b00000000000000010010010000000011;
ROM[4570] <= 32'b00000000011101000010001110110011;
ROM[4571] <= 32'b01000000011100000000001110110011;
ROM[4572] <= 32'b00000000000100111000001110010011;
ROM[4573] <= 32'b00000000000000111000101001100011;
ROM[4574] <= 32'b00000000000000000101001110110111;
ROM[4575] <= 32'b10011000010000111000001110010011;
ROM[4576] <= 32'b00000000111000111000001110110011;
ROM[4577] <= 32'b00000000000000111000000011100111;
ROM[4578] <= 32'b00000000100000011010001110000011;
ROM[4579] <= 32'b00000000011100010010000000100011;
ROM[4580] <= 32'b00000000010000010000000100010011;
ROM[4581] <= 32'b00000000010000000000001110010011;
ROM[4582] <= 32'b00000000011100010010000000100011;
ROM[4583] <= 32'b00000000010000010000000100010011;
ROM[4584] <= 32'b00000000000000000100001110110111;
ROM[4585] <= 32'b01111110110000111000001110010011;
ROM[4586] <= 32'b00000000111000111000001110110011;
ROM[4587] <= 32'b00000000011100010010000000100011;
ROM[4588] <= 32'b00000000010000010000000100010011;
ROM[4589] <= 32'b00000000001100010010000000100011;
ROM[4590] <= 32'b00000000010000010000000100010011;
ROM[4591] <= 32'b00000000010000010010000000100011;
ROM[4592] <= 32'b00000000010000010000000100010011;
ROM[4593] <= 32'b00000000010100010010000000100011;
ROM[4594] <= 32'b00000000010000010000000100010011;
ROM[4595] <= 32'b00000000011000010010000000100011;
ROM[4596] <= 32'b00000000010000010000000100010011;
ROM[4597] <= 32'b00000001010000000000001110010011;
ROM[4598] <= 32'b00000000100000111000001110010011;
ROM[4599] <= 32'b01000000011100010000001110110011;
ROM[4600] <= 32'b00000000011100000000001000110011;
ROM[4601] <= 32'b00000000001000000000000110110011;
ROM[4602] <= 32'b00001110110100000100000011101111;
ROM[4603] <= 32'b11111111110000010000000100010011;
ROM[4604] <= 32'b00000000000000010010001110000011;
ROM[4605] <= 32'b00000100011100011010010000100011;
ROM[4606] <= 32'b00000100100000011010001110000011;
ROM[4607] <= 32'b00000000011100010010000000100011;
ROM[4608] <= 32'b00000000010000010000000100010011;
ROM[4609] <= 32'b00000000000000011010001110000011;
ROM[4610] <= 32'b11111111110000010000000100010011;
ROM[4611] <= 32'b00000000000000010010010000000011;
ROM[4612] <= 32'b00000000011101000000001110110011;
ROM[4613] <= 32'b00000000000000111000001100010011;
ROM[4614] <= 32'b00000000110100110000010000110011;
ROM[4615] <= 32'b00000000000001000010001110000011;
ROM[4616] <= 32'b00000010011100011010111000100011;
ROM[4617] <= 32'b00000011110000011010001110000011;
ROM[4618] <= 32'b00000000011100010010000000100011;
ROM[4619] <= 32'b00000000010000010000000100010011;
ROM[4620] <= 32'b00000000110000011010001110000011;
ROM[4621] <= 32'b00000000011100010010000000100011;
ROM[4622] <= 32'b00000000010000010000000100010011;
ROM[4623] <= 32'b00000000000000000101001110110111;
ROM[4624] <= 32'b10001000100000111000001110010011;
ROM[4625] <= 32'b00000000111000111000001110110011;
ROM[4626] <= 32'b00000000011100010010000000100011;
ROM[4627] <= 32'b00000000010000010000000100010011;
ROM[4628] <= 32'b00000000001100010010000000100011;
ROM[4629] <= 32'b00000000010000010000000100010011;
ROM[4630] <= 32'b00000000010000010010000000100011;
ROM[4631] <= 32'b00000000010000010000000100010011;
ROM[4632] <= 32'b00000000010100010010000000100011;
ROM[4633] <= 32'b00000000010000010000000100010011;
ROM[4634] <= 32'b00000000011000010010000000100011;
ROM[4635] <= 32'b00000000010000010000000100010011;
ROM[4636] <= 32'b00000001010000000000001110010011;
ROM[4637] <= 32'b00000000100000111000001110010011;
ROM[4638] <= 32'b01000000011100010000001110110011;
ROM[4639] <= 32'b00000000011100000000001000110011;
ROM[4640] <= 32'b00000000001000000000000110110011;
ROM[4641] <= 32'b00100100000000001101000011101111;
ROM[4642] <= 32'b11111111110000010000000100010011;
ROM[4643] <= 32'b00000000000000010010001110000011;
ROM[4644] <= 32'b00000010011100011010011000100011;
ROM[4645] <= 32'b00000010110000011010001110000011;
ROM[4646] <= 32'b00000000011100010010000000100011;
ROM[4647] <= 32'b00000000010000010000000100010011;
ROM[4648] <= 32'b00000010000000011010001110000011;
ROM[4649] <= 32'b11111111110000010000000100010011;
ROM[4650] <= 32'b00000000000000010010010000000011;
ROM[4651] <= 32'b00000000011101000010010010110011;
ROM[4652] <= 32'b00000000100000111010010100110011;
ROM[4653] <= 32'b00000000101001001000001110110011;
ROM[4654] <= 32'b00000000000100111000001110010011;
ROM[4655] <= 32'b00000000000100111111001110010011;
ROM[4656] <= 32'b00000000000000111000101001100011;
ROM[4657] <= 32'b00000000000000000101001110110111;
ROM[4658] <= 32'b10001101100000111000001110010011;
ROM[4659] <= 32'b00000000111000111000001110110011;
ROM[4660] <= 32'b00000000000000111000000011100111;
ROM[4661] <= 32'b00001000110000000000000011101111;
ROM[4662] <= 32'b00000000000100000000001110010011;
ROM[4663] <= 32'b00000010011100011010101000100011;
ROM[4664] <= 32'b00000001110000011010001110000011;
ROM[4665] <= 32'b00000000011100010010000000100011;
ROM[4666] <= 32'b00000000010000010000000100010011;
ROM[4667] <= 32'b00000000110000011010001110000011;
ROM[4668] <= 32'b00000000011100010010000000100011;
ROM[4669] <= 32'b00000000010000010000000100010011;
ROM[4670] <= 32'b00000010000000011010001110000011;
ROM[4671] <= 32'b00000000011100010010000000100011;
ROM[4672] <= 32'b00000000010000010000000100010011;
ROM[4673] <= 32'b00000000000000000101001110110111;
ROM[4674] <= 32'b10010101000000111000001110010011;
ROM[4675] <= 32'b00000000111000111000001110110011;
ROM[4676] <= 32'b00000000011100010010000000100011;
ROM[4677] <= 32'b00000000010000010000000100010011;
ROM[4678] <= 32'b00000000001100010010000000100011;
ROM[4679] <= 32'b00000000010000010000000100010011;
ROM[4680] <= 32'b00000000010000010010000000100011;
ROM[4681] <= 32'b00000000010000010000000100010011;
ROM[4682] <= 32'b00000000010100010010000000100011;
ROM[4683] <= 32'b00000000010000010000000100010011;
ROM[4684] <= 32'b00000000011000010010000000100011;
ROM[4685] <= 32'b00000000010000010000000100010011;
ROM[4686] <= 32'b00000001010000000000001110010011;
ROM[4687] <= 32'b00000000110000111000001110010011;
ROM[4688] <= 32'b01000000011100010000001110110011;
ROM[4689] <= 32'b00000000011100000000001000110011;
ROM[4690] <= 32'b00000000001000000000000110110011;
ROM[4691] <= 32'b00100110010000001101000011101111;
ROM[4692] <= 32'b11111111110000010000000100010011;
ROM[4693] <= 32'b00000000000000010010001110000011;
ROM[4694] <= 32'b00000000011101100010000000100011;
ROM[4695] <= 32'b00000000010000000000000011101111;
ROM[4696] <= 32'b00000000110000011010001110000011;
ROM[4697] <= 32'b00000000011100010010000000100011;
ROM[4698] <= 32'b00000000010000010000000100010011;
ROM[4699] <= 32'b00000000000100000000001110010011;
ROM[4700] <= 32'b11111111110000010000000100010011;
ROM[4701] <= 32'b00000000000000010010010000000011;
ROM[4702] <= 32'b00000000011101000000001110110011;
ROM[4703] <= 32'b00000000011100011010011000100011;
ROM[4704] <= 32'b11011101000111111111000011101111;
ROM[4705] <= 32'b00000011010000011010001110000011;
ROM[4706] <= 32'b00000000011100010010000000100011;
ROM[4707] <= 32'b00000000010000010000000100010011;
ROM[4708] <= 32'b00000000000000000000001110010011;
ROM[4709] <= 32'b11111111110000010000000100010011;
ROM[4710] <= 32'b00000000000000010010010000000011;
ROM[4711] <= 32'b00000000011101000010010010110011;
ROM[4712] <= 32'b00000000100000111010010100110011;
ROM[4713] <= 32'b00000000101001001000001110110011;
ROM[4714] <= 32'b00000000000100111000001110010011;
ROM[4715] <= 32'b00000000000100111111001110010011;
ROM[4716] <= 32'b00000000000000111000101001100011;
ROM[4717] <= 32'b00000000000000000101001110110111;
ROM[4718] <= 32'b10011100100000111000001110010011;
ROM[4719] <= 32'b00000000111000111000001110110011;
ROM[4720] <= 32'b00000000000000111000000011100111;
ROM[4721] <= 32'b01000110010000000000000011101111;
ROM[4722] <= 32'b00000001100000011010001110000011;
ROM[4723] <= 32'b00000000011100010010000000100011;
ROM[4724] <= 32'b00000000010000010000000100010011;
ROM[4725] <= 32'b00000000000100000000001110010011;
ROM[4726] <= 32'b11111111110000010000000100010011;
ROM[4727] <= 32'b00000000000000010010010000000011;
ROM[4728] <= 32'b00000000011101000010010010110011;
ROM[4729] <= 32'b00000000100000111010010100110011;
ROM[4730] <= 32'b00000000101001001000001110110011;
ROM[4731] <= 32'b00000000000100111000001110010011;
ROM[4732] <= 32'b00000000000100111111001110010011;
ROM[4733] <= 32'b00000000000000111000101001100011;
ROM[4734] <= 32'b00000000000000000101001110110111;
ROM[4735] <= 32'b10100000110000111000001110010011;
ROM[4736] <= 32'b00000000111000111000001110110011;
ROM[4737] <= 32'b00000000000000111000000011100111;
ROM[4738] <= 32'b00100111100000000000000011101111;
ROM[4739] <= 32'b00000110110000011010001110000011;
ROM[4740] <= 32'b00000000011100010010000000100011;
ROM[4741] <= 32'b00000000010000010000000100010011;
ROM[4742] <= 32'b00000000000000000101001110110111;
ROM[4743] <= 32'b10100110010000111000001110010011;
ROM[4744] <= 32'b00000000111000111000001110110011;
ROM[4745] <= 32'b00000000011100010010000000100011;
ROM[4746] <= 32'b00000000010000010000000100010011;
ROM[4747] <= 32'b00000000001100010010000000100011;
ROM[4748] <= 32'b00000000010000010000000100010011;
ROM[4749] <= 32'b00000000010000010010000000100011;
ROM[4750] <= 32'b00000000010000010000000100010011;
ROM[4751] <= 32'b00000000010100010010000000100011;
ROM[4752] <= 32'b00000000010000010000000100010011;
ROM[4753] <= 32'b00000000011000010010000000100011;
ROM[4754] <= 32'b00000000010000010000000100010011;
ROM[4755] <= 32'b00000001010000000000001110010011;
ROM[4756] <= 32'b00000000010000111000001110010011;
ROM[4757] <= 32'b01000000011100010000001110110011;
ROM[4758] <= 32'b00000000011100000000001000110011;
ROM[4759] <= 32'b00000000001000000000000110110011;
ROM[4760] <= 32'b01000101010100001011000011101111;
ROM[4761] <= 32'b11111111110000010000000100010011;
ROM[4762] <= 32'b00000000000000010010001110000011;
ROM[4763] <= 32'b00000000011101100010000000100011;
ROM[4764] <= 32'b00000000000000000101001110110111;
ROM[4765] <= 32'b10101011110000111000001110010011;
ROM[4766] <= 32'b00000000111000111000001110110011;
ROM[4767] <= 32'b00000000011100010010000000100011;
ROM[4768] <= 32'b00000000010000010000000100010011;
ROM[4769] <= 32'b00000000001100010010000000100011;
ROM[4770] <= 32'b00000000010000010000000100010011;
ROM[4771] <= 32'b00000000010000010010000000100011;
ROM[4772] <= 32'b00000000010000010000000100010011;
ROM[4773] <= 32'b00000000010100010010000000100011;
ROM[4774] <= 32'b00000000010000010000000100010011;
ROM[4775] <= 32'b00000000011000010010000000100011;
ROM[4776] <= 32'b00000000010000010000000100010011;
ROM[4777] <= 32'b00000001010000000000001110010011;
ROM[4778] <= 32'b00000000000000111000001110010011;
ROM[4779] <= 32'b01000000011100010000001110110011;
ROM[4780] <= 32'b00000000011100000000001000110011;
ROM[4781] <= 32'b00000000001000000000000110110011;
ROM[4782] <= 32'b01111010110100001011000011101111;
ROM[4783] <= 32'b11111111110000010000000100010011;
ROM[4784] <= 32'b00000000000000010010001110000011;
ROM[4785] <= 32'b00000000011101100010000000100011;
ROM[4786] <= 32'b00000111000000011010001110000011;
ROM[4787] <= 32'b00000000011100010010000000100011;
ROM[4788] <= 32'b00000000010000010000000100010011;
ROM[4789] <= 32'b00000000000000000101001110110111;
ROM[4790] <= 32'b10110010000000111000001110010011;
ROM[4791] <= 32'b00000000111000111000001110110011;
ROM[4792] <= 32'b00000000011100010010000000100011;
ROM[4793] <= 32'b00000000010000010000000100010011;
ROM[4794] <= 32'b00000000001100010010000000100011;
ROM[4795] <= 32'b00000000010000010000000100010011;
ROM[4796] <= 32'b00000000010000010010000000100011;
ROM[4797] <= 32'b00000000010000010000000100010011;
ROM[4798] <= 32'b00000000010100010010000000100011;
ROM[4799] <= 32'b00000000010000010000000100010011;
ROM[4800] <= 32'b00000000011000010010000000100011;
ROM[4801] <= 32'b00000000010000010000000100010011;
ROM[4802] <= 32'b00000001010000000000001110010011;
ROM[4803] <= 32'b00000000010000111000001110010011;
ROM[4804] <= 32'b01000000011100010000001110110011;
ROM[4805] <= 32'b00000000011100000000001000110011;
ROM[4806] <= 32'b00000000001000000000000110110011;
ROM[4807] <= 32'b00111001100100001011000011101111;
ROM[4808] <= 32'b11111111110000010000000100010011;
ROM[4809] <= 32'b00000000000000010010001110000011;
ROM[4810] <= 32'b00000000011101100010000000100011;
ROM[4811] <= 32'b00000000100000011010001110000011;
ROM[4812] <= 32'b00000000011100010010000000100011;
ROM[4813] <= 32'b00000000010000010000000100010011;
ROM[4814] <= 32'b00000000010000000000001110010011;
ROM[4815] <= 32'b00000000011100010010000000100011;
ROM[4816] <= 32'b00000000010000010000000100010011;
ROM[4817] <= 32'b00000000000000000101001110110111;
ROM[4818] <= 32'b10111001000000111000001110010011;
ROM[4819] <= 32'b00000000111000111000001110110011;
ROM[4820] <= 32'b00000000011100010010000000100011;
ROM[4821] <= 32'b00000000010000010000000100010011;
ROM[4822] <= 32'b00000000001100010010000000100011;
ROM[4823] <= 32'b00000000010000010000000100010011;
ROM[4824] <= 32'b00000000010000010010000000100011;
ROM[4825] <= 32'b00000000010000010000000100010011;
ROM[4826] <= 32'b00000000010100010010000000100011;
ROM[4827] <= 32'b00000000010000010000000100010011;
ROM[4828] <= 32'b00000000011000010010000000100011;
ROM[4829] <= 32'b00000000010000010000000100010011;
ROM[4830] <= 32'b00000001010000000000001110010011;
ROM[4831] <= 32'b00000000100000111000001110010011;
ROM[4832] <= 32'b01000000011100010000001110110011;
ROM[4833] <= 32'b00000000011100000000001000110011;
ROM[4834] <= 32'b00000000001000000000000110110011;
ROM[4835] <= 32'b01010100100000000100000011101111;
ROM[4836] <= 32'b11111111110000010000000100010011;
ROM[4837] <= 32'b00000000000000010010001110000011;
ROM[4838] <= 32'b00000100011100011010010000100011;
ROM[4839] <= 32'b00000100100000011010001110000011;
ROM[4840] <= 32'b00000000011100010010000000100011;
ROM[4841] <= 32'b00000000010000010000000100010011;
ROM[4842] <= 32'b00000000000000011010001110000011;
ROM[4843] <= 32'b11111111110000010000000100010011;
ROM[4844] <= 32'b00000000000000010010010000000011;
ROM[4845] <= 32'b00000000011101000000001110110011;
ROM[4846] <= 32'b00000000000000111000001100010011;
ROM[4847] <= 32'b00000000110100110000010000110011;
ROM[4848] <= 32'b00000000000001000010001110000011;
ROM[4849] <= 32'b00000000011100010010000000100011;
ROM[4850] <= 32'b00000000010000010000000100010011;
ROM[4851] <= 32'b00000000000000000101001110110111;
ROM[4852] <= 32'b11000001100000111000001110010011;
ROM[4853] <= 32'b00000000111000111000001110110011;
ROM[4854] <= 32'b00000000011100010010000000100011;
ROM[4855] <= 32'b00000000010000010000000100010011;
ROM[4856] <= 32'b00000000001100010010000000100011;
ROM[4857] <= 32'b00000000010000010000000100010011;
ROM[4858] <= 32'b00000000010000010010000000100011;
ROM[4859] <= 32'b00000000010000010000000100010011;
ROM[4860] <= 32'b00000000010100010010000000100011;
ROM[4861] <= 32'b00000000010000010000000100010011;
ROM[4862] <= 32'b00000000011000010010000000100011;
ROM[4863] <= 32'b00000000010000010000000100010011;
ROM[4864] <= 32'b00000001010000000000001110010011;
ROM[4865] <= 32'b00000000010000111000001110010011;
ROM[4866] <= 32'b01000000011100010000001110110011;
ROM[4867] <= 32'b00000000011100000000001000110011;
ROM[4868] <= 32'b00000000001000000000000110110011;
ROM[4869] <= 32'b00101010000100001011000011101111;
ROM[4870] <= 32'b11111111110000010000000100010011;
ROM[4871] <= 32'b00000000000000010010001110000011;
ROM[4872] <= 32'b00000000011101100010000000100011;
ROM[4873] <= 32'b00000000000000000101001110110111;
ROM[4874] <= 32'b11000111000000111000001110010011;
ROM[4875] <= 32'b00000000111000111000001110110011;
ROM[4876] <= 32'b00000000011100010010000000100011;
ROM[4877] <= 32'b00000000010000010000000100010011;
ROM[4878] <= 32'b00000000001100010010000000100011;
ROM[4879] <= 32'b00000000010000010000000100010011;
ROM[4880] <= 32'b00000000010000010010000000100011;
ROM[4881] <= 32'b00000000010000010000000100010011;
ROM[4882] <= 32'b00000000010100010010000000100011;
ROM[4883] <= 32'b00000000010000010000000100010011;
ROM[4884] <= 32'b00000000011000010010000000100011;
ROM[4885] <= 32'b00000000010000010000000100010011;
ROM[4886] <= 32'b00000001010000000000001110010011;
ROM[4887] <= 32'b00000000000000111000001110010011;
ROM[4888] <= 32'b01000000011100010000001110110011;
ROM[4889] <= 32'b00000000011100000000001000110011;
ROM[4890] <= 32'b00000000001000000000000110110011;
ROM[4891] <= 32'b01011111100100001011000011101111;
ROM[4892] <= 32'b11111111110000010000000100010011;
ROM[4893] <= 32'b00000000000000010010001110000011;
ROM[4894] <= 32'b00000000011101100010000000100011;
ROM[4895] <= 32'b00011000100000000000000011101111;
ROM[4896] <= 32'b00000110110000011010001110000011;
ROM[4897] <= 32'b00000000011100010010000000100011;
ROM[4898] <= 32'b00000000010000010000000100010011;
ROM[4899] <= 32'b00000000000000000101001110110111;
ROM[4900] <= 32'b11001101100000111000001110010011;
ROM[4901] <= 32'b00000000111000111000001110110011;
ROM[4902] <= 32'b00000000011100010010000000100011;
ROM[4903] <= 32'b00000000010000010000000100010011;
ROM[4904] <= 32'b00000000001100010010000000100011;
ROM[4905] <= 32'b00000000010000010000000100010011;
ROM[4906] <= 32'b00000000010000010010000000100011;
ROM[4907] <= 32'b00000000010000010000000100010011;
ROM[4908] <= 32'b00000000010100010010000000100011;
ROM[4909] <= 32'b00000000010000010000000100010011;
ROM[4910] <= 32'b00000000011000010010000000100011;
ROM[4911] <= 32'b00000000010000010000000100010011;
ROM[4912] <= 32'b00000001010000000000001110010011;
ROM[4913] <= 32'b00000000010000111000001110010011;
ROM[4914] <= 32'b01000000011100010000001110110011;
ROM[4915] <= 32'b00000000011100000000001000110011;
ROM[4916] <= 32'b00000000001000000000000110110011;
ROM[4917] <= 32'b00011110000100001011000011101111;
ROM[4918] <= 32'b11111111110000010000000100010011;
ROM[4919] <= 32'b00000000000000010010001110000011;
ROM[4920] <= 32'b00000000011101100010000000100011;
ROM[4921] <= 32'b00000001100000011010001110000011;
ROM[4922] <= 32'b00000000011100010010000000100011;
ROM[4923] <= 32'b00000000010000010000000100010011;
ROM[4924] <= 32'b00000000000000000101001110110111;
ROM[4925] <= 32'b11010011110000111000001110010011;
ROM[4926] <= 32'b00000000111000111000001110110011;
ROM[4927] <= 32'b00000000011100010010000000100011;
ROM[4928] <= 32'b00000000010000010000000100010011;
ROM[4929] <= 32'b00000000001100010010000000100011;
ROM[4930] <= 32'b00000000010000010000000100010011;
ROM[4931] <= 32'b00000000010000010010000000100011;
ROM[4932] <= 32'b00000000010000010000000100010011;
ROM[4933] <= 32'b00000000010100010010000000100011;
ROM[4934] <= 32'b00000000010000010000000100010011;
ROM[4935] <= 32'b00000000011000010010000000100011;
ROM[4936] <= 32'b00000000010000010000000100010011;
ROM[4937] <= 32'b00000001010000000000001110010011;
ROM[4938] <= 32'b00000000010000111000001110010011;
ROM[4939] <= 32'b01000000011100010000001110110011;
ROM[4940] <= 32'b00000000011100000000001000110011;
ROM[4941] <= 32'b00000000001000000000000110110011;
ROM[4942] <= 32'b00110100010100001011000011101111;
ROM[4943] <= 32'b11111111110000010000000100010011;
ROM[4944] <= 32'b00000000000000010010001110000011;
ROM[4945] <= 32'b00000000011101100010000000100011;
ROM[4946] <= 32'b00000001100000011010001110000011;
ROM[4947] <= 32'b00000000011100010010000000100011;
ROM[4948] <= 32'b00000000010000010000000100010011;
ROM[4949] <= 32'b00000000000000000101001110110111;
ROM[4950] <= 32'b11011010000000111000001110010011;
ROM[4951] <= 32'b00000000111000111000001110110011;
ROM[4952] <= 32'b00000000011100010010000000100011;
ROM[4953] <= 32'b00000000010000010000000100010011;
ROM[4954] <= 32'b00000000001100010010000000100011;
ROM[4955] <= 32'b00000000010000010000000100010011;
ROM[4956] <= 32'b00000000010000010010000000100011;
ROM[4957] <= 32'b00000000010000010000000100010011;
ROM[4958] <= 32'b00000000010100010010000000100011;
ROM[4959] <= 32'b00000000010000010000000100010011;
ROM[4960] <= 32'b00000000011000010010000000100011;
ROM[4961] <= 32'b00000000010000010000000100010011;
ROM[4962] <= 32'b00000001010000000000001110010011;
ROM[4963] <= 32'b00000000010000111000001110010011;
ROM[4964] <= 32'b01000000011100010000001110110011;
ROM[4965] <= 32'b00000000011100000000001000110011;
ROM[4966] <= 32'b00000000001000000000000110110011;
ROM[4967] <= 32'b00010001100100001011000011101111;
ROM[4968] <= 32'b11111111110000010000000100010011;
ROM[4969] <= 32'b00000000000000010010001110000011;
ROM[4970] <= 32'b00000000011101100010000000100011;
ROM[4971] <= 32'b00000000000000000101001110110111;
ROM[4972] <= 32'b11011111100000111000001110010011;
ROM[4973] <= 32'b00000000111000111000001110110011;
ROM[4974] <= 32'b00000000011100010010000000100011;
ROM[4975] <= 32'b00000000010000010000000100010011;
ROM[4976] <= 32'b00000000001100010010000000100011;
ROM[4977] <= 32'b00000000010000010000000100010011;
ROM[4978] <= 32'b00000000010000010010000000100011;
ROM[4979] <= 32'b00000000010000010000000100010011;
ROM[4980] <= 32'b00000000010100010010000000100011;
ROM[4981] <= 32'b00000000010000010000000100010011;
ROM[4982] <= 32'b00000000011000010010000000100011;
ROM[4983] <= 32'b00000000010000010000000100010011;
ROM[4984] <= 32'b00000001010000000000001110010011;
ROM[4985] <= 32'b00000000000000111000001110010011;
ROM[4986] <= 32'b01000000011100010000001110110011;
ROM[4987] <= 32'b00000000011100000000001000110011;
ROM[4988] <= 32'b00000000001000000000000110110011;
ROM[4989] <= 32'b01000111000100001011000011101111;
ROM[4990] <= 32'b11111111110000010000000100010011;
ROM[4991] <= 32'b00000000000000010010001110000011;
ROM[4992] <= 32'b00000000011101100010000000100011;
ROM[4993] <= 32'b00000001100000011010001110000011;
ROM[4994] <= 32'b00000000011100010010000000100011;
ROM[4995] <= 32'b00000000010000010000000100010011;
ROM[4996] <= 32'b00000000000100000000001110010011;
ROM[4997] <= 32'b11111111110000010000000100010011;
ROM[4998] <= 32'b00000000000000010010010000000011;
ROM[4999] <= 32'b01000000011101000000001110110011;
ROM[5000] <= 32'b00000000011100011010110000100011;
ROM[5001] <= 32'b00110101110000000000000011101111;
ROM[5002] <= 32'b00000000000000000000001110010011;
ROM[5003] <= 32'b00000010011100011010110000100011;
ROM[5004] <= 32'b00000000000000000000001110010011;
ROM[5005] <= 32'b00000000011100011010011000100011;
ROM[5006] <= 32'b00000000110000011010001110000011;
ROM[5007] <= 32'b00000000011100010010000000100011;
ROM[5008] <= 32'b00000000010000010000000100010011;
ROM[5009] <= 32'b00000001000000011010001110000011;
ROM[5010] <= 32'b11111111110000010000000100010011;
ROM[5011] <= 32'b00000000000000010010010000000011;
ROM[5012] <= 32'b00000000011101000010001110110011;
ROM[5013] <= 32'b01000000011100000000001110110011;
ROM[5014] <= 32'b00000000000100111000001110010011;
ROM[5015] <= 32'b00000000000000111000101001100011;
ROM[5016] <= 32'b00000000000000000101001110110111;
ROM[5017] <= 32'b11110101010000111000001110010011;
ROM[5018] <= 32'b00000000111000111000001110110011;
ROM[5019] <= 32'b00000000000000111000000011100111;
ROM[5020] <= 32'b00000001110000011010001110000011;
ROM[5021] <= 32'b00000000011100010010000000100011;
ROM[5022] <= 32'b00000000010000010000000100010011;
ROM[5023] <= 32'b00000000110000011010001110000011;
ROM[5024] <= 32'b00000000011100010010000000100011;
ROM[5025] <= 32'b00000000010000010000000100010011;
ROM[5026] <= 32'b00000000000000000101001110110111;
ROM[5027] <= 32'b11101101010000111000001110010011;
ROM[5028] <= 32'b00000000111000111000001110110011;
ROM[5029] <= 32'b00000000011100010010000000100011;
ROM[5030] <= 32'b00000000010000010000000100010011;
ROM[5031] <= 32'b00000000001100010010000000100011;
ROM[5032] <= 32'b00000000010000010000000100010011;
ROM[5033] <= 32'b00000000010000010010000000100011;
ROM[5034] <= 32'b00000000010000010000000100010011;
ROM[5035] <= 32'b00000000010100010010000000100011;
ROM[5036] <= 32'b00000000010000010000000100010011;
ROM[5037] <= 32'b00000000011000010010000000100011;
ROM[5038] <= 32'b00000000010000010000000100010011;
ROM[5039] <= 32'b00000001010000000000001110010011;
ROM[5040] <= 32'b00000000100000111000001110010011;
ROM[5041] <= 32'b01000000011100010000001110110011;
ROM[5042] <= 32'b00000000011100000000001000110011;
ROM[5043] <= 32'b00000000001000000000000110110011;
ROM[5044] <= 32'b00111111010100001100000011101111;
ROM[5045] <= 32'b11111111110000010000000100010011;
ROM[5046] <= 32'b00000000000000010010001110000011;
ROM[5047] <= 32'b00000010011100011010011000100011;
ROM[5048] <= 32'b00000010110000011010001110000011;
ROM[5049] <= 32'b00000000011100010010000000100011;
ROM[5050] <= 32'b00000000010000010000000100010011;
ROM[5051] <= 32'b00000011000000011010001110000011;
ROM[5052] <= 32'b11111111110000010000000100010011;
ROM[5053] <= 32'b00000000000000010010010000000011;
ROM[5054] <= 32'b00000000011101000010010010110011;
ROM[5055] <= 32'b00000000100000111010010100110011;
ROM[5056] <= 32'b00000000101001001000001110110011;
ROM[5057] <= 32'b00000000000100111000001110010011;
ROM[5058] <= 32'b00000000000100111111001110010011;
ROM[5059] <= 32'b00000000000000111000101001100011;
ROM[5060] <= 32'b00000000000000000101001110110111;
ROM[5061] <= 32'b11110010010000111000001110010011;
ROM[5062] <= 32'b00000000111000111000001110110011;
ROM[5063] <= 32'b00000000000000111000000011100111;
ROM[5064] <= 32'b00000001000000000000000011101111;
ROM[5065] <= 32'b00000000000100000000001110010011;
ROM[5066] <= 32'b00000010011100011010110000100011;
ROM[5067] <= 32'b00000000010000000000000011101111;
ROM[5068] <= 32'b00000000110000011010001110000011;
ROM[5069] <= 32'b00000000011100010010000000100011;
ROM[5070] <= 32'b00000000010000010000000100010011;
ROM[5071] <= 32'b00000000000100000000001110010011;
ROM[5072] <= 32'b11111111110000010000000100010011;
ROM[5073] <= 32'b00000000000000010010010000000011;
ROM[5074] <= 32'b00000000011101000000001110110011;
ROM[5075] <= 32'b00000000011100011010011000100011;
ROM[5076] <= 32'b11101110100111111111000011101111;
ROM[5077] <= 32'b00000011100000011010001110000011;
ROM[5078] <= 32'b00000000011100010010000000100011;
ROM[5079] <= 32'b00000000010000010000000100010011;
ROM[5080] <= 32'b00000000000000000000001110010011;
ROM[5081] <= 32'b11111111110000010000000100010011;
ROM[5082] <= 32'b00000000000000010010010000000011;
ROM[5083] <= 32'b00000000011101000010010010110011;
ROM[5084] <= 32'b00000000100000111010010100110011;
ROM[5085] <= 32'b00000000101001001000001110110011;
ROM[5086] <= 32'b00000000000100111000001110010011;
ROM[5087] <= 32'b00000000000100111111001110010011;
ROM[5088] <= 32'b00000000000000111000101001100011;
ROM[5089] <= 32'b00000000000000000101001110110111;
ROM[5090] <= 32'b11111001100000111000001110010011;
ROM[5091] <= 32'b00000000111000111000001110110011;
ROM[5092] <= 32'b00000000000000111000000011100111;
ROM[5093] <= 32'b00011110110000000000000011101111;
ROM[5094] <= 32'b00000000000100000000001110010011;
ROM[5095] <= 32'b00000010011100011010001000100011;
ROM[5096] <= 32'b00000111010000011010001110000011;
ROM[5097] <= 32'b00000000011100010010000000100011;
ROM[5098] <= 32'b00000000010000010000000100010011;
ROM[5099] <= 32'b00000000000000000101001110110111;
ROM[5100] <= 32'b11111111100000111000001110010011;
ROM[5101] <= 32'b00000000111000111000001110110011;
ROM[5102] <= 32'b00000000011100010010000000100011;
ROM[5103] <= 32'b00000000010000010000000100010011;
ROM[5104] <= 32'b00000000001100010010000000100011;
ROM[5105] <= 32'b00000000010000010000000100010011;
ROM[5106] <= 32'b00000000010000010010000000100011;
ROM[5107] <= 32'b00000000010000010000000100010011;
ROM[5108] <= 32'b00000000010100010010000000100011;
ROM[5109] <= 32'b00000000010000010000000100010011;
ROM[5110] <= 32'b00000000011000010010000000100011;
ROM[5111] <= 32'b00000000010000010000000100010011;
ROM[5112] <= 32'b00000001010000000000001110010011;
ROM[5113] <= 32'b00000000010000111000001110010011;
ROM[5114] <= 32'b01000000011100010000001110110011;
ROM[5115] <= 32'b00000000011100000000001000110011;
ROM[5116] <= 32'b00000000001000000000000110110011;
ROM[5117] <= 32'b01101100000000001011000011101111;
ROM[5118] <= 32'b11111111110000010000000100010011;
ROM[5119] <= 32'b00000000000000010010001110000011;
ROM[5120] <= 32'b00000000011101100010000000100011;
ROM[5121] <= 32'b00000000000000000101001110110111;
ROM[5122] <= 32'b00000101000000111000001110010011;
ROM[5123] <= 32'b00000000111000111000001110110011;
ROM[5124] <= 32'b00000000011100010010000000100011;
ROM[5125] <= 32'b00000000010000010000000100010011;
ROM[5126] <= 32'b00000000001100010010000000100011;
ROM[5127] <= 32'b00000000010000010000000100010011;
ROM[5128] <= 32'b00000000010000010010000000100011;
ROM[5129] <= 32'b00000000010000010000000100010011;
ROM[5130] <= 32'b00000000010100010010000000100011;
ROM[5131] <= 32'b00000000010000010000000100010011;
ROM[5132] <= 32'b00000000011000010010000000100011;
ROM[5133] <= 32'b00000000010000010000000100010011;
ROM[5134] <= 32'b00000001010000000000001110010011;
ROM[5135] <= 32'b00000000000000111000001110010011;
ROM[5136] <= 32'b01000000011100010000001110110011;
ROM[5137] <= 32'b00000000011100000000001000110011;
ROM[5138] <= 32'b00000000001000000000000110110011;
ROM[5139] <= 32'b00100001100100001011000011101111;
ROM[5140] <= 32'b11111111110000010000000100010011;
ROM[5141] <= 32'b00000000000000010010001110000011;
ROM[5142] <= 32'b00000000011101100010000000100011;
ROM[5143] <= 32'b00000111000000011010001110000011;
ROM[5144] <= 32'b00000000011100010010000000100011;
ROM[5145] <= 32'b00000000010000010000000100010011;
ROM[5146] <= 32'b00000000000000000101001110110111;
ROM[5147] <= 32'b00001011010000111000001110010011;
ROM[5148] <= 32'b00000000111000111000001110110011;
ROM[5149] <= 32'b00000000011100010010000000100011;
ROM[5150] <= 32'b00000000010000010000000100010011;
ROM[5151] <= 32'b00000000001100010010000000100011;
ROM[5152] <= 32'b00000000010000010000000100010011;
ROM[5153] <= 32'b00000000010000010010000000100011;
ROM[5154] <= 32'b00000000010000010000000100010011;
ROM[5155] <= 32'b00000000010100010010000000100011;
ROM[5156] <= 32'b00000000010000010000000100010011;
ROM[5157] <= 32'b00000000011000010010000000100011;
ROM[5158] <= 32'b00000000010000010000000100010011;
ROM[5159] <= 32'b00000001010000000000001110010011;
ROM[5160] <= 32'b00000000010000111000001110010011;
ROM[5161] <= 32'b01000000011100010000001110110011;
ROM[5162] <= 32'b00000000011100000000001000110011;
ROM[5163] <= 32'b00000000001000000000000110110011;
ROM[5164] <= 32'b01100000010000001011000011101111;
ROM[5165] <= 32'b11111111110000010000000100010011;
ROM[5166] <= 32'b00000000000000010010001110000011;
ROM[5167] <= 32'b00000000011101100010000000100011;
ROM[5168] <= 32'b00000001110000011010001110000011;
ROM[5169] <= 32'b00000000011100010010000000100011;
ROM[5170] <= 32'b00000000010000010000000100010011;
ROM[5171] <= 32'b00000000000000000101001110110111;
ROM[5172] <= 32'b00010001100000111000001110010011;
ROM[5173] <= 32'b00000000111000111000001110110011;
ROM[5174] <= 32'b00000000011100010010000000100011;
ROM[5175] <= 32'b00000000010000010000000100010011;
ROM[5176] <= 32'b00000000001100010010000000100011;
ROM[5177] <= 32'b00000000010000010000000100010011;
ROM[5178] <= 32'b00000000010000010010000000100011;
ROM[5179] <= 32'b00000000010000010000000100010011;
ROM[5180] <= 32'b00000000010100010010000000100011;
ROM[5181] <= 32'b00000000010000010000000100010011;
ROM[5182] <= 32'b00000000011000010010000000100011;
ROM[5183] <= 32'b00000000010000010000000100010011;
ROM[5184] <= 32'b00000001010000000000001110010011;
ROM[5185] <= 32'b00000000010000111000001110010011;
ROM[5186] <= 32'b01000000011100010000001110110011;
ROM[5187] <= 32'b00000000011100000000001000110011;
ROM[5188] <= 32'b00000000001000000000000110110011;
ROM[5189] <= 32'b01011010000000001011000011101111;
ROM[5190] <= 32'b11111111110000010000000100010011;
ROM[5191] <= 32'b00000000000000010010001110000011;
ROM[5192] <= 32'b00000000011101100010000000100011;
ROM[5193] <= 32'b00000000000000000101001110110111;
ROM[5194] <= 32'b00010111000000111000001110010011;
ROM[5195] <= 32'b00000000111000111000001110110011;
ROM[5196] <= 32'b00000000011100010010000000100011;
ROM[5197] <= 32'b00000000010000010000000100010011;
ROM[5198] <= 32'b00000000001100010010000000100011;
ROM[5199] <= 32'b00000000010000010000000100010011;
ROM[5200] <= 32'b00000000010000010010000000100011;
ROM[5201] <= 32'b00000000010000010000000100010011;
ROM[5202] <= 32'b00000000010100010010000000100011;
ROM[5203] <= 32'b00000000010000010000000100010011;
ROM[5204] <= 32'b00000000011000010010000000100011;
ROM[5205] <= 32'b00000000010000010000000100010011;
ROM[5206] <= 32'b00000001010000000000001110010011;
ROM[5207] <= 32'b00000000000000111000001110010011;
ROM[5208] <= 32'b01000000011100010000001110110011;
ROM[5209] <= 32'b00000000011100000000001000110011;
ROM[5210] <= 32'b00000000001000000000000110110011;
ROM[5211] <= 32'b00001111100100001011000011101111;
ROM[5212] <= 32'b11111111110000010000000100010011;
ROM[5213] <= 32'b00000000000000010010001110000011;
ROM[5214] <= 32'b00000000011101100010000000100011;
ROM[5215] <= 32'b00000000010000000000000011101111;
ROM[5216] <= 32'b00000000000000000000001110010011;
ROM[5217] <= 32'b00000000011100011010101000100011;
ROM[5218] <= 32'b00000010010000011010001110000011;
ROM[5219] <= 32'b00000000011100010010000000100011;
ROM[5220] <= 32'b00000000010000010000000100010011;
ROM[5221] <= 32'b00000000000000000000001110010011;
ROM[5222] <= 32'b11111111110000010000000100010011;
ROM[5223] <= 32'b00000000000000010010010000000011;
ROM[5224] <= 32'b00000000011101000010010010110011;
ROM[5225] <= 32'b00000000100000111010010100110011;
ROM[5226] <= 32'b00000000101001001000001110110011;
ROM[5227] <= 32'b00000000000100111000001110010011;
ROM[5228] <= 32'b00000000000100111111001110010011;
ROM[5229] <= 32'b00000000000000111000101001100011;
ROM[5230] <= 32'b00000000000000000101001110110111;
ROM[5231] <= 32'b00011100110000111000001110010011;
ROM[5232] <= 32'b00000000111000111000001110110011;
ROM[5233] <= 32'b00000000000000111000000011100111;
ROM[5234] <= 32'b00000100100000000000000011101111;
ROM[5235] <= 32'b00000001100000011010001110000011;
ROM[5236] <= 32'b00000000011100010010000000100011;
ROM[5237] <= 32'b00000000010000010000000100010011;
ROM[5238] <= 32'b00000000000000000000001110010011;
ROM[5239] <= 32'b11111111110000010000000100010011;
ROM[5240] <= 32'b00000000000000010010010000000011;
ROM[5241] <= 32'b00000000100000111010001110110011;
ROM[5242] <= 32'b00000000000000111000101001100011;
ROM[5243] <= 32'b00000000000000000101001110110111;
ROM[5244] <= 32'b00100000000000111000001110010011;
ROM[5245] <= 32'b00000000111000111000001110110011;
ROM[5246] <= 32'b00000000000000111000000011100111;
ROM[5247] <= 32'b00000001000000000000000011101111;
ROM[5248] <= 32'b00000000000100000000001110010011;
ROM[5249] <= 32'b00000000011100011010101000100011;
ROM[5250] <= 32'b00000000010000000000000011101111;
ROM[5251] <= 32'b00000000010000000000000011101111;
ROM[5252] <= 32'b00000000000000000101001110110111;
ROM[5253] <= 32'b00100101110000111000001110010011;
ROM[5254] <= 32'b00000000111000111000001110110011;
ROM[5255] <= 32'b00000000011100010010000000100011;
ROM[5256] <= 32'b00000000010000010000000100010011;
ROM[5257] <= 32'b00000000001100010010000000100011;
ROM[5258] <= 32'b00000000010000010000000100010011;
ROM[5259] <= 32'b00000000010000010010000000100011;
ROM[5260] <= 32'b00000000010000010000000100010011;
ROM[5261] <= 32'b00000000010100010010000000100011;
ROM[5262] <= 32'b00000000010000010000000100010011;
ROM[5263] <= 32'b00000000011000010010000000100011;
ROM[5264] <= 32'b00000000010000010000000100010011;
ROM[5265] <= 32'b00000001010000000000001110010011;
ROM[5266] <= 32'b00000000000000111000001110010011;
ROM[5267] <= 32'b01000000011100010000001110110011;
ROM[5268] <= 32'b00000000011100000000001000110011;
ROM[5269] <= 32'b00000000001000000000000110110011;
ROM[5270] <= 32'b00000000110100001011000011101111;
ROM[5271] <= 32'b11111111110000010000000100010011;
ROM[5272] <= 32'b00000000000000010010001110000011;
ROM[5273] <= 32'b00000000011101100010000000100011;
ROM[5274] <= 32'b10100000000011111111000011101111;
ROM[5275] <= 32'b00000000100000011010001110000011;
ROM[5276] <= 32'b00000000011100010010000000100011;
ROM[5277] <= 32'b00000000010000010000000100010011;
ROM[5278] <= 32'b00000000000100000000001110010011;
ROM[5279] <= 32'b11111111110000010000000100010011;
ROM[5280] <= 32'b00000000000000010010010000000011;
ROM[5281] <= 32'b00000000011101000000001110110011;
ROM[5282] <= 32'b00000000011100011010010000100011;
ROM[5283] <= 32'b10101010110111111101000011101111;
ROM[5284] <= 32'b00000000000000000000001110010011;
ROM[5285] <= 32'b00000000011100010010000000100011;
ROM[5286] <= 32'b00000000010000010000000100010011;
ROM[5287] <= 32'b00000001010000000000001110010011;
ROM[5288] <= 32'b01000000011100011000001110110011;
ROM[5289] <= 32'b00000000000000111010000010000011;
ROM[5290] <= 32'b11111111110000010000000100010011;
ROM[5291] <= 32'b00000000000000010010001110000011;
ROM[5292] <= 32'b00000000011100100010000000100011;
ROM[5293] <= 32'b00000000010000100000000100010011;
ROM[5294] <= 32'b00000001010000000000001110010011;
ROM[5295] <= 32'b01000000011100011000001110110011;
ROM[5296] <= 32'b00000000010000111010000110000011;
ROM[5297] <= 32'b00000000100000111010001000000011;
ROM[5298] <= 32'b00000000110000111010001010000011;
ROM[5299] <= 32'b00000001000000111010001100000011;
ROM[5300] <= 32'b00000000000000001000000011100111;
ROM[5301] <= 32'b00000000000000000100001110110111;
ROM[5302] <= 32'b11111111111100111000001110010011;
ROM[5303] <= 32'b00000100011101101010000000100011;
ROM[5304] <= 32'b00000100000001101010001110000011;
ROM[5305] <= 32'b00000000011100010010000000100011;
ROM[5306] <= 32'b00000000010000010000000100010011;
ROM[5307] <= 32'b00000000010000000000001110010011;
ROM[5308] <= 32'b00000000011100010010000000100011;
ROM[5309] <= 32'b00000000010000010000000100010011;
ROM[5310] <= 32'b00000000000000000101001110110111;
ROM[5311] <= 32'b00110100010000111000001110010011;
ROM[5312] <= 32'b00000000111000111000001110110011;
ROM[5313] <= 32'b00000000011100010010000000100011;
ROM[5314] <= 32'b00000000010000010000000100010011;
ROM[5315] <= 32'b00000000001100010010000000100011;
ROM[5316] <= 32'b00000000010000010000000100010011;
ROM[5317] <= 32'b00000000010000010010000000100011;
ROM[5318] <= 32'b00000000010000010000000100010011;
ROM[5319] <= 32'b00000000010100010010000000100011;
ROM[5320] <= 32'b00000000010000010000000100010011;
ROM[5321] <= 32'b00000000011000010010000000100011;
ROM[5322] <= 32'b00000000010000010000000100010011;
ROM[5323] <= 32'b00000001010000000000001110010011;
ROM[5324] <= 32'b00000000100000111000001110010011;
ROM[5325] <= 32'b01000000011100010000001110110011;
ROM[5326] <= 32'b00000000011100000000001000110011;
ROM[5327] <= 32'b00000000001000000000000110110011;
ROM[5328] <= 32'b01011001010100000011000011101111;
ROM[5329] <= 32'b11111111110000010000000100010011;
ROM[5330] <= 32'b00000000000000010010001110000011;
ROM[5331] <= 32'b00000100011101101010000000100011;
ROM[5332] <= 32'b00000000000000000000001110010011;
ROM[5333] <= 32'b00000100011101101010001000100011;
ROM[5334] <= 32'b00000000000000000000001110010011;
ROM[5335] <= 32'b00000000011100010010000000100011;
ROM[5336] <= 32'b00000000010000010000000100010011;
ROM[5337] <= 32'b00000001010000000000001110010011;
ROM[5338] <= 32'b01000000011100011000001110110011;
ROM[5339] <= 32'b00000000000000111010000010000011;
ROM[5340] <= 32'b11111111110000010000000100010011;
ROM[5341] <= 32'b00000000000000010010001110000011;
ROM[5342] <= 32'b00000000011100100010000000100011;
ROM[5343] <= 32'b00000000010000100000000100010011;
ROM[5344] <= 32'b00000001010000000000001110010011;
ROM[5345] <= 32'b01000000011100011000001110110011;
ROM[5346] <= 32'b00000000010000111010000110000011;
ROM[5347] <= 32'b00000000100000111010001000000011;
ROM[5348] <= 32'b00000000110000111010001010000011;
ROM[5349] <= 32'b00000001000000111010001100000011;
ROM[5350] <= 32'b00000000000000001000000011100111;
ROM[5351] <= 32'b00000000000000000000001110010011;
ROM[5352] <= 32'b00000000011100010010000000100011;
ROM[5353] <= 32'b00000000010000010000000100010011;
ROM[5354] <= 32'b00000100000001101010001110000011;
ROM[5355] <= 32'b11111111110000010000000100010011;
ROM[5356] <= 32'b00000000000000010010010000000011;
ROM[5357] <= 32'b00000000011101000000001110110011;
ROM[5358] <= 32'b00000000000000111000001100010011;
ROM[5359] <= 32'b00000000110100110000010000110011;
ROM[5360] <= 32'b00000000000001000010001110000011;
ROM[5361] <= 32'b00000000011100010010000000100011;
ROM[5362] <= 32'b00000000010000010000000100010011;
ROM[5363] <= 32'b00000001010000000000001110010011;
ROM[5364] <= 32'b01000000011100011000001110110011;
ROM[5365] <= 32'b00000000000000111010000010000011;
ROM[5366] <= 32'b11111111110000010000000100010011;
ROM[5367] <= 32'b00000000000000010010001110000011;
ROM[5368] <= 32'b00000000011100100010000000100011;
ROM[5369] <= 32'b00000000010000100000000100010011;
ROM[5370] <= 32'b00000001010000000000001110010011;
ROM[5371] <= 32'b01000000011100011000001110110011;
ROM[5372] <= 32'b00000000010000111010000110000011;
ROM[5373] <= 32'b00000000100000111010001000000011;
ROM[5374] <= 32'b00000000110000111010001010000011;
ROM[5375] <= 32'b00000001000000111010001100000011;
ROM[5376] <= 32'b00000000000000001000000011100111;
ROM[5377] <= 32'b00000000000000010010000000100011;
ROM[5378] <= 32'b00000000010000010000000100010011;
ROM[5379] <= 32'b00000000000000010010000000100011;
ROM[5380] <= 32'b00000000010000010000000100010011;
ROM[5381] <= 32'b00000000000000000000001110010011;
ROM[5382] <= 32'b00000000011100011010001000100011;
ROM[5383] <= 32'b00000000010000011010001110000011;
ROM[5384] <= 32'b00000000011100010010000000100011;
ROM[5385] <= 32'b00000000010000010000000100010011;
ROM[5386] <= 32'b00000000000000000000001110010011;
ROM[5387] <= 32'b11111111110000010000000100010011;
ROM[5388] <= 32'b00000000000000010010010000000011;
ROM[5389] <= 32'b00000000011101000010010010110011;
ROM[5390] <= 32'b00000000100000111010010100110011;
ROM[5391] <= 32'b00000000101001001000001110110011;
ROM[5392] <= 32'b00000000000100111000001110010011;
ROM[5393] <= 32'b00000000000100111111001110010011;
ROM[5394] <= 32'b01000000011100000000001110110011;
ROM[5395] <= 32'b00000000000100111000001110010011;
ROM[5396] <= 32'b00000000000000111000101001100011;
ROM[5397] <= 32'b00000000000000000101001110110111;
ROM[5398] <= 32'b01011011000000111000001110010011;
ROM[5399] <= 32'b00000000111000111000001110110011;
ROM[5400] <= 32'b00000000000000111000000011100111;
ROM[5401] <= 32'b00000000000000000101001110110111;
ROM[5402] <= 32'b01001011000000111000001110010011;
ROM[5403] <= 32'b00000000111000111000001110110011;
ROM[5404] <= 32'b00000000011100010010000000100011;
ROM[5405] <= 32'b00000000010000010000000100010011;
ROM[5406] <= 32'b00000000001100010010000000100011;
ROM[5407] <= 32'b00000000010000010000000100010011;
ROM[5408] <= 32'b00000000010000010010000000100011;
ROM[5409] <= 32'b00000000010000010000000100010011;
ROM[5410] <= 32'b00000000010100010010000000100011;
ROM[5411] <= 32'b00000000010000010000000100010011;
ROM[5412] <= 32'b00000000011000010010000000100011;
ROM[5413] <= 32'b00000000010000010000000100010011;
ROM[5414] <= 32'b00000001010000000000001110010011;
ROM[5415] <= 32'b00000000000000111000001110010011;
ROM[5416] <= 32'b01000000011100010000001110110011;
ROM[5417] <= 32'b00000000011100000000001000110011;
ROM[5418] <= 32'b00000000001000000000000110110011;
ROM[5419] <= 32'b11101111000111111111000011101111;
ROM[5420] <= 32'b11111111110000010000000100010011;
ROM[5421] <= 32'b00000000000000010010001110000011;
ROM[5422] <= 32'b00000000011100011010000000100011;
ROM[5423] <= 32'b00000000000000011010001110000011;
ROM[5424] <= 32'b00000000011100010010000000100011;
ROM[5425] <= 32'b00000000010000010000000100010011;
ROM[5426] <= 32'b00000000100100000000001110010011;
ROM[5427] <= 32'b11111111110000010000000100010011;
ROM[5428] <= 32'b00000000000000010010010000000011;
ROM[5429] <= 32'b00000000011101000010010010110011;
ROM[5430] <= 32'b00000000100000111010010100110011;
ROM[5431] <= 32'b00000000101001001000001110110011;
ROM[5432] <= 32'b00000000000100111000001110010011;
ROM[5433] <= 32'b00000000000100111111001110010011;
ROM[5434] <= 32'b00000000000000111000101001100011;
ROM[5435] <= 32'b00000000000000000101001110110111;
ROM[5436] <= 32'b01010000000000111000001110010011;
ROM[5437] <= 32'b00000000111000111000001110110011;
ROM[5438] <= 32'b00000000000000111000000011100111;
ROM[5439] <= 32'b00000110000000000000000011101111;
ROM[5440] <= 32'b00000100010001101010001110000011;
ROM[5441] <= 32'b00000000011100010010000000100011;
ROM[5442] <= 32'b00000000010000010000000100010011;
ROM[5443] <= 32'b00000000000000000000001110010011;
ROM[5444] <= 32'b11111111110000010000000100010011;
ROM[5445] <= 32'b00000000000000010010010000000011;
ROM[5446] <= 32'b00000000011101000010010010110011;
ROM[5447] <= 32'b00000000100000111010010100110011;
ROM[5448] <= 32'b00000000101001001000001110110011;
ROM[5449] <= 32'b00000000000100111000001110010011;
ROM[5450] <= 32'b00000000000100111111001110010011;
ROM[5451] <= 32'b00000000000000111000101001100011;
ROM[5452] <= 32'b00000000000000000101001110110111;
ROM[5453] <= 32'b01010100010000111000001110010011;
ROM[5454] <= 32'b00000000111000111000001110110011;
ROM[5455] <= 32'b00000000000000111000000011100111;
ROM[5456] <= 32'b00000001000000000000000011101111;
ROM[5457] <= 32'b00000010000000000000001110010011;
ROM[5458] <= 32'b00000100011101101010001000100011;
ROM[5459] <= 32'b00000000110000000000000011101111;
ROM[5460] <= 32'b00000000000000000000001110010011;
ROM[5461] <= 32'b00000100011101101010001000100011;
ROM[5462] <= 32'b00000101010000000000000011101111;
ROM[5463] <= 32'b00000000000000011010001110000011;
ROM[5464] <= 32'b00000000011100010010000000100011;
ROM[5465] <= 32'b00000000010000010000000100010011;
ROM[5466] <= 32'b00000000000000000000001110010011;
ROM[5467] <= 32'b11111111110000010000000100010011;
ROM[5468] <= 32'b00000000000000010010010000000011;
ROM[5469] <= 32'b00000000011101000010010010110011;
ROM[5470] <= 32'b00000000100000111010010100110011;
ROM[5471] <= 32'b00000000101001001000001110110011;
ROM[5472] <= 32'b00000000000100111000001110010011;
ROM[5473] <= 32'b00000000000100111111001110010011;
ROM[5474] <= 32'b00000000000000111000101001100011;
ROM[5475] <= 32'b00000000000000000101001110110111;
ROM[5476] <= 32'b01011010000000111000001110010011;
ROM[5477] <= 32'b00000000111000111000001110110011;
ROM[5478] <= 32'b00000000000000111000000011100111;
ROM[5479] <= 32'b00000000100000000000000011101111;
ROM[5480] <= 32'b00000000110000000000000011101111;
ROM[5481] <= 32'b00000000000100000000001110010011;
ROM[5482] <= 32'b00000000011100011010001000100011;
ROM[5483] <= 32'b11100111000111111111000011101111;
ROM[5484] <= 32'b00000000000000011010001110000011;
ROM[5485] <= 32'b00000000011100010010000000100011;
ROM[5486] <= 32'b00000000010000010000000100010011;
ROM[5487] <= 32'b00000110000000000000001110010011;
ROM[5488] <= 32'b11111111110000010000000100010011;
ROM[5489] <= 32'b00000000000000010010010000000011;
ROM[5490] <= 32'b00000000100000111010001110110011;
ROM[5491] <= 32'b00000000000000111000101001100011;
ROM[5492] <= 32'b00000000000000000101001110110111;
ROM[5493] <= 32'b01011110010000111000001110010011;
ROM[5494] <= 32'b00000000111000111000001110110011;
ROM[5495] <= 32'b00000000000000111000000011100111;
ROM[5496] <= 32'b00001100010000000000000011101111;
ROM[5497] <= 32'b00000000000000011010001110000011;
ROM[5498] <= 32'b00000000011100010010000000100011;
ROM[5499] <= 32'b00000000010000010000000100010011;
ROM[5500] <= 32'b00000111101100000000001110010011;
ROM[5501] <= 32'b11111111110000010000000100010011;
ROM[5502] <= 32'b00000000000000010010010000000011;
ROM[5503] <= 32'b00000000011101000010001110110011;
ROM[5504] <= 32'b00000000000000111000101001100011;
ROM[5505] <= 32'b00000000000000000101001110110111;
ROM[5506] <= 32'b01100001100000111000001110010011;
ROM[5507] <= 32'b00000000111000111000001110110011;
ROM[5508] <= 32'b00000000000000111000000011100111;
ROM[5509] <= 32'b00001000110000000000000011101111;
ROM[5510] <= 32'b00000000000000011010001110000011;
ROM[5511] <= 32'b00000000011100010010000000100011;
ROM[5512] <= 32'b00000000010000010000000100010011;
ROM[5513] <= 32'b00000100010001101010001110000011;
ROM[5514] <= 32'b11111111110000010000000100010011;
ROM[5515] <= 32'b00000000000000010010010000000011;
ROM[5516] <= 32'b01000000011101000000001110110011;
ROM[5517] <= 32'b00000000011100011010000000100011;
ROM[5518] <= 32'b00000000000000011010001110000011;
ROM[5519] <= 32'b00000000011100010010000000100011;
ROM[5520] <= 32'b00000000010000010000000100010011;
ROM[5521] <= 32'b00000000000000000101001110110111;
ROM[5522] <= 32'b01101001000000111000001110010011;
ROM[5523] <= 32'b00000000111000111000001110110011;
ROM[5524] <= 32'b00000000011100010010000000100011;
ROM[5525] <= 32'b00000000010000010000000100010011;
ROM[5526] <= 32'b00000000001100010010000000100011;
ROM[5527] <= 32'b00000000010000010000000100010011;
ROM[5528] <= 32'b00000000010000010010000000100011;
ROM[5529] <= 32'b00000000010000010000000100010011;
ROM[5530] <= 32'b00000000010100010010000000100011;
ROM[5531] <= 32'b00000000010000010000000100010011;
ROM[5532] <= 32'b00000000011000010010000000100011;
ROM[5533] <= 32'b00000000010000010000000100010011;
ROM[5534] <= 32'b00000001010000000000001110010011;
ROM[5535] <= 32'b00000000010000111000001110010011;
ROM[5536] <= 32'b01000000011100010000001110110011;
ROM[5537] <= 32'b00000000011100000000001000110011;
ROM[5538] <= 32'b00000000001000000000000110110011;
ROM[5539] <= 32'b00101011010000001010000011101111;
ROM[5540] <= 32'b11111111110000010000000100010011;
ROM[5541] <= 32'b00000000000000010010001110000011;
ROM[5542] <= 32'b00000000011101100010000000100011;
ROM[5543] <= 32'b00000000010000000000000011101111;
ROM[5544] <= 32'b00000000010000000000000011101111;
ROM[5545] <= 32'b00000000000000011010001110000011;
ROM[5546] <= 32'b00000000011100010010000000100011;
ROM[5547] <= 32'b00000000010000010000000100010011;
ROM[5548] <= 32'b00000010111100000000001110010011;
ROM[5549] <= 32'b11111111110000010000000100010011;
ROM[5550] <= 32'b00000000000000010010010000000011;
ROM[5551] <= 32'b00000000100000111010001110110011;
ROM[5552] <= 32'b00000000000000111000101001100011;
ROM[5553] <= 32'b00000000000000000101001110110111;
ROM[5554] <= 32'b01101101100000111000001110010011;
ROM[5555] <= 32'b00000000111000111000001110110011;
ROM[5556] <= 32'b00000000000000111000000011100111;
ROM[5557] <= 32'b00001010010000000000000011101111;
ROM[5558] <= 32'b00000000000000011010001110000011;
ROM[5559] <= 32'b00000000011100010010000000100011;
ROM[5560] <= 32'b00000000010000010000000100010011;
ROM[5561] <= 32'b00000011101000000000001110010011;
ROM[5562] <= 32'b11111111110000010000000100010011;
ROM[5563] <= 32'b00000000000000010010010000000011;
ROM[5564] <= 32'b00000000011101000010001110110011;
ROM[5565] <= 32'b00000000000000111000101001100011;
ROM[5566] <= 32'b00000000000000000101001110110111;
ROM[5567] <= 32'b01110000110000111000001110010011;
ROM[5568] <= 32'b00000000111000111000001110110011;
ROM[5569] <= 32'b00000000000000111000000011100111;
ROM[5570] <= 32'b00000110110000000000000011101111;
ROM[5571] <= 32'b00000000000000011010001110000011;
ROM[5572] <= 32'b00000000011100010010000000100011;
ROM[5573] <= 32'b00000000010000010000000100010011;
ROM[5574] <= 32'b00000000000000000101001110110111;
ROM[5575] <= 32'b01110110010000111000001110010011;
ROM[5576] <= 32'b00000000111000111000001110110011;
ROM[5577] <= 32'b00000000011100010010000000100011;
ROM[5578] <= 32'b00000000010000010000000100010011;
ROM[5579] <= 32'b00000000001100010010000000100011;
ROM[5580] <= 32'b00000000010000010000000100010011;
ROM[5581] <= 32'b00000000010000010010000000100011;
ROM[5582] <= 32'b00000000010000010000000100010011;
ROM[5583] <= 32'b00000000010100010010000000100011;
ROM[5584] <= 32'b00000000010000010000000100010011;
ROM[5585] <= 32'b00000000011000010010000000100011;
ROM[5586] <= 32'b00000000010000010000000100010011;
ROM[5587] <= 32'b00000001010000000000001110010011;
ROM[5588] <= 32'b00000000010000111000001110010011;
ROM[5589] <= 32'b01000000011100010000001110110011;
ROM[5590] <= 32'b00000000011100000000001000110011;
ROM[5591] <= 32'b00000000001000000000000110110011;
ROM[5592] <= 32'b00011110000000001010000011101111;
ROM[5593] <= 32'b11111111110000010000000100010011;
ROM[5594] <= 32'b00000000000000010010001110000011;
ROM[5595] <= 32'b00000000011101100010000000100011;
ROM[5596] <= 32'b00000000010000000000000011101111;
ROM[5597] <= 32'b00000000010000000000000011101111;
ROM[5598] <= 32'b00000000000000011010001110000011;
ROM[5599] <= 32'b00000000011100010010000000100011;
ROM[5600] <= 32'b00000000010000010000000100010011;
ROM[5601] <= 32'b00000001010000000000001110010011;
ROM[5602] <= 32'b01000000011100011000001110110011;
ROM[5603] <= 32'b00000000000000111010000010000011;
ROM[5604] <= 32'b11111111110000010000000100010011;
ROM[5605] <= 32'b00000000000000010010001110000011;
ROM[5606] <= 32'b00000000011100100010000000100011;
ROM[5607] <= 32'b00000000010000100000000100010011;
ROM[5608] <= 32'b00000001010000000000001110010011;
ROM[5609] <= 32'b01000000011100011000001110110011;
ROM[5610] <= 32'b00000000010000111010000110000011;
ROM[5611] <= 32'b00000000100000111010001000000011;
ROM[5612] <= 32'b00000000110000111010001010000011;
ROM[5613] <= 32'b00000001000000111010001100000011;
ROM[5614] <= 32'b00000000000000001000000011100111;
ROM[5615] <= 32'b00000000000000010010000000100011;
ROM[5616] <= 32'b00000000010000010000000100010011;
ROM[5617] <= 32'b00000000000000010010000000100011;
ROM[5618] <= 32'b00000000010000010000000100010011;
ROM[5619] <= 32'b00000000000000100010001110000011;
ROM[5620] <= 32'b00000000011100010010000000100011;
ROM[5621] <= 32'b00000000010000010000000100010011;
ROM[5622] <= 32'b00000000000000000110001110110111;
ROM[5623] <= 32'b10000010010000111000001110010011;
ROM[5624] <= 32'b00000000111000111000001110110011;
ROM[5625] <= 32'b00000000011100010010000000100011;
ROM[5626] <= 32'b00000000010000010000000100010011;
ROM[5627] <= 32'b00000000001100010010000000100011;
ROM[5628] <= 32'b00000000010000010000000100010011;
ROM[5629] <= 32'b00000000010000010010000000100011;
ROM[5630] <= 32'b00000000010000010000000100010011;
ROM[5631] <= 32'b00000000010100010010000000100011;
ROM[5632] <= 32'b00000000010000010000000100010011;
ROM[5633] <= 32'b00000000011000010010000000100011;
ROM[5634] <= 32'b00000000010000010000000100010011;
ROM[5635] <= 32'b00000001010000000000001110010011;
ROM[5636] <= 32'b00000000010000111000001110010011;
ROM[5637] <= 32'b01000000011100010000001110110011;
ROM[5638] <= 32'b00000000011100000000001000110011;
ROM[5639] <= 32'b00000000001000000000000110110011;
ROM[5640] <= 32'b01101001010100001010000011101111;
ROM[5641] <= 32'b11111111110000010000000100010011;
ROM[5642] <= 32'b00000000000000010010001110000011;
ROM[5643] <= 32'b00000000011101100010000000100011;
ROM[5644] <= 32'b00000011001000000000001110010011;
ROM[5645] <= 32'b00000000011100010010000000100011;
ROM[5646] <= 32'b00000000010000010000000100010011;
ROM[5647] <= 32'b00000000000000000110001110110111;
ROM[5648] <= 32'b10001000100000111000001110010011;
ROM[5649] <= 32'b00000000111000111000001110110011;
ROM[5650] <= 32'b00000000011100010010000000100011;
ROM[5651] <= 32'b00000000010000010000000100010011;
ROM[5652] <= 32'b00000000001100010010000000100011;
ROM[5653] <= 32'b00000000010000010000000100010011;
ROM[5654] <= 32'b00000000010000010010000000100011;
ROM[5655] <= 32'b00000000010000010000000100010011;
ROM[5656] <= 32'b00000000010100010010000000100011;
ROM[5657] <= 32'b00000000010000010000000100010011;
ROM[5658] <= 32'b00000000011000010010000000100011;
ROM[5659] <= 32'b00000000010000010000000100010011;
ROM[5660] <= 32'b00000001010000000000001110010011;
ROM[5661] <= 32'b00000000010000111000001110010011;
ROM[5662] <= 32'b01000000011100010000001110110011;
ROM[5663] <= 32'b00000000011100000000001000110011;
ROM[5664] <= 32'b00000000001000000000000110110011;
ROM[5665] <= 32'b00000111110000001100000011101111;
ROM[5666] <= 32'b11111111110000010000000100010011;
ROM[5667] <= 32'b00000000000000010010001110000011;
ROM[5668] <= 32'b00000000011100011010000000100011;
ROM[5669] <= 32'b00000000000000000110001110110111;
ROM[5670] <= 32'b10001110000000111000001110010011;
ROM[5671] <= 32'b00000000111000111000001110110011;
ROM[5672] <= 32'b00000000011100010010000000100011;
ROM[5673] <= 32'b00000000010000010000000100010011;
ROM[5674] <= 32'b00000000001100010010000000100011;
ROM[5675] <= 32'b00000000010000010000000100010011;
ROM[5676] <= 32'b00000000010000010010000000100011;
ROM[5677] <= 32'b00000000010000010000000100010011;
ROM[5678] <= 32'b00000000010100010010000000100011;
ROM[5679] <= 32'b00000000010000010000000100010011;
ROM[5680] <= 32'b00000000011000010010000000100011;
ROM[5681] <= 32'b00000000010000010000000100010011;
ROM[5682] <= 32'b00000001010000000000001110010011;
ROM[5683] <= 32'b00000000000000111000001110010011;
ROM[5684] <= 32'b01000000011100010000001110110011;
ROM[5685] <= 32'b00000000011100000000001000110011;
ROM[5686] <= 32'b00000000001000000000000110110011;
ROM[5687] <= 32'b10110010100111111111000011101111;
ROM[5688] <= 32'b11111111110000010000000100010011;
ROM[5689] <= 32'b00000000000000010010001110000011;
ROM[5690] <= 32'b00000000011100011010001000100011;
ROM[5691] <= 32'b00000000010000011010001110000011;
ROM[5692] <= 32'b00000000011100010010000000100011;
ROM[5693] <= 32'b00000000010000010000000100010011;
ROM[5694] <= 32'b00000000000000000110001110110111;
ROM[5695] <= 32'b10010100010000111000001110010011;
ROM[5696] <= 32'b00000000111000111000001110110011;
ROM[5697] <= 32'b00000000011100010010000000100011;
ROM[5698] <= 32'b00000000010000010000000100010011;
ROM[5699] <= 32'b00000000001100010010000000100011;
ROM[5700] <= 32'b00000000010000010000000100010011;
ROM[5701] <= 32'b00000000010000010010000000100011;
ROM[5702] <= 32'b00000000010000010000000100010011;
ROM[5703] <= 32'b00000000010100010010000000100011;
ROM[5704] <= 32'b00000000010000010000000100010011;
ROM[5705] <= 32'b00000000011000010010000000100011;
ROM[5706] <= 32'b00000000010000010000000100010011;
ROM[5707] <= 32'b00000001010000000000001110010011;
ROM[5708] <= 32'b00000000000000111000001110010011;
ROM[5709] <= 32'b01000000011100010000001110110011;
ROM[5710] <= 32'b00000000011100000000001000110011;
ROM[5711] <= 32'b00000000001000000000000110110011;
ROM[5712] <= 32'b00001100100000001101000011101111;
ROM[5713] <= 32'b11111111110000010000000100010011;
ROM[5714] <= 32'b00000000000000010010001110000011;
ROM[5715] <= 32'b11111111110000010000000100010011;
ROM[5716] <= 32'b00000000000000010010010000000011;
ROM[5717] <= 32'b00000000011101000010010010110011;
ROM[5718] <= 32'b00000000100000111010010100110011;
ROM[5719] <= 32'b00000000101001001000001110110011;
ROM[5720] <= 32'b00000000000100111000001110010011;
ROM[5721] <= 32'b00000000000100111111001110010011;
ROM[5722] <= 32'b01000000011100000000001110110011;
ROM[5723] <= 32'b00000000000100111000001110010011;
ROM[5724] <= 32'b01000000011100000000001110110011;
ROM[5725] <= 32'b00000000000100111000001110010011;
ROM[5726] <= 32'b00000000000000111000101001100011;
ROM[5727] <= 32'b00000000000000000110001110110111;
ROM[5728] <= 32'b10111010110000111000001110010011;
ROM[5729] <= 32'b00000000111000111000001110110011;
ROM[5730] <= 32'b00000000000000111000000011100111;
ROM[5731] <= 32'b00000000010000011010001110000011;
ROM[5732] <= 32'b00000000011100010010000000100011;
ROM[5733] <= 32'b00000000010000010000000100010011;
ROM[5734] <= 32'b00000000000000000110001110110111;
ROM[5735] <= 32'b10011110010000111000001110010011;
ROM[5736] <= 32'b00000000111000111000001110110011;
ROM[5737] <= 32'b00000000011100010010000000100011;
ROM[5738] <= 32'b00000000010000010000000100010011;
ROM[5739] <= 32'b00000000001100010010000000100011;
ROM[5740] <= 32'b00000000010000010000000100010011;
ROM[5741] <= 32'b00000000010000010010000000100011;
ROM[5742] <= 32'b00000000010000010000000100010011;
ROM[5743] <= 32'b00000000010100010010000000100011;
ROM[5744] <= 32'b00000000010000010000000100010011;
ROM[5745] <= 32'b00000000011000010010000000100011;
ROM[5746] <= 32'b00000000010000010000000100010011;
ROM[5747] <= 32'b00000001010000000000001110010011;
ROM[5748] <= 32'b00000000000000111000001110010011;
ROM[5749] <= 32'b01000000011100010000001110110011;
ROM[5750] <= 32'b00000000011100000000001000110011;
ROM[5751] <= 32'b00000000001000000000000110110011;
ROM[5752] <= 32'b00000110110000001101000011101111;
ROM[5753] <= 32'b11111111110000010000000100010011;
ROM[5754] <= 32'b00000000000000010010001110000011;
ROM[5755] <= 32'b11111111110000010000000100010011;
ROM[5756] <= 32'b00000000000000010010010000000011;
ROM[5757] <= 32'b00000000011101000010010010110011;
ROM[5758] <= 32'b00000000100000111010010100110011;
ROM[5759] <= 32'b00000000101001001000001110110011;
ROM[5760] <= 32'b00000000000100111000001110010011;
ROM[5761] <= 32'b00000000000100111111001110010011;
ROM[5762] <= 32'b00000000000000111000101001100011;
ROM[5763] <= 32'b00000000000000000110001110110111;
ROM[5764] <= 32'b10100010000000111000001110010011;
ROM[5765] <= 32'b00000000111000111000001110110011;
ROM[5766] <= 32'b00000000000000111000000011100111;
ROM[5767] <= 32'b00001100010000000000000011101111;
ROM[5768] <= 32'b00000000000000011010001110000011;
ROM[5769] <= 32'b00000000011100010010000000100011;
ROM[5770] <= 32'b00000000010000010000000100010011;
ROM[5771] <= 32'b00000000000000000110001110110111;
ROM[5772] <= 32'b10100111100000111000001110010011;
ROM[5773] <= 32'b00000000111000111000001110110011;
ROM[5774] <= 32'b00000000011100010010000000100011;
ROM[5775] <= 32'b00000000010000010000000100010011;
ROM[5776] <= 32'b00000000001100010010000000100011;
ROM[5777] <= 32'b00000000010000010000000100010011;
ROM[5778] <= 32'b00000000010000010010000000100011;
ROM[5779] <= 32'b00000000010000010000000100010011;
ROM[5780] <= 32'b00000000010100010010000000100011;
ROM[5781] <= 32'b00000000010000010000000100010011;
ROM[5782] <= 32'b00000000011000010010000000100011;
ROM[5783] <= 32'b00000000010000010000000100010011;
ROM[5784] <= 32'b00000001010000000000001110010011;
ROM[5785] <= 32'b00000000010000111000001110010011;
ROM[5786] <= 32'b01000000011100010000001110110011;
ROM[5787] <= 32'b00000000011100000000001000110011;
ROM[5788] <= 32'b00000000001000000000000110110011;
ROM[5789] <= 32'b00111100010000001100000011101111;
ROM[5790] <= 32'b11111111110000010000000100010011;
ROM[5791] <= 32'b00000000000000010010001110000011;
ROM[5792] <= 32'b00000000011101100010000000100011;
ROM[5793] <= 32'b00000000000000000110001110110111;
ROM[5794] <= 32'b10101101000000111000001110010011;
ROM[5795] <= 32'b00000000111000111000001110110011;
ROM[5796] <= 32'b00000000011100010010000000100011;
ROM[5797] <= 32'b00000000010000010000000100010011;
ROM[5798] <= 32'b00000000001100010010000000100011;
ROM[5799] <= 32'b00000000010000010000000100010011;
ROM[5800] <= 32'b00000000010000010010000000100011;
ROM[5801] <= 32'b00000000010000010000000100010011;
ROM[5802] <= 32'b00000000010100010010000000100011;
ROM[5803] <= 32'b00000000010000010000000100010011;
ROM[5804] <= 32'b00000000011000010010000000100011;
ROM[5805] <= 32'b00000000010000010000000100010011;
ROM[5806] <= 32'b00000001010000000000001110010011;
ROM[5807] <= 32'b00000000000000111000001110010011;
ROM[5808] <= 32'b01000000011100010000001110110011;
ROM[5809] <= 32'b00000000011100000000001000110011;
ROM[5810] <= 32'b00000000001000000000000110110011;
ROM[5811] <= 32'b00010000110000001011000011101111;
ROM[5812] <= 32'b11111111110000010000000100010011;
ROM[5813] <= 32'b00000000000000010010001110000011;
ROM[5814] <= 32'b00000000011101100010000000100011;
ROM[5815] <= 32'b00000111010000000000000011101111;
ROM[5816] <= 32'b00000000000000011010001110000011;
ROM[5817] <= 32'b00000000011100010010000000100011;
ROM[5818] <= 32'b00000000010000010000000100010011;
ROM[5819] <= 32'b00000000010000011010001110000011;
ROM[5820] <= 32'b00000000011100010010000000100011;
ROM[5821] <= 32'b00000000010000010000000100010011;
ROM[5822] <= 32'b00000000000000000110001110110111;
ROM[5823] <= 32'b10110100010000111000001110010011;
ROM[5824] <= 32'b00000000111000111000001110110011;
ROM[5825] <= 32'b00000000011100010010000000100011;
ROM[5826] <= 32'b00000000010000010000000100010011;
ROM[5827] <= 32'b00000000001100010010000000100011;
ROM[5828] <= 32'b00000000010000010000000100010011;
ROM[5829] <= 32'b00000000010000010010000000100011;
ROM[5830] <= 32'b00000000010000010000000100010011;
ROM[5831] <= 32'b00000000010100010010000000100011;
ROM[5832] <= 32'b00000000010000010000000100010011;
ROM[5833] <= 32'b00000000011000010010000000100011;
ROM[5834] <= 32'b00000000010000010000000100010011;
ROM[5835] <= 32'b00000001010000000000001110010011;
ROM[5836] <= 32'b00000000100000111000001110010011;
ROM[5837] <= 32'b01000000011100010000001110110011;
ROM[5838] <= 32'b00000000011100000000001000110011;
ROM[5839] <= 32'b00000000001000000000000110110011;
ROM[5840] <= 32'b00010111110000001100000011101111;
ROM[5841] <= 32'b11111111110000010000000100010011;
ROM[5842] <= 32'b00000000000000010010001110000011;
ROM[5843] <= 32'b00000000011101100010000000100011;
ROM[5844] <= 32'b00000000000000000110001110110111;
ROM[5845] <= 32'b10111001110000111000001110010011;
ROM[5846] <= 32'b00000000111000111000001110110011;
ROM[5847] <= 32'b00000000011100010010000000100011;
ROM[5848] <= 32'b00000000010000010000000100010011;
ROM[5849] <= 32'b00000000001100010010000000100011;
ROM[5850] <= 32'b00000000010000010000000100010011;
ROM[5851] <= 32'b00000000010000010010000000100011;
ROM[5852] <= 32'b00000000010000010000000100010011;
ROM[5853] <= 32'b00000000010100010010000000100011;
ROM[5854] <= 32'b00000000010000010000000100010011;
ROM[5855] <= 32'b00000000011000010010000000100011;
ROM[5856] <= 32'b00000000010000010000000100010011;
ROM[5857] <= 32'b00000001010000000000001110010011;
ROM[5858] <= 32'b00000000000000111000001110010011;
ROM[5859] <= 32'b01000000011100010000001110110011;
ROM[5860] <= 32'b00000000011100000000001000110011;
ROM[5861] <= 32'b00000000001000000000000110110011;
ROM[5862] <= 32'b10000110110111111111000011101111;
ROM[5863] <= 32'b11111111110000010000000100010011;
ROM[5864] <= 32'b00000000000000010010001110000011;
ROM[5865] <= 32'b00000000011100011010001000100011;
ROM[5866] <= 32'b11010100010111111111000011101111;
ROM[5867] <= 32'b00000000000000011010001110000011;
ROM[5868] <= 32'b00000000011100010010000000100011;
ROM[5869] <= 32'b00000000010000010000000100010011;
ROM[5870] <= 32'b00000001010000000000001110010011;
ROM[5871] <= 32'b01000000011100011000001110110011;
ROM[5872] <= 32'b00000000000000111010000010000011;
ROM[5873] <= 32'b11111111110000010000000100010011;
ROM[5874] <= 32'b00000000000000010010001110000011;
ROM[5875] <= 32'b00000000011100100010000000100011;
ROM[5876] <= 32'b00000000010000100000000100010011;
ROM[5877] <= 32'b00000001010000000000001110010011;
ROM[5878] <= 32'b01000000011100011000001110110011;
ROM[5879] <= 32'b00000000010000111010000110000011;
ROM[5880] <= 32'b00000000100000111010001000000011;
ROM[5881] <= 32'b00000000110000111010001010000011;
ROM[5882] <= 32'b00000001000000111010001100000011;
ROM[5883] <= 32'b00000000000000001000000011100111;
ROM[5884] <= 32'b00000000000000010010000000100011;
ROM[5885] <= 32'b00000000010000010000000100010011;
ROM[5886] <= 32'b00000000000000100010001110000011;
ROM[5887] <= 32'b00000000011100010010000000100011;
ROM[5888] <= 32'b00000000010000010000000100010011;
ROM[5889] <= 32'b00000000000000000110001110110111;
ROM[5890] <= 32'b11000101000000111000001110010011;
ROM[5891] <= 32'b00000000111000111000001110110011;
ROM[5892] <= 32'b00000000011100010010000000100011;
ROM[5893] <= 32'b00000000010000010000000100010011;
ROM[5894] <= 32'b00000000001100010010000000100011;
ROM[5895] <= 32'b00000000010000010000000100010011;
ROM[5896] <= 32'b00000000010000010010000000100011;
ROM[5897] <= 32'b00000000010000010000000100010011;
ROM[5898] <= 32'b00000000010100010010000000100011;
ROM[5899] <= 32'b00000000010000010000000100010011;
ROM[5900] <= 32'b00000000011000010010000000100011;
ROM[5901] <= 32'b00000000010000010000000100010011;
ROM[5902] <= 32'b00000001010000000000001110010011;
ROM[5903] <= 32'b00000000010000111000001110010011;
ROM[5904] <= 32'b01000000011100010000001110110011;
ROM[5905] <= 32'b00000000011100000000001000110011;
ROM[5906] <= 32'b00000000001000000000000110110011;
ROM[5907] <= 32'b10110111000111111111000011101111;
ROM[5908] <= 32'b11111111110000010000000100010011;
ROM[5909] <= 32'b00000000000000010010001110000011;
ROM[5910] <= 32'b00000000011100011010000000100011;
ROM[5911] <= 32'b00000000000000011010001110000011;
ROM[5912] <= 32'b00000000011100010010000000100011;
ROM[5913] <= 32'b00000000010000010000000100010011;
ROM[5914] <= 32'b00000000000000000110001110110111;
ROM[5915] <= 32'b11001011010000111000001110010011;
ROM[5916] <= 32'b00000000111000111000001110110011;
ROM[5917] <= 32'b00000000011100010010000000100011;
ROM[5918] <= 32'b00000000010000010000000100010011;
ROM[5919] <= 32'b00000000001100010010000000100011;
ROM[5920] <= 32'b00000000010000010000000100010011;
ROM[5921] <= 32'b00000000010000010010000000100011;
ROM[5922] <= 32'b00000000010000010000000100010011;
ROM[5923] <= 32'b00000000010100010010000000100011;
ROM[5924] <= 32'b00000000010000010000000100010011;
ROM[5925] <= 32'b00000000011000010010000000100011;
ROM[5926] <= 32'b00000000010000010000000100010011;
ROM[5927] <= 32'b00000001010000000000001110010011;
ROM[5928] <= 32'b00000000010000111000001110010011;
ROM[5929] <= 32'b01000000011100010000001110110011;
ROM[5930] <= 32'b00000000011100000000001000110011;
ROM[5931] <= 32'b00000000001000000000000110110011;
ROM[5932] <= 32'b00100011100000001100000011101111;
ROM[5933] <= 32'b00000001010000000000001110010011;
ROM[5934] <= 32'b01000000011100011000001110110011;
ROM[5935] <= 32'b00000000000000111010000010000011;
ROM[5936] <= 32'b11111111110000010000000100010011;
ROM[5937] <= 32'b00000000000000010010001110000011;
ROM[5938] <= 32'b00000000011100100010000000100011;
ROM[5939] <= 32'b00000000010000100000000100010011;
ROM[5940] <= 32'b00000001010000000000001110010011;
ROM[5941] <= 32'b01000000011100011000001110110011;
ROM[5942] <= 32'b00000000010000111010000110000011;
ROM[5943] <= 32'b00000000100000111010001000000011;
ROM[5944] <= 32'b00000000110000111010001010000011;
ROM[5945] <= 32'b00000001000000111010001100000011;
ROM[5946] <= 32'b00000000000000001000000011100111;
ROM[5947] <= 32'b00000000000000010010000000100011;
ROM[5948] <= 32'b00000000010000010000000100010011;
ROM[5949] <= 32'b00000000000000010010000000100011;
ROM[5950] <= 32'b00000000010000010000000100010011;
ROM[5951] <= 32'b00000000000000010010000000100011;
ROM[5952] <= 32'b00000000010000010000000100010011;
ROM[5953] <= 32'b00000000000000010010000000100011;
ROM[5954] <= 32'b00000000010000010000000100010011;
ROM[5955] <= 32'b00000000000000010010000000100011;
ROM[5956] <= 32'b00000000010000010000000100010011;
ROM[5957] <= 32'b00000000000000010010000000100011;
ROM[5958] <= 32'b00000000010000010000000100010011;
ROM[5959] <= 32'b00000000000000010010000000100011;
ROM[5960] <= 32'b00000000010000010000000100010011;
ROM[5961] <= 32'b00000000000000010010000000100011;
ROM[5962] <= 32'b00000000010000010000000100010011;
ROM[5963] <= 32'b00000000000000010010000000100011;
ROM[5964] <= 32'b00000000010000010000000100010011;
ROM[5965] <= 32'b00000000000000010010000000100011;
ROM[5966] <= 32'b00000000010000010000000100010011;
ROM[5967] <= 32'b00000000000000010010000000100011;
ROM[5968] <= 32'b00000000010000010000000100010011;
ROM[5969] <= 32'b00000000000000010010000000100011;
ROM[5970] <= 32'b00000000010000010000000100010011;
ROM[5971] <= 32'b00000000000000010010000000100011;
ROM[5972] <= 32'b00000000010000010000000100010011;
ROM[5973] <= 32'b00000000000000010010000000100011;
ROM[5974] <= 32'b00000000010000010000000100010011;
ROM[5975] <= 32'b00000000000000010010000000100011;
ROM[5976] <= 32'b00000000010000010000000100010011;
ROM[5977] <= 32'b00000000000000010010000000100011;
ROM[5978] <= 32'b00000000010000010000000100010011;
ROM[5979] <= 32'b00000000000000010010000000100011;
ROM[5980] <= 32'b00000000010000010000000100010011;
ROM[5981] <= 32'b00000000000000010010000000100011;
ROM[5982] <= 32'b00000000010000010000000100010011;
ROM[5983] <= 32'b00000000000000010010000000100011;
ROM[5984] <= 32'b00000000010000010000000100010011;
ROM[5985] <= 32'b00000000000000010010000000100011;
ROM[5986] <= 32'b00000000010000010000000100010011;
ROM[5987] <= 32'b00000000000000010010000000100011;
ROM[5988] <= 32'b00000000010000010000000100010011;
ROM[5989] <= 32'b00000000000000010010000000100011;
ROM[5990] <= 32'b00000000010000010000000100010011;
ROM[5991] <= 32'b00000000000000010010000000100011;
ROM[5992] <= 32'b00000000010000010000000100010011;
ROM[5993] <= 32'b00000000000000010010000000100011;
ROM[5994] <= 32'b00000000010000010000000100010011;
ROM[5995] <= 32'b00000100001100000000001110010011;
ROM[5996] <= 32'b00000100011100011010010000100011;
ROM[5997] <= 32'b00000100110000000000001110010011;
ROM[5998] <= 32'b00000100011100011010001000100011;
ROM[5999] <= 32'b00000100011000000000001110010011;
ROM[6000] <= 32'b00000100011100011010100000100011;
ROM[6001] <= 32'b00000101000100000000001110010011;
ROM[6002] <= 32'b00000100011100011010101000100011;
ROM[6003] <= 32'b00000100010100000000001110010011;
ROM[6004] <= 32'b00000100011100011010011000100011;
ROM[6005] <= 32'b00000101001100000000001110010011;
ROM[6006] <= 32'b00000100011100011010110000100011;
ROM[6007] <= 32'b00000100100000000000001110010011;
ROM[6008] <= 32'b00000100011100011010111000100011;
ROM[6009] <= 32'b00000000000100000000001110010011;
ROM[6010] <= 32'b00000000011100010010000000100011;
ROM[6011] <= 32'b00000000010000010000000100010011;
ROM[6012] <= 32'b00000000000000000110001110110111;
ROM[6013] <= 32'b11100011110000111000001110010011;
ROM[6014] <= 32'b00000000111000111000001110110011;
ROM[6015] <= 32'b00000000011100010010000000100011;
ROM[6016] <= 32'b00000000010000010000000100010011;
ROM[6017] <= 32'b00000000001100010010000000100011;
ROM[6018] <= 32'b00000000010000010000000100010011;
ROM[6019] <= 32'b00000000010000010010000000100011;
ROM[6020] <= 32'b00000000010000010000000100010011;
ROM[6021] <= 32'b00000000010100010010000000100011;
ROM[6022] <= 32'b00000000010000010000000100010011;
ROM[6023] <= 32'b00000000011000010010000000100011;
ROM[6024] <= 32'b00000000010000010000000100010011;
ROM[6025] <= 32'b00000001010000000000001110010011;
ROM[6026] <= 32'b00000000010000111000001110010011;
ROM[6027] <= 32'b01000000011100010000001110110011;
ROM[6028] <= 32'b00000000011100000000001000110011;
ROM[6029] <= 32'b00000000001000000000000110110011;
ROM[6030] <= 32'b00101100100100001011000011101111;
ROM[6031] <= 32'b11111111110000010000000100010011;
ROM[6032] <= 32'b00000000000000010010001110000011;
ROM[6033] <= 32'b00000000011100011010011000100011;
ROM[6034] <= 32'b00000000110000011010001110000011;
ROM[6035] <= 32'b00000000011100010010000000100011;
ROM[6036] <= 32'b00000000010000010000000100010011;
ROM[6037] <= 32'b00000010000000000000001110010011;
ROM[6038] <= 32'b00000000011100010010000000100011;
ROM[6039] <= 32'b00000000010000010000000100010011;
ROM[6040] <= 32'b00000000000000000110001110110111;
ROM[6041] <= 32'b11101010110000111000001110010011;
ROM[6042] <= 32'b00000000111000111000001110110011;
ROM[6043] <= 32'b00000000011100010010000000100011;
ROM[6044] <= 32'b00000000010000010000000100010011;
ROM[6045] <= 32'b00000000001100010010000000100011;
ROM[6046] <= 32'b00000000010000010000000100010011;
ROM[6047] <= 32'b00000000010000010010000000100011;
ROM[6048] <= 32'b00000000010000010000000100010011;
ROM[6049] <= 32'b00000000010100010010000000100011;
ROM[6050] <= 32'b00000000010000010000000100010011;
ROM[6051] <= 32'b00000000011000010010000000100011;
ROM[6052] <= 32'b00000000010000010000000100010011;
ROM[6053] <= 32'b00000001010000000000001110010011;
ROM[6054] <= 32'b00000000100000111000001110010011;
ROM[6055] <= 32'b01000000011100010000001110110011;
ROM[6056] <= 32'b00000000011100000000001000110011;
ROM[6057] <= 32'b00000000001000000000000110110011;
ROM[6058] <= 32'b01100001010100001011000011101111;
ROM[6059] <= 32'b11111111110000010000000100010011;
ROM[6060] <= 32'b00000000000000010010001110000011;
ROM[6061] <= 32'b00000000011101100010000000100011;
ROM[6062] <= 32'b00000000110000011010001110000011;
ROM[6063] <= 32'b00000000011100011010011000100011;
ROM[6064] <= 32'b00000000100100000000001110010011;
ROM[6065] <= 32'b00000000011100010010000000100011;
ROM[6066] <= 32'b00000000010000010000000100010011;
ROM[6067] <= 32'b00000000000000000110001110110111;
ROM[6068] <= 32'b11110001100000111000001110010011;
ROM[6069] <= 32'b00000000111000111000001110110011;
ROM[6070] <= 32'b00000000011100010010000000100011;
ROM[6071] <= 32'b00000000010000010000000100010011;
ROM[6072] <= 32'b00000000001100010010000000100011;
ROM[6073] <= 32'b00000000010000010000000100010011;
ROM[6074] <= 32'b00000000010000010010000000100011;
ROM[6075] <= 32'b00000000010000010000000100010011;
ROM[6076] <= 32'b00000000010100010010000000100011;
ROM[6077] <= 32'b00000000010000010000000100010011;
ROM[6078] <= 32'b00000000011000010010000000100011;
ROM[6079] <= 32'b00000000010000010000000100010011;
ROM[6080] <= 32'b00000001010000000000001110010011;
ROM[6081] <= 32'b00000000010000111000001110010011;
ROM[6082] <= 32'b01000000011100010000001110110011;
ROM[6083] <= 32'b00000000011100000000001000110011;
ROM[6084] <= 32'b00000000001000000000000110110011;
ROM[6085] <= 32'b00011110110100001011000011101111;
ROM[6086] <= 32'b11111111110000010000000100010011;
ROM[6087] <= 32'b00000000000000010010001110000011;
ROM[6088] <= 32'b00000000011100011010010000100011;
ROM[6089] <= 32'b00000000100000011010001110000011;
ROM[6090] <= 32'b00000000011100010010000000100011;
ROM[6091] <= 32'b00000000010000010000000100010011;
ROM[6092] <= 32'b00000110010000000000001110010011;
ROM[6093] <= 32'b00000000011100010010000000100011;
ROM[6094] <= 32'b00000000010000010000000100010011;
ROM[6095] <= 32'b00000000000000000110001110110111;
ROM[6096] <= 32'b11111000100000111000001110010011;
ROM[6097] <= 32'b00000000111000111000001110110011;
ROM[6098] <= 32'b00000000011100010010000000100011;
ROM[6099] <= 32'b00000000010000010000000100010011;
ROM[6100] <= 32'b00000000001100010010000000100011;
ROM[6101] <= 32'b00000000010000010000000100010011;
ROM[6102] <= 32'b00000000010000010010000000100011;
ROM[6103] <= 32'b00000000010000010000000100010011;
ROM[6104] <= 32'b00000000010100010010000000100011;
ROM[6105] <= 32'b00000000010000010000000100010011;
ROM[6106] <= 32'b00000000011000010010000000100011;
ROM[6107] <= 32'b00000000010000010000000100010011;
ROM[6108] <= 32'b00000001010000000000001110010011;
ROM[6109] <= 32'b00000000100000111000001110010011;
ROM[6110] <= 32'b01000000011100010000001110110011;
ROM[6111] <= 32'b00000000011100000000001000110011;
ROM[6112] <= 32'b00000000001000000000000110110011;
ROM[6113] <= 32'b01010011100100001011000011101111;
ROM[6114] <= 32'b11111111110000010000000100010011;
ROM[6115] <= 32'b00000000000000010010001110000011;
ROM[6116] <= 32'b00000000011101100010000000100011;
ROM[6117] <= 32'b00000000100000011010001110000011;
ROM[6118] <= 32'b00000000011100010010000000100011;
ROM[6119] <= 32'b00000000010000010000000100010011;
ROM[6120] <= 32'b00000110000100000000001110010011;
ROM[6121] <= 32'b00000000011100010010000000100011;
ROM[6122] <= 32'b00000000010000010000000100010011;
ROM[6123] <= 32'b00000000000000000110001110110111;
ROM[6124] <= 32'b11111111100000111000001110010011;
ROM[6125] <= 32'b00000000111000111000001110110011;
ROM[6126] <= 32'b00000000011100010010000000100011;
ROM[6127] <= 32'b00000000010000010000000100010011;
ROM[6128] <= 32'b00000000001100010010000000100011;
ROM[6129] <= 32'b00000000010000010000000100010011;
ROM[6130] <= 32'b00000000010000010010000000100011;
ROM[6131] <= 32'b00000000010000010000000100010011;
ROM[6132] <= 32'b00000000010100010010000000100011;
ROM[6133] <= 32'b00000000010000010000000100010011;
ROM[6134] <= 32'b00000000011000010010000000100011;
ROM[6135] <= 32'b00000000010000010000000100010011;
ROM[6136] <= 32'b00000001010000000000001110010011;
ROM[6137] <= 32'b00000000100000111000001110010011;
ROM[6138] <= 32'b01000000011100010000001110110011;
ROM[6139] <= 32'b00000000011100000000001000110011;
ROM[6140] <= 32'b00000000001000000000000110110011;
ROM[6141] <= 32'b01001100100100001011000011101111;
ROM[6142] <= 32'b11111111110000010000000100010011;
ROM[6143] <= 32'b00000000000000010010001110000011;
ROM[6144] <= 32'b00000000011101100010000000100011;
ROM[6145] <= 32'b00000000100000011010001110000011;
ROM[6146] <= 32'b00000000011100010010000000100011;
ROM[6147] <= 32'b00000000010000010000000100010011;
ROM[6148] <= 32'b00000111011000000000001110010011;
ROM[6149] <= 32'b00000000011100010010000000100011;
ROM[6150] <= 32'b00000000010000010000000100010011;
ROM[6151] <= 32'b00000000000000000110001110110111;
ROM[6152] <= 32'b00000110100000111000001110010011;
ROM[6153] <= 32'b00000000111000111000001110110011;
ROM[6154] <= 32'b00000000011100010010000000100011;
ROM[6155] <= 32'b00000000010000010000000100010011;
ROM[6156] <= 32'b00000000001100010010000000100011;
ROM[6157] <= 32'b00000000010000010000000100010011;
ROM[6158] <= 32'b00000000010000010010000000100011;
ROM[6159] <= 32'b00000000010000010000000100010011;
ROM[6160] <= 32'b00000000010100010010000000100011;
ROM[6161] <= 32'b00000000010000010000000100010011;
ROM[6162] <= 32'b00000000011000010010000000100011;
ROM[6163] <= 32'b00000000010000010000000100010011;
ROM[6164] <= 32'b00000001010000000000001110010011;
ROM[6165] <= 32'b00000000100000111000001110010011;
ROM[6166] <= 32'b01000000011100010000001110110011;
ROM[6167] <= 32'b00000000011100000000001000110011;
ROM[6168] <= 32'b00000000001000000000000110110011;
ROM[6169] <= 32'b01000101100100001011000011101111;
ROM[6170] <= 32'b11111111110000010000000100010011;
ROM[6171] <= 32'b00000000000000010010001110000011;
ROM[6172] <= 32'b00000000011101100010000000100011;
ROM[6173] <= 32'b00000000100000011010001110000011;
ROM[6174] <= 32'b00000000011100010010000000100011;
ROM[6175] <= 32'b00000000010000010000000100010011;
ROM[6176] <= 32'b00000110100100000000001110010011;
ROM[6177] <= 32'b00000000011100010010000000100011;
ROM[6178] <= 32'b00000000010000010000000100010011;
ROM[6179] <= 32'b00000000000000000110001110110111;
ROM[6180] <= 32'b00001101100000111000001110010011;
ROM[6181] <= 32'b00000000111000111000001110110011;
ROM[6182] <= 32'b00000000011100010010000000100011;
ROM[6183] <= 32'b00000000010000010000000100010011;
ROM[6184] <= 32'b00000000001100010010000000100011;
ROM[6185] <= 32'b00000000010000010000000100010011;
ROM[6186] <= 32'b00000000010000010010000000100011;
ROM[6187] <= 32'b00000000010000010000000100010011;
ROM[6188] <= 32'b00000000010100010010000000100011;
ROM[6189] <= 32'b00000000010000010000000100010011;
ROM[6190] <= 32'b00000000011000010010000000100011;
ROM[6191] <= 32'b00000000010000010000000100010011;
ROM[6192] <= 32'b00000001010000000000001110010011;
ROM[6193] <= 32'b00000000100000111000001110010011;
ROM[6194] <= 32'b01000000011100010000001110110011;
ROM[6195] <= 32'b00000000011100000000001000110011;
ROM[6196] <= 32'b00000000001000000000000110110011;
ROM[6197] <= 32'b00111110100100001011000011101111;
ROM[6198] <= 32'b11111111110000010000000100010011;
ROM[6199] <= 32'b00000000000000010010001110000011;
ROM[6200] <= 32'b00000000011101100010000000100011;
ROM[6201] <= 32'b00000000100000011010001110000011;
ROM[6202] <= 32'b00000000011100010010000000100011;
ROM[6203] <= 32'b00000000010000010000000100010011;
ROM[6204] <= 32'b00000110111000000000001110010011;
ROM[6205] <= 32'b00000000011100010010000000100011;
ROM[6206] <= 32'b00000000010000010000000100010011;
ROM[6207] <= 32'b00000000000000000110001110110111;
ROM[6208] <= 32'b00010100100000111000001110010011;
ROM[6209] <= 32'b00000000111000111000001110110011;
ROM[6210] <= 32'b00000000011100010010000000100011;
ROM[6211] <= 32'b00000000010000010000000100010011;
ROM[6212] <= 32'b00000000001100010010000000100011;
ROM[6213] <= 32'b00000000010000010000000100010011;
ROM[6214] <= 32'b00000000010000010010000000100011;
ROM[6215] <= 32'b00000000010000010000000100010011;
ROM[6216] <= 32'b00000000010100010010000000100011;
ROM[6217] <= 32'b00000000010000010000000100010011;
ROM[6218] <= 32'b00000000011000010010000000100011;
ROM[6219] <= 32'b00000000010000010000000100010011;
ROM[6220] <= 32'b00000001010000000000001110010011;
ROM[6221] <= 32'b00000000100000111000001110010011;
ROM[6222] <= 32'b01000000011100010000001110110011;
ROM[6223] <= 32'b00000000011100000000001000110011;
ROM[6224] <= 32'b00000000001000000000000110110011;
ROM[6225] <= 32'b00110111100100001011000011101111;
ROM[6226] <= 32'b11111111110000010000000100010011;
ROM[6227] <= 32'b00000000000000010010001110000011;
ROM[6228] <= 32'b00000000011101100010000000100011;
ROM[6229] <= 32'b00000000100000011010001110000011;
ROM[6230] <= 32'b00000000011100010010000000100011;
ROM[6231] <= 32'b00000000010000010000000100010011;
ROM[6232] <= 32'b00000110001100000000001110010011;
ROM[6233] <= 32'b00000000011100010010000000100011;
ROM[6234] <= 32'b00000000010000010000000100010011;
ROM[6235] <= 32'b00000000000000000110001110110111;
ROM[6236] <= 32'b00011011100000111000001110010011;
ROM[6237] <= 32'b00000000111000111000001110110011;
ROM[6238] <= 32'b00000000011100010010000000100011;
ROM[6239] <= 32'b00000000010000010000000100010011;
ROM[6240] <= 32'b00000000001100010010000000100011;
ROM[6241] <= 32'b00000000010000010000000100010011;
ROM[6242] <= 32'b00000000010000010010000000100011;
ROM[6243] <= 32'b00000000010000010000000100010011;
ROM[6244] <= 32'b00000000010100010010000000100011;
ROM[6245] <= 32'b00000000010000010000000100010011;
ROM[6246] <= 32'b00000000011000010010000000100011;
ROM[6247] <= 32'b00000000010000010000000100010011;
ROM[6248] <= 32'b00000001010000000000001110010011;
ROM[6249] <= 32'b00000000100000111000001110010011;
ROM[6250] <= 32'b01000000011100010000001110110011;
ROM[6251] <= 32'b00000000011100000000001000110011;
ROM[6252] <= 32'b00000000001000000000000110110011;
ROM[6253] <= 32'b00110000100100001011000011101111;
ROM[6254] <= 32'b11111111110000010000000100010011;
ROM[6255] <= 32'b00000000000000010010001110000011;
ROM[6256] <= 32'b00000000011101100010000000100011;
ROM[6257] <= 32'b00000000100000011010001110000011;
ROM[6258] <= 32'b00000000011100010010000000100011;
ROM[6259] <= 32'b00000000010000010000000100010011;
ROM[6260] <= 32'b00000110100100000000001110010011;
ROM[6261] <= 32'b00000000011100010010000000100011;
ROM[6262] <= 32'b00000000010000010000000100010011;
ROM[6263] <= 32'b00000000000000000110001110110111;
ROM[6264] <= 32'b00100010100000111000001110010011;
ROM[6265] <= 32'b00000000111000111000001110110011;
ROM[6266] <= 32'b00000000011100010010000000100011;
ROM[6267] <= 32'b00000000010000010000000100010011;
ROM[6268] <= 32'b00000000001100010010000000100011;
ROM[6269] <= 32'b00000000010000010000000100010011;
ROM[6270] <= 32'b00000000010000010010000000100011;
ROM[6271] <= 32'b00000000010000010000000100010011;
ROM[6272] <= 32'b00000000010100010010000000100011;
ROM[6273] <= 32'b00000000010000010000000100010011;
ROM[6274] <= 32'b00000000011000010010000000100011;
ROM[6275] <= 32'b00000000010000010000000100010011;
ROM[6276] <= 32'b00000001010000000000001110010011;
ROM[6277] <= 32'b00000000100000111000001110010011;
ROM[6278] <= 32'b01000000011100010000001110110011;
ROM[6279] <= 32'b00000000011100000000001000110011;
ROM[6280] <= 32'b00000000001000000000000110110011;
ROM[6281] <= 32'b00101001100100001011000011101111;
ROM[6282] <= 32'b11111111110000010000000100010011;
ROM[6283] <= 32'b00000000000000010010001110000011;
ROM[6284] <= 32'b00000000011101100010000000100011;
ROM[6285] <= 32'b00000000100000011010001110000011;
ROM[6286] <= 32'b00000000011100010010000000100011;
ROM[6287] <= 32'b00000000010000010000000100010011;
ROM[6288] <= 32'b00000010010000000000001110010011;
ROM[6289] <= 32'b00000000011100010010000000100011;
ROM[6290] <= 32'b00000000010000010000000100010011;
ROM[6291] <= 32'b00000000000000000110001110110111;
ROM[6292] <= 32'b00101001100000111000001110010011;
ROM[6293] <= 32'b00000000111000111000001110110011;
ROM[6294] <= 32'b00000000011100010010000000100011;
ROM[6295] <= 32'b00000000010000010000000100010011;
ROM[6296] <= 32'b00000000001100010010000000100011;
ROM[6297] <= 32'b00000000010000010000000100010011;
ROM[6298] <= 32'b00000000010000010010000000100011;
ROM[6299] <= 32'b00000000010000010000000100010011;
ROM[6300] <= 32'b00000000010100010010000000100011;
ROM[6301] <= 32'b00000000010000010000000100010011;
ROM[6302] <= 32'b00000000011000010010000000100011;
ROM[6303] <= 32'b00000000010000010000000100010011;
ROM[6304] <= 32'b00000001010000000000001110010011;
ROM[6305] <= 32'b00000000100000111000001110010011;
ROM[6306] <= 32'b01000000011100010000001110110011;
ROM[6307] <= 32'b00000000011100000000001000110011;
ROM[6308] <= 32'b00000000001000000000000110110011;
ROM[6309] <= 32'b00100010100100001011000011101111;
ROM[6310] <= 32'b11111111110000010000000100010011;
ROM[6311] <= 32'b00000000000000010010001110000011;
ROM[6312] <= 32'b00000000011101100010000000100011;
ROM[6313] <= 32'b00000000100000011010001110000011;
ROM[6314] <= 32'b00000000011100010010000000100011;
ROM[6315] <= 32'b00000000010000010000000100010011;
ROM[6316] <= 32'b00000010000000000000001110010011;
ROM[6317] <= 32'b00000000011100010010000000100011;
ROM[6318] <= 32'b00000000010000010000000100010011;
ROM[6319] <= 32'b00000000000000000110001110110111;
ROM[6320] <= 32'b00110000100000111000001110010011;
ROM[6321] <= 32'b00000000111000111000001110110011;
ROM[6322] <= 32'b00000000011100010010000000100011;
ROM[6323] <= 32'b00000000010000010000000100010011;
ROM[6324] <= 32'b00000000001100010010000000100011;
ROM[6325] <= 32'b00000000010000010000000100010011;
ROM[6326] <= 32'b00000000010000010010000000100011;
ROM[6327] <= 32'b00000000010000010000000100010011;
ROM[6328] <= 32'b00000000010100010010000000100011;
ROM[6329] <= 32'b00000000010000010000000100010011;
ROM[6330] <= 32'b00000000011000010010000000100011;
ROM[6331] <= 32'b00000000010000010000000100010011;
ROM[6332] <= 32'b00000001010000000000001110010011;
ROM[6333] <= 32'b00000000100000111000001110010011;
ROM[6334] <= 32'b01000000011100010000001110110011;
ROM[6335] <= 32'b00000000011100000000001000110011;
ROM[6336] <= 32'b00000000001000000000000110110011;
ROM[6337] <= 32'b00011011100100001011000011101111;
ROM[6338] <= 32'b11111111110000010000000100010011;
ROM[6339] <= 32'b00000000000000010010001110000011;
ROM[6340] <= 32'b00000000011101100010000000100011;
ROM[6341] <= 32'b00000000100000011010001110000011;
ROM[6342] <= 32'b00000000011100011010010000100011;
ROM[6343] <= 32'b00000000011100000000001110010011;
ROM[6344] <= 32'b00000000011100010010000000100011;
ROM[6345] <= 32'b00000000010000010000000100010011;
ROM[6346] <= 32'b00000000000000000110001110110111;
ROM[6347] <= 32'b00110111010000111000001110010011;
ROM[6348] <= 32'b00000000111000111000001110110011;
ROM[6349] <= 32'b00000000011100010010000000100011;
ROM[6350] <= 32'b00000000010000010000000100010011;
ROM[6351] <= 32'b00000000001100010010000000100011;
ROM[6352] <= 32'b00000000010000010000000100010011;
ROM[6353] <= 32'b00000000010000010010000000100011;
ROM[6354] <= 32'b00000000010000010000000100010011;
ROM[6355] <= 32'b00000000010100010010000000100011;
ROM[6356] <= 32'b00000000010000010000000100010011;
ROM[6357] <= 32'b00000000011000010010000000100011;
ROM[6358] <= 32'b00000000010000010000000100010011;
ROM[6359] <= 32'b00000001010000000000001110010011;
ROM[6360] <= 32'b00000000010000111000001110010011;
ROM[6361] <= 32'b01000000011100010000001110110011;
ROM[6362] <= 32'b00000000011100000000001000110011;
ROM[6363] <= 32'b00000000001000000000000110110011;
ROM[6364] <= 32'b01011001000000001011000011101111;
ROM[6365] <= 32'b11111111110000010000000100010011;
ROM[6366] <= 32'b00000000000000010010001110000011;
ROM[6367] <= 32'b00000000011100011010100000100011;
ROM[6368] <= 32'b00000001000000011010001110000011;
ROM[6369] <= 32'b00000000011100010010000000100011;
ROM[6370] <= 32'b00000000010000010000000100010011;
ROM[6371] <= 32'b00000110100100000000001110010011;
ROM[6372] <= 32'b00000000011100010010000000100011;
ROM[6373] <= 32'b00000000010000010000000100010011;
ROM[6374] <= 32'b00000000000000000110001110110111;
ROM[6375] <= 32'b00111110010000111000001110010011;
ROM[6376] <= 32'b00000000111000111000001110110011;
ROM[6377] <= 32'b00000000011100010010000000100011;
ROM[6378] <= 32'b00000000010000010000000100010011;
ROM[6379] <= 32'b00000000001100010010000000100011;
ROM[6380] <= 32'b00000000010000010000000100010011;
ROM[6381] <= 32'b00000000010000010010000000100011;
ROM[6382] <= 32'b00000000010000010000000100010011;
ROM[6383] <= 32'b00000000010100010010000000100011;
ROM[6384] <= 32'b00000000010000010000000100010011;
ROM[6385] <= 32'b00000000011000010010000000100011;
ROM[6386] <= 32'b00000000010000010000000100010011;
ROM[6387] <= 32'b00000001010000000000001110010011;
ROM[6388] <= 32'b00000000100000111000001110010011;
ROM[6389] <= 32'b01000000011100010000001110110011;
ROM[6390] <= 32'b00000000011100000000001000110011;
ROM[6391] <= 32'b00000000001000000000000110110011;
ROM[6392] <= 32'b00001101110100001011000011101111;
ROM[6393] <= 32'b11111111110000010000000100010011;
ROM[6394] <= 32'b00000000000000010010001110000011;
ROM[6395] <= 32'b00000000011101100010000000100011;
ROM[6396] <= 32'b00000001000000011010001110000011;
ROM[6397] <= 32'b00000000011100010010000000100011;
ROM[6398] <= 32'b00000000010000010000000100010011;
ROM[6399] <= 32'b00000110111000000000001110010011;
ROM[6400] <= 32'b00000000011100010010000000100011;
ROM[6401] <= 32'b00000000010000010000000100010011;
ROM[6402] <= 32'b00000000000000000110001110110111;
ROM[6403] <= 32'b01000101010000111000001110010011;
ROM[6404] <= 32'b00000000111000111000001110110011;
ROM[6405] <= 32'b00000000011100010010000000100011;
ROM[6406] <= 32'b00000000010000010000000100010011;
ROM[6407] <= 32'b00000000001100010010000000100011;
ROM[6408] <= 32'b00000000010000010000000100010011;
ROM[6409] <= 32'b00000000010000010010000000100011;
ROM[6410] <= 32'b00000000010000010000000100010011;
ROM[6411] <= 32'b00000000010100010010000000100011;
ROM[6412] <= 32'b00000000010000010000000100010011;
ROM[6413] <= 32'b00000000011000010010000000100011;
ROM[6414] <= 32'b00000000010000010000000100010011;
ROM[6415] <= 32'b00000001010000000000001110010011;
ROM[6416] <= 32'b00000000100000111000001110010011;
ROM[6417] <= 32'b01000000011100010000001110110011;
ROM[6418] <= 32'b00000000011100000000001000110011;
ROM[6419] <= 32'b00000000001000000000000110110011;
ROM[6420] <= 32'b00000110110100001011000011101111;
ROM[6421] <= 32'b11111111110000010000000100010011;
ROM[6422] <= 32'b00000000000000010010001110000011;
ROM[6423] <= 32'b00000000011101100010000000100011;
ROM[6424] <= 32'b00000001000000011010001110000011;
ROM[6425] <= 32'b00000000011100010010000000100011;
ROM[6426] <= 32'b00000000010000010000000100010011;
ROM[6427] <= 32'b00000111011000000000001110010011;
ROM[6428] <= 32'b00000000011100010010000000100011;
ROM[6429] <= 32'b00000000010000010000000100010011;
ROM[6430] <= 32'b00000000000000000110001110110111;
ROM[6431] <= 32'b01001100010000111000001110010011;
ROM[6432] <= 32'b00000000111000111000001110110011;
ROM[6433] <= 32'b00000000011100010010000000100011;
ROM[6434] <= 32'b00000000010000010000000100010011;
ROM[6435] <= 32'b00000000001100010010000000100011;
ROM[6436] <= 32'b00000000010000010000000100010011;
ROM[6437] <= 32'b00000000010000010010000000100011;
ROM[6438] <= 32'b00000000010000010000000100010011;
ROM[6439] <= 32'b00000000010100010010000000100011;
ROM[6440] <= 32'b00000000010000010000000100010011;
ROM[6441] <= 32'b00000000011000010010000000100011;
ROM[6442] <= 32'b00000000010000010000000100010011;
ROM[6443] <= 32'b00000001010000000000001110010011;
ROM[6444] <= 32'b00000000100000111000001110010011;
ROM[6445] <= 32'b01000000011100010000001110110011;
ROM[6446] <= 32'b00000000011100000000001000110011;
ROM[6447] <= 32'b00000000001000000000000110110011;
ROM[6448] <= 32'b01111111110000001011000011101111;
ROM[6449] <= 32'b11111111110000010000000100010011;
ROM[6450] <= 32'b00000000000000010010001110000011;
ROM[6451] <= 32'b00000000011101100010000000100011;
ROM[6452] <= 32'b00000001000000011010001110000011;
ROM[6453] <= 32'b00000000011100010010000000100011;
ROM[6454] <= 32'b00000000010000010000000100010011;
ROM[6455] <= 32'b00000110000100000000001110010011;
ROM[6456] <= 32'b00000000011100010010000000100011;
ROM[6457] <= 32'b00000000010000010000000100010011;
ROM[6458] <= 32'b00000000000000000110001110110111;
ROM[6459] <= 32'b01010011010000111000001110010011;
ROM[6460] <= 32'b00000000111000111000001110110011;
ROM[6461] <= 32'b00000000011100010010000000100011;
ROM[6462] <= 32'b00000000010000010000000100010011;
ROM[6463] <= 32'b00000000001100010010000000100011;
ROM[6464] <= 32'b00000000010000010000000100010011;
ROM[6465] <= 32'b00000000010000010010000000100011;
ROM[6466] <= 32'b00000000010000010000000100010011;
ROM[6467] <= 32'b00000000010100010010000000100011;
ROM[6468] <= 32'b00000000010000010000000100010011;
ROM[6469] <= 32'b00000000011000010010000000100011;
ROM[6470] <= 32'b00000000010000010000000100010011;
ROM[6471] <= 32'b00000001010000000000001110010011;
ROM[6472] <= 32'b00000000100000111000001110010011;
ROM[6473] <= 32'b01000000011100010000001110110011;
ROM[6474] <= 32'b00000000011100000000001000110011;
ROM[6475] <= 32'b00000000001000000000000110110011;
ROM[6476] <= 32'b01111000110000001011000011101111;
ROM[6477] <= 32'b11111111110000010000000100010011;
ROM[6478] <= 32'b00000000000000010010001110000011;
ROM[6479] <= 32'b00000000011101100010000000100011;
ROM[6480] <= 32'b00000001000000011010001110000011;
ROM[6481] <= 32'b00000000011100010010000000100011;
ROM[6482] <= 32'b00000000010000010000000100010011;
ROM[6483] <= 32'b00000110110000000000001110010011;
ROM[6484] <= 32'b00000000011100010010000000100011;
ROM[6485] <= 32'b00000000010000010000000100010011;
ROM[6486] <= 32'b00000000000000000110001110110111;
ROM[6487] <= 32'b01011010010000111000001110010011;
ROM[6488] <= 32'b00000000111000111000001110110011;
ROM[6489] <= 32'b00000000011100010010000000100011;
ROM[6490] <= 32'b00000000010000010000000100010011;
ROM[6491] <= 32'b00000000001100010010000000100011;
ROM[6492] <= 32'b00000000010000010000000100010011;
ROM[6493] <= 32'b00000000010000010010000000100011;
ROM[6494] <= 32'b00000000010000010000000100010011;
ROM[6495] <= 32'b00000000010100010010000000100011;
ROM[6496] <= 32'b00000000010000010000000100010011;
ROM[6497] <= 32'b00000000011000010010000000100011;
ROM[6498] <= 32'b00000000010000010000000100010011;
ROM[6499] <= 32'b00000001010000000000001110010011;
ROM[6500] <= 32'b00000000100000111000001110010011;
ROM[6501] <= 32'b01000000011100010000001110110011;
ROM[6502] <= 32'b00000000011100000000001000110011;
ROM[6503] <= 32'b00000000001000000000000110110011;
ROM[6504] <= 32'b01110001110000001011000011101111;
ROM[6505] <= 32'b11111111110000010000000100010011;
ROM[6506] <= 32'b00000000000000010010001110000011;
ROM[6507] <= 32'b00000000011101100010000000100011;
ROM[6508] <= 32'b00000001000000011010001110000011;
ROM[6509] <= 32'b00000000011100010010000000100011;
ROM[6510] <= 32'b00000000010000010000000100010011;
ROM[6511] <= 32'b00000110100100000000001110010011;
ROM[6512] <= 32'b00000000011100010010000000100011;
ROM[6513] <= 32'b00000000010000010000000100010011;
ROM[6514] <= 32'b00000000000000000110001110110111;
ROM[6515] <= 32'b01100001010000111000001110010011;
ROM[6516] <= 32'b00000000111000111000001110110011;
ROM[6517] <= 32'b00000000011100010010000000100011;
ROM[6518] <= 32'b00000000010000010000000100010011;
ROM[6519] <= 32'b00000000001100010010000000100011;
ROM[6520] <= 32'b00000000010000010000000100010011;
ROM[6521] <= 32'b00000000010000010010000000100011;
ROM[6522] <= 32'b00000000010000010000000100010011;
ROM[6523] <= 32'b00000000010100010010000000100011;
ROM[6524] <= 32'b00000000010000010000000100010011;
ROM[6525] <= 32'b00000000011000010010000000100011;
ROM[6526] <= 32'b00000000010000010000000100010011;
ROM[6527] <= 32'b00000001010000000000001110010011;
ROM[6528] <= 32'b00000000100000111000001110010011;
ROM[6529] <= 32'b01000000011100010000001110110011;
ROM[6530] <= 32'b00000000011100000000001000110011;
ROM[6531] <= 32'b00000000001000000000000110110011;
ROM[6532] <= 32'b01101010110000001011000011101111;
ROM[6533] <= 32'b11111111110000010000000100010011;
ROM[6534] <= 32'b00000000000000010010001110000011;
ROM[6535] <= 32'b00000000011101100010000000100011;
ROM[6536] <= 32'b00000001000000011010001110000011;
ROM[6537] <= 32'b00000000011100010010000000100011;
ROM[6538] <= 32'b00000000010000010000000100010011;
ROM[6539] <= 32'b00000110010000000000001110010011;
ROM[6540] <= 32'b00000000011100010010000000100011;
ROM[6541] <= 32'b00000000010000010000000100010011;
ROM[6542] <= 32'b00000000000000000110001110110111;
ROM[6543] <= 32'b01101000010000111000001110010011;
ROM[6544] <= 32'b00000000111000111000001110110011;
ROM[6545] <= 32'b00000000011100010010000000100011;
ROM[6546] <= 32'b00000000010000010000000100010011;
ROM[6547] <= 32'b00000000001100010010000000100011;
ROM[6548] <= 32'b00000000010000010000000100010011;
ROM[6549] <= 32'b00000000010000010010000000100011;
ROM[6550] <= 32'b00000000010000010000000100010011;
ROM[6551] <= 32'b00000000010100010010000000100011;
ROM[6552] <= 32'b00000000010000010000000100010011;
ROM[6553] <= 32'b00000000011000010010000000100011;
ROM[6554] <= 32'b00000000010000010000000100010011;
ROM[6555] <= 32'b00000001010000000000001110010011;
ROM[6556] <= 32'b00000000100000111000001110010011;
ROM[6557] <= 32'b01000000011100010000001110110011;
ROM[6558] <= 32'b00000000011100000000001000110011;
ROM[6559] <= 32'b00000000001000000000000110110011;
ROM[6560] <= 32'b01100011110000001011000011101111;
ROM[6561] <= 32'b11111111110000010000000100010011;
ROM[6562] <= 32'b00000000000000010010001110000011;
ROM[6563] <= 32'b00000000011101100010000000100011;
ROM[6564] <= 32'b00000001000000011010001110000011;
ROM[6565] <= 32'b00000000011100011010100000100011;
ROM[6566] <= 32'b00000000000000000000001110010011;
ROM[6567] <= 32'b00000000011100011010000000100011;
ROM[6568] <= 32'b00000000000100000000001110010011;
ROM[6569] <= 32'b00000000011100011010001000100011;
ROM[6570] <= 32'b00000000011000000000001110010011;
ROM[6571] <= 32'b00000000011100010010000000100011;
ROM[6572] <= 32'b00000000010000010000000100010011;
ROM[6573] <= 32'b00000000000000000110001110110111;
ROM[6574] <= 32'b01110000000000111000001110010011;
ROM[6575] <= 32'b00000000111000111000001110110011;
ROM[6576] <= 32'b00000000011100010010000000100011;
ROM[6577] <= 32'b00000000010000010000000100010011;
ROM[6578] <= 32'b00000000001100010010000000100011;
ROM[6579] <= 32'b00000000010000010000000100010011;
ROM[6580] <= 32'b00000000010000010010000000100011;
ROM[6581] <= 32'b00000000010000010000000100010011;
ROM[6582] <= 32'b00000000010100010010000000100011;
ROM[6583] <= 32'b00000000010000010000000100010011;
ROM[6584] <= 32'b00000000011000010010000000100011;
ROM[6585] <= 32'b00000000010000010000000100010011;
ROM[6586] <= 32'b00000001010000000000001110010011;
ROM[6587] <= 32'b00000000010000111000001110010011;
ROM[6588] <= 32'b01000000011100010000001110110011;
ROM[6589] <= 32'b00000000011100000000001000110011;
ROM[6590] <= 32'b00000000001000000000000110110011;
ROM[6591] <= 32'b00100000010000001011000011101111;
ROM[6592] <= 32'b11111111110000010000000100010011;
ROM[6593] <= 32'b00000000000000010010001110000011;
ROM[6594] <= 32'b00000000011100011010101000100011;
ROM[6595] <= 32'b00000001010000011010001110000011;
ROM[6596] <= 32'b00000000011100010010000000100011;
ROM[6597] <= 32'b00000000010000010000000100010011;
ROM[6598] <= 32'b00000010000000000000001110010011;
ROM[6599] <= 32'b00000000011100010010000000100011;
ROM[6600] <= 32'b00000000010000010000000100010011;
ROM[6601] <= 32'b00000000000000000110001110110111;
ROM[6602] <= 32'b01110111000000111000001110010011;
ROM[6603] <= 32'b00000000111000111000001110110011;
ROM[6604] <= 32'b00000000011100010010000000100011;
ROM[6605] <= 32'b00000000010000010000000100010011;
ROM[6606] <= 32'b00000000001100010010000000100011;
ROM[6607] <= 32'b00000000010000010000000100010011;
ROM[6608] <= 32'b00000000010000010010000000100011;
ROM[6609] <= 32'b00000000010000010000000100010011;
ROM[6610] <= 32'b00000000010100010010000000100011;
ROM[6611] <= 32'b00000000010000010000000100010011;
ROM[6612] <= 32'b00000000011000010010000000100011;
ROM[6613] <= 32'b00000000010000010000000100010011;
ROM[6614] <= 32'b00000001010000000000001110010011;
ROM[6615] <= 32'b00000000100000111000001110010011;
ROM[6616] <= 32'b01000000011100010000001110110011;
ROM[6617] <= 32'b00000000011100000000001000110011;
ROM[6618] <= 32'b00000000001000000000000110110011;
ROM[6619] <= 32'b01010101000000001011000011101111;
ROM[6620] <= 32'b11111111110000010000000100010011;
ROM[6621] <= 32'b00000000000000010010001110000011;
ROM[6622] <= 32'b00000000011101100010000000100011;
ROM[6623] <= 32'b00000001010000011010001110000011;
ROM[6624] <= 32'b00000000011100010010000000100011;
ROM[6625] <= 32'b00000000010000010000000100010011;
ROM[6626] <= 32'b00000110011000000000001110010011;
ROM[6627] <= 32'b00000000011100010010000000100011;
ROM[6628] <= 32'b00000000010000010000000100010011;
ROM[6629] <= 32'b00000000000000000110001110110111;
ROM[6630] <= 32'b01111110000000111000001110010011;
ROM[6631] <= 32'b00000000111000111000001110110011;
ROM[6632] <= 32'b00000000011100010010000000100011;
ROM[6633] <= 32'b00000000010000010000000100010011;
ROM[6634] <= 32'b00000000001100010010000000100011;
ROM[6635] <= 32'b00000000010000010000000100010011;
ROM[6636] <= 32'b00000000010000010010000000100011;
ROM[6637] <= 32'b00000000010000010000000100010011;
ROM[6638] <= 32'b00000000010100010010000000100011;
ROM[6639] <= 32'b00000000010000010000000100010011;
ROM[6640] <= 32'b00000000011000010010000000100011;
ROM[6641] <= 32'b00000000010000010000000100010011;
ROM[6642] <= 32'b00000001010000000000001110010011;
ROM[6643] <= 32'b00000000100000111000001110010011;
ROM[6644] <= 32'b01000000011100010000001110110011;
ROM[6645] <= 32'b00000000011100000000001000110011;
ROM[6646] <= 32'b00000000001000000000000110110011;
ROM[6647] <= 32'b01001110000000001011000011101111;
ROM[6648] <= 32'b11111111110000010000000100010011;
ROM[6649] <= 32'b00000000000000010010001110000011;
ROM[6650] <= 32'b00000000011101100010000000100011;
ROM[6651] <= 32'b00000001010000011010001110000011;
ROM[6652] <= 32'b00000000011100010010000000100011;
ROM[6653] <= 32'b00000000010000010000000100010011;
ROM[6654] <= 32'b00000110100100000000001110010011;
ROM[6655] <= 32'b00000000011100010010000000100011;
ROM[6656] <= 32'b00000000010000010000000100010011;
ROM[6657] <= 32'b00000000000000000111001110110111;
ROM[6658] <= 32'b10000101000000111000001110010011;
ROM[6659] <= 32'b00000000111000111000001110110011;
ROM[6660] <= 32'b00000000011100010010000000100011;
ROM[6661] <= 32'b00000000010000010000000100010011;
ROM[6662] <= 32'b00000000001100010010000000100011;
ROM[6663] <= 32'b00000000010000010000000100010011;
ROM[6664] <= 32'b00000000010000010010000000100011;
ROM[6665] <= 32'b00000000010000010000000100010011;
ROM[6666] <= 32'b00000000010100010010000000100011;
ROM[6667] <= 32'b00000000010000010000000100010011;
ROM[6668] <= 32'b00000000011000010010000000100011;
ROM[6669] <= 32'b00000000010000010000000100010011;
ROM[6670] <= 32'b00000001010000000000001110010011;
ROM[6671] <= 32'b00000000100000111000001110010011;
ROM[6672] <= 32'b01000000011100010000001110110011;
ROM[6673] <= 32'b00000000011100000000001000110011;
ROM[6674] <= 32'b00000000001000000000000110110011;
ROM[6675] <= 32'b01000111000000001011000011101111;
ROM[6676] <= 32'b11111111110000010000000100010011;
ROM[6677] <= 32'b00000000000000010010001110000011;
ROM[6678] <= 32'b00000000011101100010000000100011;
ROM[6679] <= 32'b00000001010000011010001110000011;
ROM[6680] <= 32'b00000000011100010010000000100011;
ROM[6681] <= 32'b00000000010000010000000100010011;
ROM[6682] <= 32'b00000110001000000000001110010011;
ROM[6683] <= 32'b00000000011100010010000000100011;
ROM[6684] <= 32'b00000000010000010000000100010011;
ROM[6685] <= 32'b00000000000000000111001110110111;
ROM[6686] <= 32'b10001100000000111000001110010011;
ROM[6687] <= 32'b00000000111000111000001110110011;
ROM[6688] <= 32'b00000000011100010010000000100011;
ROM[6689] <= 32'b00000000010000010000000100010011;
ROM[6690] <= 32'b00000000001100010010000000100011;
ROM[6691] <= 32'b00000000010000010000000100010011;
ROM[6692] <= 32'b00000000010000010010000000100011;
ROM[6693] <= 32'b00000000010000010000000100010011;
ROM[6694] <= 32'b00000000010100010010000000100011;
ROM[6695] <= 32'b00000000010000010000000100010011;
ROM[6696] <= 32'b00000000011000010010000000100011;
ROM[6697] <= 32'b00000000010000010000000100010011;
ROM[6698] <= 32'b00000001010000000000001110010011;
ROM[6699] <= 32'b00000000100000111000001110010011;
ROM[6700] <= 32'b01000000011100010000001110110011;
ROM[6701] <= 32'b00000000011100000000001000110011;
ROM[6702] <= 32'b00000000001000000000000110110011;
ROM[6703] <= 32'b01000000000000001011000011101111;
ROM[6704] <= 32'b11111111110000010000000100010011;
ROM[6705] <= 32'b00000000000000010010001110000011;
ROM[6706] <= 32'b00000000011101100010000000100011;
ROM[6707] <= 32'b00000001010000011010001110000011;
ROM[6708] <= 32'b00000000011100010010000000100011;
ROM[6709] <= 32'b00000000010000010000000100010011;
ROM[6710] <= 32'b00000110111100000000001110010011;
ROM[6711] <= 32'b00000000011100010010000000100011;
ROM[6712] <= 32'b00000000010000010000000100010011;
ROM[6713] <= 32'b00000000000000000111001110110111;
ROM[6714] <= 32'b10010011000000111000001110010011;
ROM[6715] <= 32'b00000000111000111000001110110011;
ROM[6716] <= 32'b00000000011100010010000000100011;
ROM[6717] <= 32'b00000000010000010000000100010011;
ROM[6718] <= 32'b00000000001100010010000000100011;
ROM[6719] <= 32'b00000000010000010000000100010011;
ROM[6720] <= 32'b00000000010000010010000000100011;
ROM[6721] <= 32'b00000000010000010000000100010011;
ROM[6722] <= 32'b00000000010100010010000000100011;
ROM[6723] <= 32'b00000000010000010000000100010011;
ROM[6724] <= 32'b00000000011000010010000000100011;
ROM[6725] <= 32'b00000000010000010000000100010011;
ROM[6726] <= 32'b00000001010000000000001110010011;
ROM[6727] <= 32'b00000000100000111000001110010011;
ROM[6728] <= 32'b01000000011100010000001110110011;
ROM[6729] <= 32'b00000000011100000000001000110011;
ROM[6730] <= 32'b00000000001000000000000110110011;
ROM[6731] <= 32'b00111001000000001011000011101111;
ROM[6732] <= 32'b11111111110000010000000100010011;
ROM[6733] <= 32'b00000000000000010010001110000011;
ROM[6734] <= 32'b00000000011101100010000000100011;
ROM[6735] <= 32'b00000001010000011010001110000011;
ROM[6736] <= 32'b00000000011100010010000000100011;
ROM[6737] <= 32'b00000000010000010000000100010011;
ROM[6738] <= 32'b00000010000000000000001110010011;
ROM[6739] <= 32'b00000000011100010010000000100011;
ROM[6740] <= 32'b00000000010000010000000100010011;
ROM[6741] <= 32'b00000000000000000111001110110111;
ROM[6742] <= 32'b10011010000000111000001110010011;
ROM[6743] <= 32'b00000000111000111000001110110011;
ROM[6744] <= 32'b00000000011100010010000000100011;
ROM[6745] <= 32'b00000000010000010000000100010011;
ROM[6746] <= 32'b00000000001100010010000000100011;
ROM[6747] <= 32'b00000000010000010000000100010011;
ROM[6748] <= 32'b00000000010000010010000000100011;
ROM[6749] <= 32'b00000000010000010000000100010011;
ROM[6750] <= 32'b00000000010100010010000000100011;
ROM[6751] <= 32'b00000000010000010000000100010011;
ROM[6752] <= 32'b00000000011000010010000000100011;
ROM[6753] <= 32'b00000000010000010000000100010011;
ROM[6754] <= 32'b00000001010000000000001110010011;
ROM[6755] <= 32'b00000000100000111000001110010011;
ROM[6756] <= 32'b01000000011100010000001110110011;
ROM[6757] <= 32'b00000000011100000000001000110011;
ROM[6758] <= 32'b00000000001000000000000110110011;
ROM[6759] <= 32'b00110010000000001011000011101111;
ROM[6760] <= 32'b11111111110000010000000100010011;
ROM[6761] <= 32'b00000000000000010010001110000011;
ROM[6762] <= 32'b00000000011101100010000000100011;
ROM[6763] <= 32'b00000001010000011010001110000011;
ROM[6764] <= 32'b00000000011100011010101000100011;
ROM[6765] <= 32'b00000000101100000000001110010011;
ROM[6766] <= 32'b00000000011100010010000000100011;
ROM[6767] <= 32'b00000000010000010000000100010011;
ROM[6768] <= 32'b00000000000000000111001110110111;
ROM[6769] <= 32'b10100000110000111000001110010011;
ROM[6770] <= 32'b00000000111000111000001110110011;
ROM[6771] <= 32'b00000000011100010010000000100011;
ROM[6772] <= 32'b00000000010000010000000100010011;
ROM[6773] <= 32'b00000000001100010010000000100011;
ROM[6774] <= 32'b00000000010000010000000100010011;
ROM[6775] <= 32'b00000000010000010010000000100011;
ROM[6776] <= 32'b00000000010000010000000100010011;
ROM[6777] <= 32'b00000000010100010010000000100011;
ROM[6778] <= 32'b00000000010000010000000100010011;
ROM[6779] <= 32'b00000000011000010010000000100011;
ROM[6780] <= 32'b00000000010000010000000100010011;
ROM[6781] <= 32'b00000001010000000000001110010011;
ROM[6782] <= 32'b00000000010000111000001110010011;
ROM[6783] <= 32'b01000000011100010000001110110011;
ROM[6784] <= 32'b00000000011100000000001000110011;
ROM[6785] <= 32'b00000000001000000000000110110011;
ROM[6786] <= 32'b01101111100100001010000011101111;
ROM[6787] <= 32'b11111111110000010000000100010011;
ROM[6788] <= 32'b00000000000000010010001110000011;
ROM[6789] <= 32'b00000000011100011010110000100011;
ROM[6790] <= 32'b00000001100000011010001110000011;
ROM[6791] <= 32'b00000000011100010010000000100011;
ROM[6792] <= 32'b00000000010000010000000100010011;
ROM[6793] <= 32'b00000010000000000000001110010011;
ROM[6794] <= 32'b00000000011100010010000000100011;
ROM[6795] <= 32'b00000000010000010000000100010011;
ROM[6796] <= 32'b00000000000000000111001110110111;
ROM[6797] <= 32'b10100111110000111000001110010011;
ROM[6798] <= 32'b00000000111000111000001110110011;
ROM[6799] <= 32'b00000000011100010010000000100011;
ROM[6800] <= 32'b00000000010000010000000100010011;
ROM[6801] <= 32'b00000000001100010010000000100011;
ROM[6802] <= 32'b00000000010000010000000100010011;
ROM[6803] <= 32'b00000000010000010010000000100011;
ROM[6804] <= 32'b00000000010000010000000100010011;
ROM[6805] <= 32'b00000000010100010010000000100011;
ROM[6806] <= 32'b00000000010000010000000100010011;
ROM[6807] <= 32'b00000000011000010010000000100011;
ROM[6808] <= 32'b00000000010000010000000100010011;
ROM[6809] <= 32'b00000001010000000000001110010011;
ROM[6810] <= 32'b00000000100000111000001110010011;
ROM[6811] <= 32'b01000000011100010000001110110011;
ROM[6812] <= 32'b00000000011100000000001000110011;
ROM[6813] <= 32'b00000000001000000000000110110011;
ROM[6814] <= 32'b00100100010000001011000011101111;
ROM[6815] <= 32'b11111111110000010000000100010011;
ROM[6816] <= 32'b00000000000000010010001110000011;
ROM[6817] <= 32'b00000000011101100010000000100011;
ROM[6818] <= 32'b00000001100000011010001110000011;
ROM[6819] <= 32'b00000000011100010010000000100011;
ROM[6820] <= 32'b00000000010000010000000100010011;
ROM[6821] <= 32'b00000111001100000000001110010011;
ROM[6822] <= 32'b00000000011100010010000000100011;
ROM[6823] <= 32'b00000000010000010000000100010011;
ROM[6824] <= 32'b00000000000000000111001110110111;
ROM[6825] <= 32'b10101110110000111000001110010011;
ROM[6826] <= 32'b00000000111000111000001110110011;
ROM[6827] <= 32'b00000000011100010010000000100011;
ROM[6828] <= 32'b00000000010000010000000100010011;
ROM[6829] <= 32'b00000000001100010010000000100011;
ROM[6830] <= 32'b00000000010000010000000100010011;
ROM[6831] <= 32'b00000000010000010010000000100011;
ROM[6832] <= 32'b00000000010000010000000100010011;
ROM[6833] <= 32'b00000000010100010010000000100011;
ROM[6834] <= 32'b00000000010000010000000100010011;
ROM[6835] <= 32'b00000000011000010010000000100011;
ROM[6836] <= 32'b00000000010000010000000100010011;
ROM[6837] <= 32'b00000001010000000000001110010011;
ROM[6838] <= 32'b00000000100000111000001110010011;
ROM[6839] <= 32'b01000000011100010000001110110011;
ROM[6840] <= 32'b00000000011100000000001000110011;
ROM[6841] <= 32'b00000000001000000000000110110011;
ROM[6842] <= 32'b00011101010000001011000011101111;
ROM[6843] <= 32'b11111111110000010000000100010011;
ROM[6844] <= 32'b00000000000000010010001110000011;
ROM[6845] <= 32'b00000000011101100010000000100011;
ROM[6846] <= 32'b00000001100000011010001110000011;
ROM[6847] <= 32'b00000000011100010010000000100011;
ROM[6848] <= 32'b00000000010000010000000100010011;
ROM[6849] <= 32'b00000110111000000000001110010011;
ROM[6850] <= 32'b00000000011100010010000000100011;
ROM[6851] <= 32'b00000000010000010000000100010011;
ROM[6852] <= 32'b00000000000000000111001110110111;
ROM[6853] <= 32'b10110101110000111000001110010011;
ROM[6854] <= 32'b00000000111000111000001110110011;
ROM[6855] <= 32'b00000000011100010010000000100011;
ROM[6856] <= 32'b00000000010000010000000100010011;
ROM[6857] <= 32'b00000000001100010010000000100011;
ROM[6858] <= 32'b00000000010000010000000100010011;
ROM[6859] <= 32'b00000000010000010010000000100011;
ROM[6860] <= 32'b00000000010000010000000100010011;
ROM[6861] <= 32'b00000000010100010010000000100011;
ROM[6862] <= 32'b00000000010000010000000100010011;
ROM[6863] <= 32'b00000000011000010010000000100011;
ROM[6864] <= 32'b00000000010000010000000100010011;
ROM[6865] <= 32'b00000001010000000000001110010011;
ROM[6866] <= 32'b00000000100000111000001110010011;
ROM[6867] <= 32'b01000000011100010000001110110011;
ROM[6868] <= 32'b00000000011100000000001000110011;
ROM[6869] <= 32'b00000000001000000000000110110011;
ROM[6870] <= 32'b00010110010000001011000011101111;
ROM[6871] <= 32'b11111111110000010000000100010011;
ROM[6872] <= 32'b00000000000000010010001110000011;
ROM[6873] <= 32'b00000000011101100010000000100011;
ROM[6874] <= 32'b00000001100000011010001110000011;
ROM[6875] <= 32'b00000000011100010010000000100011;
ROM[6876] <= 32'b00000000010000010000000100010011;
ROM[6877] <= 32'b00000110000100000000001110010011;
ROM[6878] <= 32'b00000000011100010010000000100011;
ROM[6879] <= 32'b00000000010000010000000100010011;
ROM[6880] <= 32'b00000000000000000111001110110111;
ROM[6881] <= 32'b10111100110000111000001110010011;
ROM[6882] <= 32'b00000000111000111000001110110011;
ROM[6883] <= 32'b00000000011100010010000000100011;
ROM[6884] <= 32'b00000000010000010000000100010011;
ROM[6885] <= 32'b00000000001100010010000000100011;
ROM[6886] <= 32'b00000000010000010000000100010011;
ROM[6887] <= 32'b00000000010000010010000000100011;
ROM[6888] <= 32'b00000000010000010000000100010011;
ROM[6889] <= 32'b00000000010100010010000000100011;
ROM[6890] <= 32'b00000000010000010000000100010011;
ROM[6891] <= 32'b00000000011000010010000000100011;
ROM[6892] <= 32'b00000000010000010000000100010011;
ROM[6893] <= 32'b00000001010000000000001110010011;
ROM[6894] <= 32'b00000000100000111000001110010011;
ROM[6895] <= 32'b01000000011100010000001110110011;
ROM[6896] <= 32'b00000000011100000000001000110011;
ROM[6897] <= 32'b00000000001000000000000110110011;
ROM[6898] <= 32'b00001111010000001011000011101111;
ROM[6899] <= 32'b11111111110000010000000100010011;
ROM[6900] <= 32'b00000000000000010010001110000011;
ROM[6901] <= 32'b00000000011101100010000000100011;
ROM[6902] <= 32'b00000001100000011010001110000011;
ROM[6903] <= 32'b00000000011100010010000000100011;
ROM[6904] <= 32'b00000000010000010000000100010011;
ROM[6905] <= 32'b00000110101100000000001110010011;
ROM[6906] <= 32'b00000000011100010010000000100011;
ROM[6907] <= 32'b00000000010000010000000100010011;
ROM[6908] <= 32'b00000000000000000111001110110111;
ROM[6909] <= 32'b11000011110000111000001110010011;
ROM[6910] <= 32'b00000000111000111000001110110011;
ROM[6911] <= 32'b00000000011100010010000000100011;
ROM[6912] <= 32'b00000000010000010000000100010011;
ROM[6913] <= 32'b00000000001100010010000000100011;
ROM[6914] <= 32'b00000000010000010000000100010011;
ROM[6915] <= 32'b00000000010000010010000000100011;
ROM[6916] <= 32'b00000000010000010000000100010011;
ROM[6917] <= 32'b00000000010100010010000000100011;
ROM[6918] <= 32'b00000000010000010000000100010011;
ROM[6919] <= 32'b00000000011000010010000000100011;
ROM[6920] <= 32'b00000000010000010000000100010011;
ROM[6921] <= 32'b00000001010000000000001110010011;
ROM[6922] <= 32'b00000000100000111000001110010011;
ROM[6923] <= 32'b01000000011100010000001110110011;
ROM[6924] <= 32'b00000000011100000000001000110011;
ROM[6925] <= 32'b00000000001000000000000110110011;
ROM[6926] <= 32'b00001000010000001011000011101111;
ROM[6927] <= 32'b11111111110000010000000100010011;
ROM[6928] <= 32'b00000000000000010010001110000011;
ROM[6929] <= 32'b00000000011101100010000000100011;
ROM[6930] <= 32'b00000001100000011010001110000011;
ROM[6931] <= 32'b00000000011100010010000000100011;
ROM[6932] <= 32'b00000000010000010000000100010011;
ROM[6933] <= 32'b00000110010100000000001110010011;
ROM[6934] <= 32'b00000000011100010010000000100011;
ROM[6935] <= 32'b00000000010000010000000100010011;
ROM[6936] <= 32'b00000000000000000111001110110111;
ROM[6937] <= 32'b11001010110000111000001110010011;
ROM[6938] <= 32'b00000000111000111000001110110011;
ROM[6939] <= 32'b00000000011100010010000000100011;
ROM[6940] <= 32'b00000000010000010000000100010011;
ROM[6941] <= 32'b00000000001100010010000000100011;
ROM[6942] <= 32'b00000000010000010000000100010011;
ROM[6943] <= 32'b00000000010000010010000000100011;
ROM[6944] <= 32'b00000000010000010000000100010011;
ROM[6945] <= 32'b00000000010100010010000000100011;
ROM[6946] <= 32'b00000000010000010000000100010011;
ROM[6947] <= 32'b00000000011000010010000000100011;
ROM[6948] <= 32'b00000000010000010000000100010011;
ROM[6949] <= 32'b00000001010000000000001110010011;
ROM[6950] <= 32'b00000000100000111000001110010011;
ROM[6951] <= 32'b01000000011100010000001110110011;
ROM[6952] <= 32'b00000000011100000000001000110011;
ROM[6953] <= 32'b00000000001000000000000110110011;
ROM[6954] <= 32'b00000001010000001011000011101111;
ROM[6955] <= 32'b11111111110000010000000100010011;
ROM[6956] <= 32'b00000000000000010010001110000011;
ROM[6957] <= 32'b00000000011101100010000000100011;
ROM[6958] <= 32'b00000001100000011010001110000011;
ROM[6959] <= 32'b00000000011100010010000000100011;
ROM[6960] <= 32'b00000000010000010000000100010011;
ROM[6961] <= 32'b00000110011100000000001110010011;
ROM[6962] <= 32'b00000000011100010010000000100011;
ROM[6963] <= 32'b00000000010000010000000100010011;
ROM[6964] <= 32'b00000000000000000111001110110111;
ROM[6965] <= 32'b11010001110000111000001110010011;
ROM[6966] <= 32'b00000000111000111000001110110011;
ROM[6967] <= 32'b00000000011100010010000000100011;
ROM[6968] <= 32'b00000000010000010000000100010011;
ROM[6969] <= 32'b00000000001100010010000000100011;
ROM[6970] <= 32'b00000000010000010000000100010011;
ROM[6971] <= 32'b00000000010000010010000000100011;
ROM[6972] <= 32'b00000000010000010000000100010011;
ROM[6973] <= 32'b00000000010100010010000000100011;
ROM[6974] <= 32'b00000000010000010000000100010011;
ROM[6975] <= 32'b00000000011000010010000000100011;
ROM[6976] <= 32'b00000000010000010000000100010011;
ROM[6977] <= 32'b00000001010000000000001110010011;
ROM[6978] <= 32'b00000000100000111000001110010011;
ROM[6979] <= 32'b01000000011100010000001110110011;
ROM[6980] <= 32'b00000000011100000000001000110011;
ROM[6981] <= 32'b00000000001000000000000110110011;
ROM[6982] <= 32'b01111010010100001010000011101111;
ROM[6983] <= 32'b11111111110000010000000100010011;
ROM[6984] <= 32'b00000000000000010010001110000011;
ROM[6985] <= 32'b00000000011101100010000000100011;
ROM[6986] <= 32'b00000001100000011010001110000011;
ROM[6987] <= 32'b00000000011100010010000000100011;
ROM[6988] <= 32'b00000000010000010000000100010011;
ROM[6989] <= 32'b00000110000100000000001110010011;
ROM[6990] <= 32'b00000000011100010010000000100011;
ROM[6991] <= 32'b00000000010000010000000100010011;
ROM[6992] <= 32'b00000000000000000111001110110111;
ROM[6993] <= 32'b11011000110000111000001110010011;
ROM[6994] <= 32'b00000000111000111000001110110011;
ROM[6995] <= 32'b00000000011100010010000000100011;
ROM[6996] <= 32'b00000000010000010000000100010011;
ROM[6997] <= 32'b00000000001100010010000000100011;
ROM[6998] <= 32'b00000000010000010000000100010011;
ROM[6999] <= 32'b00000000010000010010000000100011;
ROM[7000] <= 32'b00000000010000010000000100010011;
ROM[7001] <= 32'b00000000010100010010000000100011;
ROM[7002] <= 32'b00000000010000010000000100010011;
ROM[7003] <= 32'b00000000011000010010000000100011;
ROM[7004] <= 32'b00000000010000010000000100010011;
ROM[7005] <= 32'b00000001010000000000001110010011;
ROM[7006] <= 32'b00000000100000111000001110010011;
ROM[7007] <= 32'b01000000011100010000001110110011;
ROM[7008] <= 32'b00000000011100000000001000110011;
ROM[7009] <= 32'b00000000001000000000000110110011;
ROM[7010] <= 32'b01110011010100001010000011101111;
ROM[7011] <= 32'b11111111110000010000000100010011;
ROM[7012] <= 32'b00000000000000010010001110000011;
ROM[7013] <= 32'b00000000011101100010000000100011;
ROM[7014] <= 32'b00000001100000011010001110000011;
ROM[7015] <= 32'b00000000011100010010000000100011;
ROM[7016] <= 32'b00000000010000010000000100010011;
ROM[7017] <= 32'b00000110110100000000001110010011;
ROM[7018] <= 32'b00000000011100010010000000100011;
ROM[7019] <= 32'b00000000010000010000000100010011;
ROM[7020] <= 32'b00000000000000000111001110110111;
ROM[7021] <= 32'b11011111110000111000001110010011;
ROM[7022] <= 32'b00000000111000111000001110110011;
ROM[7023] <= 32'b00000000011100010010000000100011;
ROM[7024] <= 32'b00000000010000010000000100010011;
ROM[7025] <= 32'b00000000001100010010000000100011;
ROM[7026] <= 32'b00000000010000010000000100010011;
ROM[7027] <= 32'b00000000010000010010000000100011;
ROM[7028] <= 32'b00000000010000010000000100010011;
ROM[7029] <= 32'b00000000010100010010000000100011;
ROM[7030] <= 32'b00000000010000010000000100010011;
ROM[7031] <= 32'b00000000011000010010000000100011;
ROM[7032] <= 32'b00000000010000010000000100010011;
ROM[7033] <= 32'b00000001010000000000001110010011;
ROM[7034] <= 32'b00000000100000111000001110010011;
ROM[7035] <= 32'b01000000011100010000001110110011;
ROM[7036] <= 32'b00000000011100000000001000110011;
ROM[7037] <= 32'b00000000001000000000000110110011;
ROM[7038] <= 32'b01101100010100001010000011101111;
ROM[7039] <= 32'b11111111110000010000000100010011;
ROM[7040] <= 32'b00000000000000010010001110000011;
ROM[7041] <= 32'b00000000011101100010000000100011;
ROM[7042] <= 32'b00000001100000011010001110000011;
ROM[7043] <= 32'b00000000011100010010000000100011;
ROM[7044] <= 32'b00000000010000010000000100010011;
ROM[7045] <= 32'b00000110010100000000001110010011;
ROM[7046] <= 32'b00000000011100010010000000100011;
ROM[7047] <= 32'b00000000010000010000000100010011;
ROM[7048] <= 32'b00000000000000000111001110110111;
ROM[7049] <= 32'b11100110110000111000001110010011;
ROM[7050] <= 32'b00000000111000111000001110110011;
ROM[7051] <= 32'b00000000011100010010000000100011;
ROM[7052] <= 32'b00000000010000010000000100010011;
ROM[7053] <= 32'b00000000001100010010000000100011;
ROM[7054] <= 32'b00000000010000010000000100010011;
ROM[7055] <= 32'b00000000010000010010000000100011;
ROM[7056] <= 32'b00000000010000010000000100010011;
ROM[7057] <= 32'b00000000010100010010000000100011;
ROM[7058] <= 32'b00000000010000010000000100010011;
ROM[7059] <= 32'b00000000011000010010000000100011;
ROM[7060] <= 32'b00000000010000010000000100010011;
ROM[7061] <= 32'b00000001010000000000001110010011;
ROM[7062] <= 32'b00000000100000111000001110010011;
ROM[7063] <= 32'b01000000011100010000001110110011;
ROM[7064] <= 32'b00000000011100000000001000110011;
ROM[7065] <= 32'b00000000001000000000000110110011;
ROM[7066] <= 32'b01100101010100001010000011101111;
ROM[7067] <= 32'b11111111110000010000000100010011;
ROM[7068] <= 32'b00000000000000010010001110000011;
ROM[7069] <= 32'b00000000011101100010000000100011;
ROM[7070] <= 32'b00000001100000011010001110000011;
ROM[7071] <= 32'b00000000011100010010000000100011;
ROM[7072] <= 32'b00000000010000010000000100010011;
ROM[7073] <= 32'b00000010000000000000001110010011;
ROM[7074] <= 32'b00000000011100010010000000100011;
ROM[7075] <= 32'b00000000010000010000000100010011;
ROM[7076] <= 32'b00000000000000000111001110110111;
ROM[7077] <= 32'b11101101110000111000001110010011;
ROM[7078] <= 32'b00000000111000111000001110110011;
ROM[7079] <= 32'b00000000011100010010000000100011;
ROM[7080] <= 32'b00000000010000010000000100010011;
ROM[7081] <= 32'b00000000001100010010000000100011;
ROM[7082] <= 32'b00000000010000010000000100010011;
ROM[7083] <= 32'b00000000010000010010000000100011;
ROM[7084] <= 32'b00000000010000010000000100010011;
ROM[7085] <= 32'b00000000010100010010000000100011;
ROM[7086] <= 32'b00000000010000010000000100010011;
ROM[7087] <= 32'b00000000011000010010000000100011;
ROM[7088] <= 32'b00000000010000010000000100010011;
ROM[7089] <= 32'b00000001010000000000001110010011;
ROM[7090] <= 32'b00000000100000111000001110010011;
ROM[7091] <= 32'b01000000011100010000001110110011;
ROM[7092] <= 32'b00000000011100000000001000110011;
ROM[7093] <= 32'b00000000001000000000000110110011;
ROM[7094] <= 32'b01011110010100001010000011101111;
ROM[7095] <= 32'b11111111110000010000000100010011;
ROM[7096] <= 32'b00000000000000010010001110000011;
ROM[7097] <= 32'b00000000011101100010000000100011;
ROM[7098] <= 32'b00000001100000011010001110000011;
ROM[7099] <= 32'b00000000011100011010110000100011;
ROM[7100] <= 32'b00000000011100000000001110010011;
ROM[7101] <= 32'b00000000011100010010000000100011;
ROM[7102] <= 32'b00000000010000010000000100010011;
ROM[7103] <= 32'b00000000000000000111001110110111;
ROM[7104] <= 32'b11110100100000111000001110010011;
ROM[7105] <= 32'b00000000111000111000001110110011;
ROM[7106] <= 32'b00000000011100010010000000100011;
ROM[7107] <= 32'b00000000010000010000000100010011;
ROM[7108] <= 32'b00000000001100010010000000100011;
ROM[7109] <= 32'b00000000010000010000000100010011;
ROM[7110] <= 32'b00000000010000010010000000100011;
ROM[7111] <= 32'b00000000010000010000000100010011;
ROM[7112] <= 32'b00000000010100010010000000100011;
ROM[7113] <= 32'b00000000010000010000000100010011;
ROM[7114] <= 32'b00000000011000010010000000100011;
ROM[7115] <= 32'b00000000010000010000000100010011;
ROM[7116] <= 32'b00000001010000000000001110010011;
ROM[7117] <= 32'b00000000010000111000001110010011;
ROM[7118] <= 32'b01000000011100010000001110110011;
ROM[7119] <= 32'b00000000011100000000001000110011;
ROM[7120] <= 32'b00000000001000000000000110110011;
ROM[7121] <= 32'b00011011110100001010000011101111;
ROM[7122] <= 32'b11111111110000010000000100010011;
ROM[7123] <= 32'b00000000000000010010001110000011;
ROM[7124] <= 32'b00000000011100011010111000100011;
ROM[7125] <= 32'b00000001110000011010001110000011;
ROM[7126] <= 32'b00000000011100010010000000100011;
ROM[7127] <= 32'b00000000010000010000000100010011;
ROM[7128] <= 32'b00000010000000000000001110010011;
ROM[7129] <= 32'b00000000011100010010000000100011;
ROM[7130] <= 32'b00000000010000010000000100010011;
ROM[7131] <= 32'b00000000000000000111001110110111;
ROM[7132] <= 32'b11111011100000111000001110010011;
ROM[7133] <= 32'b00000000111000111000001110110011;
ROM[7134] <= 32'b00000000011100010010000000100011;
ROM[7135] <= 32'b00000000010000010000000100010011;
ROM[7136] <= 32'b00000000001100010010000000100011;
ROM[7137] <= 32'b00000000010000010000000100010011;
ROM[7138] <= 32'b00000000010000010010000000100011;
ROM[7139] <= 32'b00000000010000010000000100010011;
ROM[7140] <= 32'b00000000010100010010000000100011;
ROM[7141] <= 32'b00000000010000010000000100010011;
ROM[7142] <= 32'b00000000011000010010000000100011;
ROM[7143] <= 32'b00000000010000010000000100010011;
ROM[7144] <= 32'b00000001010000000000001110010011;
ROM[7145] <= 32'b00000000100000111000001110010011;
ROM[7146] <= 32'b01000000011100010000001110110011;
ROM[7147] <= 32'b00000000011100000000001000110011;
ROM[7148] <= 32'b00000000001000000000000110110011;
ROM[7149] <= 32'b01010000100100001010000011101111;
ROM[7150] <= 32'b11111111110000010000000100010011;
ROM[7151] <= 32'b00000000000000010010001110000011;
ROM[7152] <= 32'b00000000011101100010000000100011;
ROM[7153] <= 32'b00000001110000011010001110000011;
ROM[7154] <= 32'b00000000011100010010000000100011;
ROM[7155] <= 32'b00000000010000010000000100010011;
ROM[7156] <= 32'b00000111000100000000001110010011;
ROM[7157] <= 32'b00000000011100010010000000100011;
ROM[7158] <= 32'b00000000010000010000000100010011;
ROM[7159] <= 32'b00000000000000000111001110110111;
ROM[7160] <= 32'b00000010100000111000001110010011;
ROM[7161] <= 32'b00000000111000111000001110110011;
ROM[7162] <= 32'b00000000011100010010000000100011;
ROM[7163] <= 32'b00000000010000010000000100010011;
ROM[7164] <= 32'b00000000001100010010000000100011;
ROM[7165] <= 32'b00000000010000010000000100010011;
ROM[7166] <= 32'b00000000010000010010000000100011;
ROM[7167] <= 32'b00000000010000010000000100010011;
ROM[7168] <= 32'b00000000010100010010000000100011;
ROM[7169] <= 32'b00000000010000010000000100010011;
ROM[7170] <= 32'b00000000011000010010000000100011;
ROM[7171] <= 32'b00000000010000010000000100010011;
ROM[7172] <= 32'b00000001010000000000001110010011;
ROM[7173] <= 32'b00000000100000111000001110010011;
ROM[7174] <= 32'b01000000011100010000001110110011;
ROM[7175] <= 32'b00000000011100000000001000110011;
ROM[7176] <= 32'b00000000001000000000000110110011;
ROM[7177] <= 32'b01001001100100001010000011101111;
ROM[7178] <= 32'b11111111110000010000000100010011;
ROM[7179] <= 32'b00000000000000010010001110000011;
ROM[7180] <= 32'b00000000011101100010000000100011;
ROM[7181] <= 32'b00000001110000011010001110000011;
ROM[7182] <= 32'b00000000011100010010000000100011;
ROM[7183] <= 32'b00000000010000010000000100010011;
ROM[7184] <= 32'b00000111001100000000001110010011;
ROM[7185] <= 32'b00000000011100010010000000100011;
ROM[7186] <= 32'b00000000010000010000000100010011;
ROM[7187] <= 32'b00000000000000000111001110110111;
ROM[7188] <= 32'b00001001100000111000001110010011;
ROM[7189] <= 32'b00000000111000111000001110110011;
ROM[7190] <= 32'b00000000011100010010000000100011;
ROM[7191] <= 32'b00000000010000010000000100010011;
ROM[7192] <= 32'b00000000001100010010000000100011;
ROM[7193] <= 32'b00000000010000010000000100010011;
ROM[7194] <= 32'b00000000010000010010000000100011;
ROM[7195] <= 32'b00000000010000010000000100010011;
ROM[7196] <= 32'b00000000010100010010000000100011;
ROM[7197] <= 32'b00000000010000010000000100010011;
ROM[7198] <= 32'b00000000011000010010000000100011;
ROM[7199] <= 32'b00000000010000010000000100010011;
ROM[7200] <= 32'b00000001010000000000001110010011;
ROM[7201] <= 32'b00000000100000111000001110010011;
ROM[7202] <= 32'b01000000011100010000001110110011;
ROM[7203] <= 32'b00000000011100000000001000110011;
ROM[7204] <= 32'b00000000001000000000000110110011;
ROM[7205] <= 32'b01000010100100001010000011101111;
ROM[7206] <= 32'b11111111110000010000000100010011;
ROM[7207] <= 32'b00000000000000010010001110000011;
ROM[7208] <= 32'b00000000011101100010000000100011;
ROM[7209] <= 32'b00000001110000011010001110000011;
ROM[7210] <= 32'b00000000011100010010000000100011;
ROM[7211] <= 32'b00000000010000010000000100010011;
ROM[7212] <= 32'b00000110111100000000001110010011;
ROM[7213] <= 32'b00000000011100010010000000100011;
ROM[7214] <= 32'b00000000010000010000000100010011;
ROM[7215] <= 32'b00000000000000000111001110110111;
ROM[7216] <= 32'b00010000100000111000001110010011;
ROM[7217] <= 32'b00000000111000111000001110110011;
ROM[7218] <= 32'b00000000011100010010000000100011;
ROM[7219] <= 32'b00000000010000010000000100010011;
ROM[7220] <= 32'b00000000001100010010000000100011;
ROM[7221] <= 32'b00000000010000010000000100010011;
ROM[7222] <= 32'b00000000010000010010000000100011;
ROM[7223] <= 32'b00000000010000010000000100010011;
ROM[7224] <= 32'b00000000010100010010000000100011;
ROM[7225] <= 32'b00000000010000010000000100010011;
ROM[7226] <= 32'b00000000011000010010000000100011;
ROM[7227] <= 32'b00000000010000010000000100010011;
ROM[7228] <= 32'b00000001010000000000001110010011;
ROM[7229] <= 32'b00000000100000111000001110010011;
ROM[7230] <= 32'b01000000011100010000001110110011;
ROM[7231] <= 32'b00000000011100000000001000110011;
ROM[7232] <= 32'b00000000001000000000000110110011;
ROM[7233] <= 32'b00111011100100001010000011101111;
ROM[7234] <= 32'b11111111110000010000000100010011;
ROM[7235] <= 32'b00000000000000010010001110000011;
ROM[7236] <= 32'b00000000011101100010000000100011;
ROM[7237] <= 32'b00000001110000011010001110000011;
ROM[7238] <= 32'b00000000011100010010000000100011;
ROM[7239] <= 32'b00000000010000010000000100010011;
ROM[7240] <= 32'b00000111001000000000001110010011;
ROM[7241] <= 32'b00000000011100010010000000100011;
ROM[7242] <= 32'b00000000010000010000000100010011;
ROM[7243] <= 32'b00000000000000000111001110110111;
ROM[7244] <= 32'b00010111100000111000001110010011;
ROM[7245] <= 32'b00000000111000111000001110110011;
ROM[7246] <= 32'b00000000011100010010000000100011;
ROM[7247] <= 32'b00000000010000010000000100010011;
ROM[7248] <= 32'b00000000001100010010000000100011;
ROM[7249] <= 32'b00000000010000010000000100010011;
ROM[7250] <= 32'b00000000010000010010000000100011;
ROM[7251] <= 32'b00000000010000010000000100010011;
ROM[7252] <= 32'b00000000010100010010000000100011;
ROM[7253] <= 32'b00000000010000010000000100010011;
ROM[7254] <= 32'b00000000011000010010000000100011;
ROM[7255] <= 32'b00000000010000010000000100010011;
ROM[7256] <= 32'b00000001010000000000001110010011;
ROM[7257] <= 32'b00000000100000111000001110010011;
ROM[7258] <= 32'b01000000011100010000001110110011;
ROM[7259] <= 32'b00000000011100000000001000110011;
ROM[7260] <= 32'b00000000001000000000000110110011;
ROM[7261] <= 32'b00110100100100001010000011101111;
ROM[7262] <= 32'b11111111110000010000000100010011;
ROM[7263] <= 32'b00000000000000010010001110000011;
ROM[7264] <= 32'b00000000011101100010000000100011;
ROM[7265] <= 32'b00000001110000011010001110000011;
ROM[7266] <= 32'b00000000011100010010000000100011;
ROM[7267] <= 32'b00000000010000010000000100010011;
ROM[7268] <= 32'b00000111010000000000001110010011;
ROM[7269] <= 32'b00000000011100010010000000100011;
ROM[7270] <= 32'b00000000010000010000000100010011;
ROM[7271] <= 32'b00000000000000000111001110110111;
ROM[7272] <= 32'b00011110100000111000001110010011;
ROM[7273] <= 32'b00000000111000111000001110110011;
ROM[7274] <= 32'b00000000011100010010000000100011;
ROM[7275] <= 32'b00000000010000010000000100010011;
ROM[7276] <= 32'b00000000001100010010000000100011;
ROM[7277] <= 32'b00000000010000010000000100010011;
ROM[7278] <= 32'b00000000010000010010000000100011;
ROM[7279] <= 32'b00000000010000010000000100010011;
ROM[7280] <= 32'b00000000010100010010000000100011;
ROM[7281] <= 32'b00000000010000010000000100010011;
ROM[7282] <= 32'b00000000011000010010000000100011;
ROM[7283] <= 32'b00000000010000010000000100010011;
ROM[7284] <= 32'b00000001010000000000001110010011;
ROM[7285] <= 32'b00000000100000111000001110010011;
ROM[7286] <= 32'b01000000011100010000001110110011;
ROM[7287] <= 32'b00000000011100000000001000110011;
ROM[7288] <= 32'b00000000001000000000000110110011;
ROM[7289] <= 32'b00101101100100001010000011101111;
ROM[7290] <= 32'b11111111110000010000000100010011;
ROM[7291] <= 32'b00000000000000010010001110000011;
ROM[7292] <= 32'b00000000011101100010000000100011;
ROM[7293] <= 32'b00000001110000011010001110000011;
ROM[7294] <= 32'b00000000011100010010000000100011;
ROM[7295] <= 32'b00000000010000010000000100010011;
ROM[7296] <= 32'b00000010000000000000001110010011;
ROM[7297] <= 32'b00000000011100010010000000100011;
ROM[7298] <= 32'b00000000010000010000000100010011;
ROM[7299] <= 32'b00000000000000000111001110110111;
ROM[7300] <= 32'b00100101100000111000001110010011;
ROM[7301] <= 32'b00000000111000111000001110110011;
ROM[7302] <= 32'b00000000011100010010000000100011;
ROM[7303] <= 32'b00000000010000010000000100010011;
ROM[7304] <= 32'b00000000001100010010000000100011;
ROM[7305] <= 32'b00000000010000010000000100010011;
ROM[7306] <= 32'b00000000010000010010000000100011;
ROM[7307] <= 32'b00000000010000010000000100010011;
ROM[7308] <= 32'b00000000010100010010000000100011;
ROM[7309] <= 32'b00000000010000010000000100010011;
ROM[7310] <= 32'b00000000011000010010000000100011;
ROM[7311] <= 32'b00000000010000010000000100010011;
ROM[7312] <= 32'b00000001010000000000001110010011;
ROM[7313] <= 32'b00000000100000111000001110010011;
ROM[7314] <= 32'b01000000011100010000001110110011;
ROM[7315] <= 32'b00000000011100000000001000110011;
ROM[7316] <= 32'b00000000001000000000000110110011;
ROM[7317] <= 32'b00100110100100001010000011101111;
ROM[7318] <= 32'b11111111110000010000000100010011;
ROM[7319] <= 32'b00000000000000010010001110000011;
ROM[7320] <= 32'b00000000011101100010000000100011;
ROM[7321] <= 32'b00000001110000011010001110000011;
ROM[7322] <= 32'b00000000011100011010111000100011;
ROM[7323] <= 32'b00000000100100000000001110010011;
ROM[7324] <= 32'b00000000011100010010000000100011;
ROM[7325] <= 32'b00000000010000010000000100010011;
ROM[7326] <= 32'b00000000000000000111001110110111;
ROM[7327] <= 32'b00101100010000111000001110010011;
ROM[7328] <= 32'b00000000111000111000001110110011;
ROM[7329] <= 32'b00000000011100010010000000100011;
ROM[7330] <= 32'b00000000010000010000000100010011;
ROM[7331] <= 32'b00000000001100010010000000100011;
ROM[7332] <= 32'b00000000010000010000000100010011;
ROM[7333] <= 32'b00000000010000010010000000100011;
ROM[7334] <= 32'b00000000010000010000000100010011;
ROM[7335] <= 32'b00000000010100010010000000100011;
ROM[7336] <= 32'b00000000010000010000000100010011;
ROM[7337] <= 32'b00000000011000010010000000100011;
ROM[7338] <= 32'b00000000010000010000000100010011;
ROM[7339] <= 32'b00000001010000000000001110010011;
ROM[7340] <= 32'b00000000010000111000001110010011;
ROM[7341] <= 32'b01000000011100010000001110110011;
ROM[7342] <= 32'b00000000011100000000001000110011;
ROM[7343] <= 32'b00000000001000000000000110110011;
ROM[7344] <= 32'b01100100000000001010000011101111;
ROM[7345] <= 32'b11111111110000010000000100010011;
ROM[7346] <= 32'b00000000000000010010001110000011;
ROM[7347] <= 32'b00000010011100011010000000100011;
ROM[7348] <= 32'b00000010000000011010001110000011;
ROM[7349] <= 32'b00000000011100010010000000100011;
ROM[7350] <= 32'b00000000010000010000000100010011;
ROM[7351] <= 32'b00000010000000000000001110010011;
ROM[7352] <= 32'b00000000011100010010000000100011;
ROM[7353] <= 32'b00000000010000010000000100010011;
ROM[7354] <= 32'b00000000000000000111001110110111;
ROM[7355] <= 32'b00110011010000111000001110010011;
ROM[7356] <= 32'b00000000111000111000001110110011;
ROM[7357] <= 32'b00000000011100010010000000100011;
ROM[7358] <= 32'b00000000010000010000000100010011;
ROM[7359] <= 32'b00000000001100010010000000100011;
ROM[7360] <= 32'b00000000010000010000000100010011;
ROM[7361] <= 32'b00000000010000010010000000100011;
ROM[7362] <= 32'b00000000010000010000000100010011;
ROM[7363] <= 32'b00000000010100010010000000100011;
ROM[7364] <= 32'b00000000010000010000000100010011;
ROM[7365] <= 32'b00000000011000010010000000100011;
ROM[7366] <= 32'b00000000010000010000000100010011;
ROM[7367] <= 32'b00000001010000000000001110010011;
ROM[7368] <= 32'b00000000100000111000001110010011;
ROM[7369] <= 32'b01000000011100010000001110110011;
ROM[7370] <= 32'b00000000011100000000001000110011;
ROM[7371] <= 32'b00000000001000000000000110110011;
ROM[7372] <= 32'b00011000110100001010000011101111;
ROM[7373] <= 32'b11111111110000010000000100010011;
ROM[7374] <= 32'b00000000000000010010001110000011;
ROM[7375] <= 32'b00000000011101100010000000100011;
ROM[7376] <= 32'b00000010000000011010001110000011;
ROM[7377] <= 32'b00000000011100010010000000100011;
ROM[7378] <= 32'b00000000010000010000000100010011;
ROM[7379] <= 32'b00000110100000000000001110010011;
ROM[7380] <= 32'b00000000011100010010000000100011;
ROM[7381] <= 32'b00000000010000010000000100010011;
ROM[7382] <= 32'b00000000000000000111001110110111;
ROM[7383] <= 32'b00111010010000111000001110010011;
ROM[7384] <= 32'b00000000111000111000001110110011;
ROM[7385] <= 32'b00000000011100010010000000100011;
ROM[7386] <= 32'b00000000010000010000000100010011;
ROM[7387] <= 32'b00000000001100010010000000100011;
ROM[7388] <= 32'b00000000010000010000000100010011;
ROM[7389] <= 32'b00000000010000010010000000100011;
ROM[7390] <= 32'b00000000010000010000000100010011;
ROM[7391] <= 32'b00000000010100010010000000100011;
ROM[7392] <= 32'b00000000010000010000000100010011;
ROM[7393] <= 32'b00000000011000010010000000100011;
ROM[7394] <= 32'b00000000010000010000000100010011;
ROM[7395] <= 32'b00000001010000000000001110010011;
ROM[7396] <= 32'b00000000100000111000001110010011;
ROM[7397] <= 32'b01000000011100010000001110110011;
ROM[7398] <= 32'b00000000011100000000001000110011;
ROM[7399] <= 32'b00000000001000000000000110110011;
ROM[7400] <= 32'b00010001110100001010000011101111;
ROM[7401] <= 32'b11111111110000010000000100010011;
ROM[7402] <= 32'b00000000000000010010001110000011;
ROM[7403] <= 32'b00000000011101100010000000100011;
ROM[7404] <= 32'b00000010000000011010001110000011;
ROM[7405] <= 32'b00000000011100010010000000100011;
ROM[7406] <= 32'b00000000010000010000000100010011;
ROM[7407] <= 32'b00000110000100000000001110010011;
ROM[7408] <= 32'b00000000011100010010000000100011;
ROM[7409] <= 32'b00000000010000010000000100010011;
ROM[7410] <= 32'b00000000000000000111001110110111;
ROM[7411] <= 32'b01000001010000111000001110010011;
ROM[7412] <= 32'b00000000111000111000001110110011;
ROM[7413] <= 32'b00000000011100010010000000100011;
ROM[7414] <= 32'b00000000010000010000000100010011;
ROM[7415] <= 32'b00000000001100010010000000100011;
ROM[7416] <= 32'b00000000010000010000000100010011;
ROM[7417] <= 32'b00000000010000010010000000100011;
ROM[7418] <= 32'b00000000010000010000000100010011;
ROM[7419] <= 32'b00000000010100010010000000100011;
ROM[7420] <= 32'b00000000010000010000000100010011;
ROM[7421] <= 32'b00000000011000010010000000100011;
ROM[7422] <= 32'b00000000010000010000000100010011;
ROM[7423] <= 32'b00000001010000000000001110010011;
ROM[7424] <= 32'b00000000100000111000001110010011;
ROM[7425] <= 32'b01000000011100010000001110110011;
ROM[7426] <= 32'b00000000011100000000001000110011;
ROM[7427] <= 32'b00000000001000000000000110110011;
ROM[7428] <= 32'b00001010110100001010000011101111;
ROM[7429] <= 32'b11111111110000010000000100010011;
ROM[7430] <= 32'b00000000000000010010001110000011;
ROM[7431] <= 32'b00000000011101100010000000100011;
ROM[7432] <= 32'b00000010000000011010001110000011;
ROM[7433] <= 32'b00000000011100010010000000100011;
ROM[7434] <= 32'b00000000010000010000000100010011;
ROM[7435] <= 32'b00000110111000000000001110010011;
ROM[7436] <= 32'b00000000011100010010000000100011;
ROM[7437] <= 32'b00000000010000010000000100010011;
ROM[7438] <= 32'b00000000000000000111001110110111;
ROM[7439] <= 32'b01001000010000111000001110010011;
ROM[7440] <= 32'b00000000111000111000001110110011;
ROM[7441] <= 32'b00000000011100010010000000100011;
ROM[7442] <= 32'b00000000010000010000000100010011;
ROM[7443] <= 32'b00000000001100010010000000100011;
ROM[7444] <= 32'b00000000010000010000000100010011;
ROM[7445] <= 32'b00000000010000010010000000100011;
ROM[7446] <= 32'b00000000010000010000000100010011;
ROM[7447] <= 32'b00000000010100010010000000100011;
ROM[7448] <= 32'b00000000010000010000000100010011;
ROM[7449] <= 32'b00000000011000010010000000100011;
ROM[7450] <= 32'b00000000010000010000000100010011;
ROM[7451] <= 32'b00000001010000000000001110010011;
ROM[7452] <= 32'b00000000100000111000001110010011;
ROM[7453] <= 32'b01000000011100010000001110110011;
ROM[7454] <= 32'b00000000011100000000001000110011;
ROM[7455] <= 32'b00000000001000000000000110110011;
ROM[7456] <= 32'b00000011110100001010000011101111;
ROM[7457] <= 32'b11111111110000010000000100010011;
ROM[7458] <= 32'b00000000000000010010001110000011;
ROM[7459] <= 32'b00000000011101100010000000100011;
ROM[7460] <= 32'b00000010000000011010001110000011;
ROM[7461] <= 32'b00000000011100010010000000100011;
ROM[7462] <= 32'b00000000010000010000000100010011;
ROM[7463] <= 32'b00000110011100000000001110010011;
ROM[7464] <= 32'b00000000011100010010000000100011;
ROM[7465] <= 32'b00000000010000010000000100010011;
ROM[7466] <= 32'b00000000000000000111001110110111;
ROM[7467] <= 32'b01001111010000111000001110010011;
ROM[7468] <= 32'b00000000111000111000001110110011;
ROM[7469] <= 32'b00000000011100010010000000100011;
ROM[7470] <= 32'b00000000010000010000000100010011;
ROM[7471] <= 32'b00000000001100010010000000100011;
ROM[7472] <= 32'b00000000010000010000000100010011;
ROM[7473] <= 32'b00000000010000010010000000100011;
ROM[7474] <= 32'b00000000010000010000000100010011;
ROM[7475] <= 32'b00000000010100010010000000100011;
ROM[7476] <= 32'b00000000010000010000000100010011;
ROM[7477] <= 32'b00000000011000010010000000100011;
ROM[7478] <= 32'b00000000010000010000000100010011;
ROM[7479] <= 32'b00000001010000000000001110010011;
ROM[7480] <= 32'b00000000100000111000001110010011;
ROM[7481] <= 32'b01000000011100010000001110110011;
ROM[7482] <= 32'b00000000011100000000001000110011;
ROM[7483] <= 32'b00000000001000000000000110110011;
ROM[7484] <= 32'b01111100110000001010000011101111;
ROM[7485] <= 32'b11111111110000010000000100010011;
ROM[7486] <= 32'b00000000000000010010001110000011;
ROM[7487] <= 32'b00000000011101100010000000100011;
ROM[7488] <= 32'b00000010000000011010001110000011;
ROM[7489] <= 32'b00000000011100010010000000100011;
ROM[7490] <= 32'b00000000010000010000000100010011;
ROM[7491] <= 32'b00000110110100000000001110010011;
ROM[7492] <= 32'b00000000011100010010000000100011;
ROM[7493] <= 32'b00000000010000010000000100010011;
ROM[7494] <= 32'b00000000000000000111001110110111;
ROM[7495] <= 32'b01010110010000111000001110010011;
ROM[7496] <= 32'b00000000111000111000001110110011;
ROM[7497] <= 32'b00000000011100010010000000100011;
ROM[7498] <= 32'b00000000010000010000000100010011;
ROM[7499] <= 32'b00000000001100010010000000100011;
ROM[7500] <= 32'b00000000010000010000000100010011;
ROM[7501] <= 32'b00000000010000010010000000100011;
ROM[7502] <= 32'b00000000010000010000000100010011;
ROM[7503] <= 32'b00000000010100010010000000100011;
ROM[7504] <= 32'b00000000010000010000000100010011;
ROM[7505] <= 32'b00000000011000010010000000100011;
ROM[7506] <= 32'b00000000010000010000000100010011;
ROM[7507] <= 32'b00000001010000000000001110010011;
ROM[7508] <= 32'b00000000100000111000001110010011;
ROM[7509] <= 32'b01000000011100010000001110110011;
ROM[7510] <= 32'b00000000011100000000001000110011;
ROM[7511] <= 32'b00000000001000000000000110110011;
ROM[7512] <= 32'b01110101110000001010000011101111;
ROM[7513] <= 32'b11111111110000010000000100010011;
ROM[7514] <= 32'b00000000000000010010001110000011;
ROM[7515] <= 32'b00000000011101100010000000100011;
ROM[7516] <= 32'b00000010000000011010001110000011;
ROM[7517] <= 32'b00000000011100010010000000100011;
ROM[7518] <= 32'b00000000010000010000000100010011;
ROM[7519] <= 32'b00000110000100000000001110010011;
ROM[7520] <= 32'b00000000011100010010000000100011;
ROM[7521] <= 32'b00000000010000010000000100010011;
ROM[7522] <= 32'b00000000000000000111001110110111;
ROM[7523] <= 32'b01011101010000111000001110010011;
ROM[7524] <= 32'b00000000111000111000001110110011;
ROM[7525] <= 32'b00000000011100010010000000100011;
ROM[7526] <= 32'b00000000010000010000000100010011;
ROM[7527] <= 32'b00000000001100010010000000100011;
ROM[7528] <= 32'b00000000010000010000000100010011;
ROM[7529] <= 32'b00000000010000010010000000100011;
ROM[7530] <= 32'b00000000010000010000000100010011;
ROM[7531] <= 32'b00000000010100010010000000100011;
ROM[7532] <= 32'b00000000010000010000000100010011;
ROM[7533] <= 32'b00000000011000010010000000100011;
ROM[7534] <= 32'b00000000010000010000000100010011;
ROM[7535] <= 32'b00000001010000000000001110010011;
ROM[7536] <= 32'b00000000100000111000001110010011;
ROM[7537] <= 32'b01000000011100010000001110110011;
ROM[7538] <= 32'b00000000011100000000001000110011;
ROM[7539] <= 32'b00000000001000000000000110110011;
ROM[7540] <= 32'b01101110110000001010000011101111;
ROM[7541] <= 32'b11111111110000010000000100010011;
ROM[7542] <= 32'b00000000000000010010001110000011;
ROM[7543] <= 32'b00000000011101100010000000100011;
ROM[7544] <= 32'b00000010000000011010001110000011;
ROM[7545] <= 32'b00000000011100010010000000100011;
ROM[7546] <= 32'b00000000010000010000000100010011;
ROM[7547] <= 32'b00000110111000000000001110010011;
ROM[7548] <= 32'b00000000011100010010000000100011;
ROM[7549] <= 32'b00000000010000010000000100010011;
ROM[7550] <= 32'b00000000000000000111001110110111;
ROM[7551] <= 32'b01100100010000111000001110010011;
ROM[7552] <= 32'b00000000111000111000001110110011;
ROM[7553] <= 32'b00000000011100010010000000100011;
ROM[7554] <= 32'b00000000010000010000000100010011;
ROM[7555] <= 32'b00000000001100010010000000100011;
ROM[7556] <= 32'b00000000010000010000000100010011;
ROM[7557] <= 32'b00000000010000010010000000100011;
ROM[7558] <= 32'b00000000010000010000000100010011;
ROM[7559] <= 32'b00000000010100010010000000100011;
ROM[7560] <= 32'b00000000010000010000000100010011;
ROM[7561] <= 32'b00000000011000010010000000100011;
ROM[7562] <= 32'b00000000010000010000000100010011;
ROM[7563] <= 32'b00000001010000000000001110010011;
ROM[7564] <= 32'b00000000100000111000001110010011;
ROM[7565] <= 32'b01000000011100010000001110110011;
ROM[7566] <= 32'b00000000011100000000001000110011;
ROM[7567] <= 32'b00000000001000000000000110110011;
ROM[7568] <= 32'b01100111110000001010000011101111;
ROM[7569] <= 32'b11111111110000010000000100010011;
ROM[7570] <= 32'b00000000000000010010001110000011;
ROM[7571] <= 32'b00000000011101100010000000100011;
ROM[7572] <= 32'b00000010000000011010001110000011;
ROM[7573] <= 32'b00000000011100010010000000100011;
ROM[7574] <= 32'b00000000010000010000000100010011;
ROM[7575] <= 32'b00000010000000000000001110010011;
ROM[7576] <= 32'b00000000011100010010000000100011;
ROM[7577] <= 32'b00000000010000010000000100010011;
ROM[7578] <= 32'b00000000000000000111001110110111;
ROM[7579] <= 32'b01101011010000111000001110010011;
ROM[7580] <= 32'b00000000111000111000001110110011;
ROM[7581] <= 32'b00000000011100010010000000100011;
ROM[7582] <= 32'b00000000010000010000000100010011;
ROM[7583] <= 32'b00000000001100010010000000100011;
ROM[7584] <= 32'b00000000010000010000000100010011;
ROM[7585] <= 32'b00000000010000010010000000100011;
ROM[7586] <= 32'b00000000010000010000000100010011;
ROM[7587] <= 32'b00000000010100010010000000100011;
ROM[7588] <= 32'b00000000010000010000000100010011;
ROM[7589] <= 32'b00000000011000010010000000100011;
ROM[7590] <= 32'b00000000010000010000000100010011;
ROM[7591] <= 32'b00000001010000000000001110010011;
ROM[7592] <= 32'b00000000100000111000001110010011;
ROM[7593] <= 32'b01000000011100010000001110110011;
ROM[7594] <= 32'b00000000011100000000001000110011;
ROM[7595] <= 32'b00000000001000000000000110110011;
ROM[7596] <= 32'b01100000110000001010000011101111;
ROM[7597] <= 32'b11111111110000010000000100010011;
ROM[7598] <= 32'b00000000000000010010001110000011;
ROM[7599] <= 32'b00000000011101100010000000100011;
ROM[7600] <= 32'b00000010000000011010001110000011;
ROM[7601] <= 32'b00000010011100011010000000100011;
ROM[7602] <= 32'b00000001010000011010001110000011;
ROM[7603] <= 32'b00000000011100010010000000100011;
ROM[7604] <= 32'b00000000010000010000000100010011;
ROM[7605] <= 32'b00000000000000000111001110110111;
ROM[7606] <= 32'b01110010000000111000001110010011;
ROM[7607] <= 32'b00000000111000111000001110110011;
ROM[7608] <= 32'b00000000011100010010000000100011;
ROM[7609] <= 32'b00000000010000010000000100010011;
ROM[7610] <= 32'b00000000001100010010000000100011;
ROM[7611] <= 32'b00000000010000010000000100010011;
ROM[7612] <= 32'b00000000010000010010000000100011;
ROM[7613] <= 32'b00000000010000010000000100010011;
ROM[7614] <= 32'b00000000010100010010000000100011;
ROM[7615] <= 32'b00000000010000010000000100010011;
ROM[7616] <= 32'b00000000011000010010000000100011;
ROM[7617] <= 32'b00000000010000010000000100010011;
ROM[7618] <= 32'b00000001010000000000001110010011;
ROM[7619] <= 32'b00000000010000111000001110010011;
ROM[7620] <= 32'b01000000011100010000001110110011;
ROM[7621] <= 32'b00000000011100000000001000110011;
ROM[7622] <= 32'b00000000001000000000000110110011;
ROM[7623] <= 32'b01111001100100001000000011101111;
ROM[7624] <= 32'b11111111110000010000000100010011;
ROM[7625] <= 32'b00000000000000010010001110000011;
ROM[7626] <= 32'b00000000011101100010000000100011;
ROM[7627] <= 32'b00000000000000011010001110000011;
ROM[7628] <= 32'b00000000011100010010000000100011;
ROM[7629] <= 32'b00000000010000010000000100010011;
ROM[7630] <= 32'b00000000010000011010001110000011;
ROM[7631] <= 32'b11111111110000010000000100010011;
ROM[7632] <= 32'b00000000000000010010010000000011;
ROM[7633] <= 32'b00000000011101000010001110110011;
ROM[7634] <= 32'b01000000011100000000001110110011;
ROM[7635] <= 32'b00000000000100111000001110010011;
ROM[7636] <= 32'b00000000000000111000101001100011;
ROM[7637] <= 32'b00000000000000001000001110110111;
ROM[7638] <= 32'b00010011100000111000001110010011;
ROM[7639] <= 32'b00000000111000111000001110110011;
ROM[7640] <= 32'b00000000000000111000000011100111;
ROM[7641] <= 32'b00000000100000011010001110000011;
ROM[7642] <= 32'b00000000011100010010000000100011;
ROM[7643] <= 32'b00000000010000010000000100010011;
ROM[7644] <= 32'b00000000000000000111001110110111;
ROM[7645] <= 32'b01111011110000111000001110010011;
ROM[7646] <= 32'b00000000111000111000001110110011;
ROM[7647] <= 32'b00000000011100010010000000100011;
ROM[7648] <= 32'b00000000010000010000000100010011;
ROM[7649] <= 32'b00000000001100010010000000100011;
ROM[7650] <= 32'b00000000010000010000000100010011;
ROM[7651] <= 32'b00000000010000010010000000100011;
ROM[7652] <= 32'b00000000010000010000000100010011;
ROM[7653] <= 32'b00000000010100010010000000100011;
ROM[7654] <= 32'b00000000010000010000000100010011;
ROM[7655] <= 32'b00000000011000010010000000100011;
ROM[7656] <= 32'b00000000010000010000000100010011;
ROM[7657] <= 32'b00000001010000000000001110010011;
ROM[7658] <= 32'b00000000010000111000001110010011;
ROM[7659] <= 32'b01000000011100010000001110110011;
ROM[7660] <= 32'b00000000011100000000001000110011;
ROM[7661] <= 32'b00000000001000000000000110110011;
ROM[7662] <= 32'b10000000010011111110000011101111;
ROM[7663] <= 32'b11111111110000010000000100010011;
ROM[7664] <= 32'b00000000000000010010001110000011;
ROM[7665] <= 32'b00000010011100011010001000100011;
ROM[7666] <= 32'b00000010010000011010001110000011;
ROM[7667] <= 32'b00000000011100010010000000100011;
ROM[7668] <= 32'b00000000010000010000000100010011;
ROM[7669] <= 32'b00000000000000000000001110010011;
ROM[7670] <= 32'b00000000011100010010000000100011;
ROM[7671] <= 32'b00000000010000010000000100010011;
ROM[7672] <= 32'b00000000000000001000001110110111;
ROM[7673] <= 32'b10000010110000111000001110010011;
ROM[7674] <= 32'b00000000111000111000001110110011;
ROM[7675] <= 32'b00000000011100010010000000100011;
ROM[7676] <= 32'b00000000010000010000000100010011;
ROM[7677] <= 32'b00000000001100010010000000100011;
ROM[7678] <= 32'b00000000010000010000000100010011;
ROM[7679] <= 32'b00000000010000010010000000100011;
ROM[7680] <= 32'b00000000010000010000000100010011;
ROM[7681] <= 32'b00000000010100010010000000100011;
ROM[7682] <= 32'b00000000010000010000000100010011;
ROM[7683] <= 32'b00000000011000010010000000100011;
ROM[7684] <= 32'b00000000010000010000000100010011;
ROM[7685] <= 32'b00000001010000000000001110010011;
ROM[7686] <= 32'b00000000100000111000001110010011;
ROM[7687] <= 32'b01000000011100010000001110110011;
ROM[7688] <= 32'b00000000011100000000001000110011;
ROM[7689] <= 32'b00000000001000000000000110110011;
ROM[7690] <= 32'b00101001110000001010000011101111;
ROM[7691] <= 32'b11111111110000010000000100010011;
ROM[7692] <= 32'b00000000000000010010001110000011;
ROM[7693] <= 32'b00000100011100011010000000100011;
ROM[7694] <= 32'b00000100000000011010001110000011;
ROM[7695] <= 32'b00000000011100010010000000100011;
ROM[7696] <= 32'b00000000010000010000000100010011;
ROM[7697] <= 32'b00000100010000011010001110000011;
ROM[7698] <= 32'b11111111110000010000000100010011;
ROM[7699] <= 32'b00000000000000010010010000000011;
ROM[7700] <= 32'b00000000011101000010010010110011;
ROM[7701] <= 32'b00000000100000111010010100110011;
ROM[7702] <= 32'b00000000101001001000001110110011;
ROM[7703] <= 32'b00000000000100111000001110010011;
ROM[7704] <= 32'b00000000000100111111001110010011;
ROM[7705] <= 32'b00000000000000111000101001100011;
ROM[7706] <= 32'b00000000000000001000001110110111;
ROM[7707] <= 32'b10000111110000111000001110010011;
ROM[7708] <= 32'b00000000111000111000001110110011;
ROM[7709] <= 32'b00000000000000111000000011100111;
ROM[7710] <= 32'b00011111000000000000000011101111;
ROM[7711] <= 32'b00000000000000001000001110110111;
ROM[7712] <= 32'b10001100100000111000001110010011;
ROM[7713] <= 32'b00000000111000111000001110110011;
ROM[7714] <= 32'b00000000011100010010000000100011;
ROM[7715] <= 32'b00000000010000010000000100010011;
ROM[7716] <= 32'b00000000001100010010000000100011;
ROM[7717] <= 32'b00000000010000010000000100010011;
ROM[7718] <= 32'b00000000010000010010000000100011;
ROM[7719] <= 32'b00000000010000010000000100010011;
ROM[7720] <= 32'b00000000010100010010000000100011;
ROM[7721] <= 32'b00000000010000010000000100010011;
ROM[7722] <= 32'b00000000011000010010000000100011;
ROM[7723] <= 32'b00000000010000010000000100010011;
ROM[7724] <= 32'b00000001010000000000001110010011;
ROM[7725] <= 32'b00000000000000111000001110010011;
ROM[7726] <= 32'b01000000011100010000001110110011;
ROM[7727] <= 32'b00000000011100000000001000110011;
ROM[7728] <= 32'b00000000001000000000000110110011;
ROM[7729] <= 32'b00011010000000001001000011101111;
ROM[7730] <= 32'b11111111110000010000000100010011;
ROM[7731] <= 32'b00000000000000010010001110000011;
ROM[7732] <= 32'b00000000011101100010000000100011;
ROM[7733] <= 32'b00000001010000011010001110000011;
ROM[7734] <= 32'b00000000011100010010000000100011;
ROM[7735] <= 32'b00000000010000010000000100010011;
ROM[7736] <= 32'b00000000000000001000001110110111;
ROM[7737] <= 32'b10010010110000111000001110010011;
ROM[7738] <= 32'b00000000111000111000001110110011;
ROM[7739] <= 32'b00000000011100010010000000100011;
ROM[7740] <= 32'b00000000010000010000000100010011;
ROM[7741] <= 32'b00000000001100010010000000100011;
ROM[7742] <= 32'b00000000010000010000000100010011;
ROM[7743] <= 32'b00000000010000010010000000100011;
ROM[7744] <= 32'b00000000010000010000000100010011;
ROM[7745] <= 32'b00000000010100010010000000100011;
ROM[7746] <= 32'b00000000010000010000000100010011;
ROM[7747] <= 32'b00000000011000010010000000100011;
ROM[7748] <= 32'b00000000010000010000000100010011;
ROM[7749] <= 32'b00000001010000000000001110010011;
ROM[7750] <= 32'b00000000010000111000001110010011;
ROM[7751] <= 32'b01000000011100010000001110110011;
ROM[7752] <= 32'b00000000011100000000001000110011;
ROM[7753] <= 32'b00000000001000000000000110110011;
ROM[7754] <= 32'b01011000110100001000000011101111;
ROM[7755] <= 32'b11111111110000010000000100010011;
ROM[7756] <= 32'b00000000000000010010001110000011;
ROM[7757] <= 32'b00000000011101100010000000100011;
ROM[7758] <= 32'b00000001100000011010001110000011;
ROM[7759] <= 32'b00000000011100010010000000100011;
ROM[7760] <= 32'b00000000010000010000000100010011;
ROM[7761] <= 32'b00000000000000001000001110110111;
ROM[7762] <= 32'b10011001000000111000001110010011;
ROM[7763] <= 32'b00000000111000111000001110110011;
ROM[7764] <= 32'b00000000011100010010000000100011;
ROM[7765] <= 32'b00000000010000010000000100010011;
ROM[7766] <= 32'b00000000001100010010000000100011;
ROM[7767] <= 32'b00000000010000010000000100010011;
ROM[7768] <= 32'b00000000010000010010000000100011;
ROM[7769] <= 32'b00000000010000010000000100010011;
ROM[7770] <= 32'b00000000010100010010000000100011;
ROM[7771] <= 32'b00000000010000010000000100010011;
ROM[7772] <= 32'b00000000011000010010000000100011;
ROM[7773] <= 32'b00000000010000010000000100010011;
ROM[7774] <= 32'b00000001010000000000001110010011;
ROM[7775] <= 32'b00000000010000111000001110010011;
ROM[7776] <= 32'b01000000011100010000001110110011;
ROM[7777] <= 32'b00000000011100000000001000110011;
ROM[7778] <= 32'b00000000001000000000000110110011;
ROM[7779] <= 32'b01010010100100001000000011101111;
ROM[7780] <= 32'b11111111110000010000000100010011;
ROM[7781] <= 32'b00000000000000010010001110000011;
ROM[7782] <= 32'b00000000011101100010000000100011;
ROM[7783] <= 32'b00000001110000011010001110000011;
ROM[7784] <= 32'b00000000011100010010000000100011;
ROM[7785] <= 32'b00000000010000010000000100010011;
ROM[7786] <= 32'b00000000000000001000001110110111;
ROM[7787] <= 32'b10011111010000111000001110010011;
ROM[7788] <= 32'b00000000111000111000001110110011;
ROM[7789] <= 32'b00000000011100010010000000100011;
ROM[7790] <= 32'b00000000010000010000000100010011;
ROM[7791] <= 32'b00000000001100010010000000100011;
ROM[7792] <= 32'b00000000010000010000000100010011;
ROM[7793] <= 32'b00000000010000010010000000100011;
ROM[7794] <= 32'b00000000010000010000000100010011;
ROM[7795] <= 32'b00000000010100010010000000100011;
ROM[7796] <= 32'b00000000010000010000000100010011;
ROM[7797] <= 32'b00000000011000010010000000100011;
ROM[7798] <= 32'b00000000010000010000000100010011;
ROM[7799] <= 32'b00000001010000000000001110010011;
ROM[7800] <= 32'b00000000010000111000001110010011;
ROM[7801] <= 32'b01000000011100010000001110110011;
ROM[7802] <= 32'b00000000011100000000001000110011;
ROM[7803] <= 32'b00000000001000000000000110110011;
ROM[7804] <= 32'b01001100010100001000000011101111;
ROM[7805] <= 32'b11111111110000010000000100010011;
ROM[7806] <= 32'b00000000000000010010001110000011;
ROM[7807] <= 32'b00000000011101100010000000100011;
ROM[7808] <= 32'b00000010000000011010001110000011;
ROM[7809] <= 32'b00000000011100010010000000100011;
ROM[7810] <= 32'b00000000010000010000000100010011;
ROM[7811] <= 32'b00000000000000001000001110110111;
ROM[7812] <= 32'b10100101100000111000001110010011;
ROM[7813] <= 32'b00000000111000111000001110110011;
ROM[7814] <= 32'b00000000011100010010000000100011;
ROM[7815] <= 32'b00000000010000010000000100010011;
ROM[7816] <= 32'b00000000001100010010000000100011;
ROM[7817] <= 32'b00000000010000010000000100010011;
ROM[7818] <= 32'b00000000010000010010000000100011;
ROM[7819] <= 32'b00000000010000010000000100010011;
ROM[7820] <= 32'b00000000010100010010000000100011;
ROM[7821] <= 32'b00000000010000010000000100010011;
ROM[7822] <= 32'b00000000011000010010000000100011;
ROM[7823] <= 32'b00000000010000010000000100010011;
ROM[7824] <= 32'b00000001010000000000001110010011;
ROM[7825] <= 32'b00000000010000111000001110010011;
ROM[7826] <= 32'b01000000011100010000001110110011;
ROM[7827] <= 32'b00000000011100000000001000110011;
ROM[7828] <= 32'b00000000001000000000000110110011;
ROM[7829] <= 32'b01000110000100001000000011101111;
ROM[7830] <= 32'b11111111110000010000000100010011;
ROM[7831] <= 32'b00000000000000010010001110000011;
ROM[7832] <= 32'b00000000011101100010000000100011;
ROM[7833] <= 32'b01100111100000000000000011101111;
ROM[7834] <= 32'b00000100000000011010001110000011;
ROM[7835] <= 32'b00000000011100010010000000100011;
ROM[7836] <= 32'b00000000010000010000000100010011;
ROM[7837] <= 32'b00000100100000011010001110000011;
ROM[7838] <= 32'b11111111110000010000000100010011;
ROM[7839] <= 32'b00000000000000010010010000000011;
ROM[7840] <= 32'b00000000011101000010010010110011;
ROM[7841] <= 32'b00000000100000111010010100110011;
ROM[7842] <= 32'b00000000101001001000001110110011;
ROM[7843] <= 32'b00000000000100111000001110010011;
ROM[7844] <= 32'b00000000000100111111001110010011;
ROM[7845] <= 32'b00000000000000111000101001100011;
ROM[7846] <= 32'b00000000000000001000001110110111;
ROM[7847] <= 32'b10101010110000111000001110010011;
ROM[7848] <= 32'b00000000111000111000001110110011;
ROM[7849] <= 32'b00000000000000111000000011100111;
ROM[7850] <= 32'b00001101000000000000000011101111;
ROM[7851] <= 32'b00000000000000001000001110110111;
ROM[7852] <= 32'b10101111100000111000001110010011;
ROM[7853] <= 32'b00000000111000111000001110110011;
ROM[7854] <= 32'b00000000011100010010000000100011;
ROM[7855] <= 32'b00000000010000010000000100010011;
ROM[7856] <= 32'b00000000001100010010000000100011;
ROM[7857] <= 32'b00000000010000010000000100010011;
ROM[7858] <= 32'b00000000010000010010000000100011;
ROM[7859] <= 32'b00000000010000010000000100010011;
ROM[7860] <= 32'b00000000010100010010000000100011;
ROM[7861] <= 32'b00000000010000010000000100010011;
ROM[7862] <= 32'b00000000011000010010000000100011;
ROM[7863] <= 32'b00000000010000010000000100010011;
ROM[7864] <= 32'b00000001010000000000001110010011;
ROM[7865] <= 32'b00000000000000111000001110010011;
ROM[7866] <= 32'b01000000011100010000001110110011;
ROM[7867] <= 32'b00000000011100000000001000110011;
ROM[7868] <= 32'b00000000001000000000000110110011;
ROM[7869] <= 32'b01001011110100001001000011101111;
ROM[7870] <= 32'b11111111110000010000000100010011;
ROM[7871] <= 32'b00000000000000010010001110000011;
ROM[7872] <= 32'b00000000011101100010000000100011;
ROM[7873] <= 32'b00000000000000000000001110010011;
ROM[7874] <= 32'b00000000011100010010000000100011;
ROM[7875] <= 32'b00000000010000010000000100010011;
ROM[7876] <= 32'b00000000000000000000001110010011;
ROM[7877] <= 32'b00000000011100010010000000100011;
ROM[7878] <= 32'b00000000010000010000000100010011;
ROM[7879] <= 32'b00000000000000001000001110110111;
ROM[7880] <= 32'b10110110100000111000001110010011;
ROM[7881] <= 32'b00000000111000111000001110110011;
ROM[7882] <= 32'b00000000011100010010000000100011;
ROM[7883] <= 32'b00000000010000010000000100010011;
ROM[7884] <= 32'b00000000001100010010000000100011;
ROM[7885] <= 32'b00000000010000010000000100010011;
ROM[7886] <= 32'b00000000010000010010000000100011;
ROM[7887] <= 32'b00000000010000010000000100010011;
ROM[7888] <= 32'b00000000010100010010000000100011;
ROM[7889] <= 32'b00000000010000010000000100010011;
ROM[7890] <= 32'b00000000011000010010000000100011;
ROM[7891] <= 32'b00000000010000010000000100010011;
ROM[7892] <= 32'b00000001010000000000001110010011;
ROM[7893] <= 32'b00000000100000111000001110010011;
ROM[7894] <= 32'b01000000011100010000001110110011;
ROM[7895] <= 32'b00000000011100000000001000110011;
ROM[7896] <= 32'b00000000001000000000000110110011;
ROM[7897] <= 32'b01011000100100000111000011101111;
ROM[7898] <= 32'b11111111110000010000000100010011;
ROM[7899] <= 32'b00000000000000010010001110000011;
ROM[7900] <= 32'b00000000011101100010000000100011;
ROM[7901] <= 32'b01010110100000000000000011101111;
ROM[7902] <= 32'b00000100000000011010001110000011;
ROM[7903] <= 32'b00000000011100010010000000100011;
ROM[7904] <= 32'b00000000010000010000000100010011;
ROM[7905] <= 32'b00000100110000011010001110000011;
ROM[7906] <= 32'b11111111110000010000000100010011;
ROM[7907] <= 32'b00000000000000010010010000000011;
ROM[7908] <= 32'b00000000011101000010010010110011;
ROM[7909] <= 32'b00000000100000111010010100110011;
ROM[7910] <= 32'b00000000101001001000001110110011;
ROM[7911] <= 32'b00000000000100111000001110010011;
ROM[7912] <= 32'b00000000000100111111001110010011;
ROM[7913] <= 32'b00000000000000111000101001100011;
ROM[7914] <= 32'b00000000000000001000001110110111;
ROM[7915] <= 32'b10111011110000111000001110010011;
ROM[7916] <= 32'b00000000111000111000001110110011;
ROM[7917] <= 32'b00000000000000111000000011100111;
ROM[7918] <= 32'b00000001000000000000000011101111;
ROM[7919] <= 32'b00000000001000000000001110010011;
ROM[7920] <= 32'b00000000011100011010000000100011;
ROM[7921] <= 32'b01010001100000000000000011101111;
ROM[7922] <= 32'b00000100000000011010001110000011;
ROM[7923] <= 32'b00000000011100010010000000100011;
ROM[7924] <= 32'b00000000010000010000000100010011;
ROM[7925] <= 32'b00000101000000011010001110000011;
ROM[7926] <= 32'b11111111110000010000000100010011;
ROM[7927] <= 32'b00000000000000010010010000000011;
ROM[7928] <= 32'b00000000011101000010010010110011;
ROM[7929] <= 32'b00000000100000111010010100110011;
ROM[7930] <= 32'b00000000101001001000001110110011;
ROM[7931] <= 32'b00000000000100111000001110010011;
ROM[7932] <= 32'b00000000000100111111001110010011;
ROM[7933] <= 32'b00000000000000111000101001100011;
ROM[7934] <= 32'b00000000000000001000001110110111;
ROM[7935] <= 32'b11000000110000111000001110010011;
ROM[7936] <= 32'b00000000111000111000001110110011;
ROM[7937] <= 32'b00000000000000111000000011100111;
ROM[7938] <= 32'b01000011010000000000000011101111;
ROM[7939] <= 32'b00000000001100000000001110010011;
ROM[7940] <= 32'b00000000011100010010000000100011;
ROM[7941] <= 32'b00000000010000010000000100010011;
ROM[7942] <= 32'b00000000000000001000001110110111;
ROM[7943] <= 32'b11000110010000111000001110010011;
ROM[7944] <= 32'b00000000111000111000001110110011;
ROM[7945] <= 32'b00000000011100010010000000100011;
ROM[7946] <= 32'b00000000010000010000000100010011;
ROM[7947] <= 32'b00000000001100010010000000100011;
ROM[7948] <= 32'b00000000010000010000000100010011;
ROM[7949] <= 32'b00000000010000010010000000100011;
ROM[7950] <= 32'b00000000010000010000000100010011;
ROM[7951] <= 32'b00000000010100010010000000100011;
ROM[7952] <= 32'b00000000010000010000000100010011;
ROM[7953] <= 32'b00000000011000010010000000100011;
ROM[7954] <= 32'b00000000010000010000000100010011;
ROM[7955] <= 32'b00000001010000000000001110010011;
ROM[7956] <= 32'b00000000010000111000001110010011;
ROM[7957] <= 32'b01000000011100010000001110110011;
ROM[7958] <= 32'b00000000011100000000001000110011;
ROM[7959] <= 32'b00000000001000000000000110110011;
ROM[7960] <= 32'b01001010000100001001000011101111;
ROM[7961] <= 32'b11111111110000010000000100010011;
ROM[7962] <= 32'b00000000000000010010001110000011;
ROM[7963] <= 32'b00000010011100011010111000100011;
ROM[7964] <= 32'b00000011110000011010001110000011;
ROM[7965] <= 32'b00000000011100010010000000100011;
ROM[7966] <= 32'b00000000010000010000000100010011;
ROM[7967] <= 32'b00000110111000000000001110010011;
ROM[7968] <= 32'b00000000011100010010000000100011;
ROM[7969] <= 32'b00000000010000010000000100010011;
ROM[7970] <= 32'b00000000000000001000001110110111;
ROM[7971] <= 32'b11001101010000111000001110010011;
ROM[7972] <= 32'b00000000111000111000001110110011;
ROM[7973] <= 32'b00000000011100010010000000100011;
ROM[7974] <= 32'b00000000010000010000000100010011;
ROM[7975] <= 32'b00000000001100010010000000100011;
ROM[7976] <= 32'b00000000010000010000000100010011;
ROM[7977] <= 32'b00000000010000010010000000100011;
ROM[7978] <= 32'b00000000010000010000000100010011;
ROM[7979] <= 32'b00000000010100010010000000100011;
ROM[7980] <= 32'b00000000010000010000000100010011;
ROM[7981] <= 32'b00000000011000010010000000100011;
ROM[7982] <= 32'b00000000010000010000000100010011;
ROM[7983] <= 32'b00000001010000000000001110010011;
ROM[7984] <= 32'b00000000100000111000001110010011;
ROM[7985] <= 32'b01000000011100010000001110110011;
ROM[7986] <= 32'b00000000011100000000001000110011;
ROM[7987] <= 32'b00000000001000000000000110110011;
ROM[7988] <= 32'b01111110110100001001000011101111;
ROM[7989] <= 32'b11111111110000010000000100010011;
ROM[7990] <= 32'b00000000000000010010001110000011;
ROM[7991] <= 32'b00000000011101100010000000100011;
ROM[7992] <= 32'b00000011110000011010001110000011;
ROM[7993] <= 32'b00000000011100010010000000100011;
ROM[7994] <= 32'b00000000010000010000000100010011;
ROM[7995] <= 32'b00000011101000000000001110010011;
ROM[7996] <= 32'b00000000011100010010000000100011;
ROM[7997] <= 32'b00000000010000010000000100010011;
ROM[7998] <= 32'b00000000000000001000001110110111;
ROM[7999] <= 32'b11010100010000111000001110010011;
ROM[8000] <= 32'b00000000111000111000001110110011;
ROM[8001] <= 32'b00000000011100010010000000100011;
ROM[8002] <= 32'b00000000010000010000000100010011;
ROM[8003] <= 32'b00000000001100010010000000100011;
ROM[8004] <= 32'b00000000010000010000000100010011;
ROM[8005] <= 32'b00000000010000010010000000100011;
ROM[8006] <= 32'b00000000010000010000000100010011;
ROM[8007] <= 32'b00000000010100010010000000100011;
ROM[8008] <= 32'b00000000010000010000000100010011;
ROM[8009] <= 32'b00000000011000010010000000100011;
ROM[8010] <= 32'b00000000010000010000000100010011;
ROM[8011] <= 32'b00000001010000000000001110010011;
ROM[8012] <= 32'b00000000100000111000001110010011;
ROM[8013] <= 32'b01000000011100010000001110110011;
ROM[8014] <= 32'b00000000011100000000001000110011;
ROM[8015] <= 32'b00000000001000000000000110110011;
ROM[8016] <= 32'b01110111110100001001000011101111;
ROM[8017] <= 32'b11111111110000010000000100010011;
ROM[8018] <= 32'b00000000000000010010001110000011;
ROM[8019] <= 32'b00000000011101100010000000100011;
ROM[8020] <= 32'b00000011110000011010001110000011;
ROM[8021] <= 32'b00000000011100010010000000100011;
ROM[8022] <= 32'b00000000010000010000000100010011;
ROM[8023] <= 32'b00000010000000000000001110010011;
ROM[8024] <= 32'b00000000011100010010000000100011;
ROM[8025] <= 32'b00000000010000010000000100010011;
ROM[8026] <= 32'b00000000000000001000001110110111;
ROM[8027] <= 32'b11011011010000111000001110010011;
ROM[8028] <= 32'b00000000111000111000001110110011;
ROM[8029] <= 32'b00000000011100010010000000100011;
ROM[8030] <= 32'b00000000010000010000000100010011;
ROM[8031] <= 32'b00000000001100010010000000100011;
ROM[8032] <= 32'b00000000010000010000000100010011;
ROM[8033] <= 32'b00000000010000010010000000100011;
ROM[8034] <= 32'b00000000010000010000000100010011;
ROM[8035] <= 32'b00000000010100010010000000100011;
ROM[8036] <= 32'b00000000010000010000000100010011;
ROM[8037] <= 32'b00000000011000010010000000100011;
ROM[8038] <= 32'b00000000010000010000000100010011;
ROM[8039] <= 32'b00000001010000000000001110010011;
ROM[8040] <= 32'b00000000100000111000001110010011;
ROM[8041] <= 32'b01000000011100010000001110110011;
ROM[8042] <= 32'b00000000011100000000001000110011;
ROM[8043] <= 32'b00000000001000000000000110110011;
ROM[8044] <= 32'b01110000110100001001000011101111;
ROM[8045] <= 32'b11111111110000010000000100010011;
ROM[8046] <= 32'b00000000000000010010001110000011;
ROM[8047] <= 32'b00000000011101100010000000100011;
ROM[8048] <= 32'b00000011110000011010001110000011;
ROM[8049] <= 32'b00000010011100011010111000100011;
ROM[8050] <= 32'b00000011110000011010001110000011;
ROM[8051] <= 32'b00000000011100010010000000100011;
ROM[8052] <= 32'b00000000010000010000000100010011;
ROM[8053] <= 32'b00000000000000001000001110110111;
ROM[8054] <= 32'b11100010000000111000001110010011;
ROM[8055] <= 32'b00000000111000111000001110110011;
ROM[8056] <= 32'b00000000011100010010000000100011;
ROM[8057] <= 32'b00000000010000010000000100010011;
ROM[8058] <= 32'b00000000001100010010000000100011;
ROM[8059] <= 32'b00000000010000010000000100010011;
ROM[8060] <= 32'b00000000010000010010000000100011;
ROM[8061] <= 32'b00000000010000010000000100010011;
ROM[8062] <= 32'b00000000010100010010000000100011;
ROM[8063] <= 32'b00000000010000010000000100010011;
ROM[8064] <= 32'b00000000011000010010000000100011;
ROM[8065] <= 32'b00000000010000010000000100010011;
ROM[8066] <= 32'b00000001010000000000001110010011;
ROM[8067] <= 32'b00000000010000111000001110010011;
ROM[8068] <= 32'b01000000011100010000001110110011;
ROM[8069] <= 32'b00000000011100000000001000110011;
ROM[8070] <= 32'b00000000001000000000000110110011;
ROM[8071] <= 32'b11011101010111111101000011101111;
ROM[8072] <= 32'b11111111110000010000000100010011;
ROM[8073] <= 32'b00000000000000010010001110000011;
ROM[8074] <= 32'b00000010011100011010010000100011;
ROM[8075] <= 32'b00000000000000000000001110010011;
ROM[8076] <= 32'b00000010011100011010011000100011;
ROM[8077] <= 32'b00000000000100000000001110010011;
ROM[8078] <= 32'b00000010011100011010100000100011;
ROM[8079] <= 32'b00000010100000011010001110000011;
ROM[8080] <= 32'b00000000011100010010000000100011;
ROM[8081] <= 32'b00000000010000010000000100010011;
ROM[8082] <= 32'b00000000000100000000001110010011;
ROM[8083] <= 32'b11111111110000010000000100010011;
ROM[8084] <= 32'b00000000000000010010010000000011;
ROM[8085] <= 32'b00000000011101000010010010110011;
ROM[8086] <= 32'b00000000100000111010010100110011;
ROM[8087] <= 32'b00000000101001001000001110110011;
ROM[8088] <= 32'b00000000000100111000001110010011;
ROM[8089] <= 32'b00000000000100111111001110010011;
ROM[8090] <= 32'b00000000000000111000101001100011;
ROM[8091] <= 32'b00000000000000001000001110110111;
ROM[8092] <= 32'b11101000000000111000001110010011;
ROM[8093] <= 32'b00000000111000111000001110110011;
ROM[8094] <= 32'b00000000000000111000000011100111;
ROM[8095] <= 32'b00000110110000000000000011101111;
ROM[8096] <= 32'b00000011000000011010001110000011;
ROM[8097] <= 32'b00000000011100010010000000100011;
ROM[8098] <= 32'b00000000010000010000000100010011;
ROM[8099] <= 32'b00000000000000001000001110110111;
ROM[8100] <= 32'b11101101100000111000001110010011;
ROM[8101] <= 32'b00000000111000111000001110110011;
ROM[8102] <= 32'b00000000011100010010000000100011;
ROM[8103] <= 32'b00000000010000010000000100010011;
ROM[8104] <= 32'b00000000001100010010000000100011;
ROM[8105] <= 32'b00000000010000010000000100010011;
ROM[8106] <= 32'b00000000010000010010000000100011;
ROM[8107] <= 32'b00000000010000010000000100010011;
ROM[8108] <= 32'b00000000010100010010000000100011;
ROM[8109] <= 32'b00000000010000010000000100010011;
ROM[8110] <= 32'b00000000011000010010000000100011;
ROM[8111] <= 32'b00000000010000010000000100010011;
ROM[8112] <= 32'b00000001010000000000001110010011;
ROM[8113] <= 32'b00000000010000111000001110010011;
ROM[8114] <= 32'b01000000011100010000001110110011;
ROM[8115] <= 32'b00000000011100000000001000110011;
ROM[8116] <= 32'b00000000001000000000000110110011;
ROM[8117] <= 32'b00011010100100001000000011101111;
ROM[8118] <= 32'b11111111110000010000000100010011;
ROM[8119] <= 32'b00000000000000010010001110000011;
ROM[8120] <= 32'b00000000011101100010000000100011;
ROM[8121] <= 32'b00000000010000000000000011101111;
ROM[8122] <= 32'b00000000001000000000001110010011;
ROM[8123] <= 32'b00000010011100011010110000100011;
ROM[8124] <= 32'b00000011100000011010001110000011;
ROM[8125] <= 32'b00000000011100010010000000100011;
ROM[8126] <= 32'b00000000010000010000000100010011;
ROM[8127] <= 32'b00000010100000011010001110000011;
ROM[8128] <= 32'b11111111110000010000000100010011;
ROM[8129] <= 32'b00000000000000010010010000000011;
ROM[8130] <= 32'b00000000011101000010001110110011;
ROM[8131] <= 32'b01000000011100000000001110110011;
ROM[8132] <= 32'b00000000000100111000001110010011;
ROM[8133] <= 32'b00000000000000111000101001100011;
ROM[8134] <= 32'b00000000000000001000001110110111;
ROM[8135] <= 32'b11110111110000111000001110010011;
ROM[8136] <= 32'b00000000111000111000001110110011;
ROM[8137] <= 32'b00000000000000111000000011100111;
ROM[8138] <= 32'b00000010110000011010001110000011;
ROM[8139] <= 32'b00000000011100010010000000100011;
ROM[8140] <= 32'b00000000010000010000000100010011;
ROM[8141] <= 32'b00000011000000011010001110000011;
ROM[8142] <= 32'b11111111110000010000000100010011;
ROM[8143] <= 32'b00000000000000010010010000000011;
ROM[8144] <= 32'b00000000011101000000001110110011;
ROM[8145] <= 32'b00000010011100011010101000100011;
ROM[8146] <= 32'b00000011000000011010001110000011;
ROM[8147] <= 32'b00000010011100011010011000100011;
ROM[8148] <= 32'b00000011010000011010001110000011;
ROM[8149] <= 32'b00000010011100011010100000100011;
ROM[8150] <= 32'b00000011100000011010001110000011;
ROM[8151] <= 32'b00000000011100010010000000100011;
ROM[8152] <= 32'b00000000010000010000000100010011;
ROM[8153] <= 32'b00000000000100000000001110010011;
ROM[8154] <= 32'b11111111110000010000000100010011;
ROM[8155] <= 32'b00000000000000010010010000000011;
ROM[8156] <= 32'b00000000011101000000001110110011;
ROM[8157] <= 32'b00000010011100011010110000100011;
ROM[8158] <= 32'b11110111100111111111000011101111;
ROM[8159] <= 32'b00000000000000001000001110110111;
ROM[8160] <= 32'b11111100100000111000001110010011;
ROM[8161] <= 32'b00000000111000111000001110110011;
ROM[8162] <= 32'b00000000011100010010000000100011;
ROM[8163] <= 32'b00000000010000010000000100010011;
ROM[8164] <= 32'b00000000001100010010000000100011;
ROM[8165] <= 32'b00000000010000010000000100010011;
ROM[8166] <= 32'b00000000010000010010000000100011;
ROM[8167] <= 32'b00000000010000010000000100010011;
ROM[8168] <= 32'b00000000010100010010000000100011;
ROM[8169] <= 32'b00000000010000010000000100010011;
ROM[8170] <= 32'b00000000011000010010000000100011;
ROM[8171] <= 32'b00000000010000010000000100010011;
ROM[8172] <= 32'b00000001010000000000001110010011;
ROM[8173] <= 32'b00000000000000111000001110010011;
ROM[8174] <= 32'b01000000011100010000001110110011;
ROM[8175] <= 32'b00000000011100000000001000110011;
ROM[8176] <= 32'b00000000001000000000000110110011;
ROM[8177] <= 32'b00101010000100001000000011101111;
ROM[8178] <= 32'b11111111110000010000000100010011;
ROM[8179] <= 32'b00000000000000010010001110000011;
ROM[8180] <= 32'b00000000011101100010000000100011;
ROM[8181] <= 32'b00000011010000011010001110000011;
ROM[8182] <= 32'b00000000011100010010000000100011;
ROM[8183] <= 32'b00000000010000010000000100010011;
ROM[8184] <= 32'b00000000000000001000001110110111;
ROM[8185] <= 32'b00000010110000111000001110010011;
ROM[8186] <= 32'b00000000111000111000001110110011;
ROM[8187] <= 32'b00000000011100010010000000100011;
ROM[8188] <= 32'b00000000010000010000000100010011;
ROM[8189] <= 32'b00000000001100010010000000100011;
ROM[8190] <= 32'b00000000010000010000000100010011;
ROM[8191] <= 32'b00000000010000010010000000100011;
ROM[8192] <= 32'b00000000010000010000000100010011;
ROM[8193] <= 32'b00000000010100010010000000100011;
ROM[8194] <= 32'b00000000010000010000000100010011;
ROM[8195] <= 32'b00000000011000010010000000100011;
ROM[8196] <= 32'b00000000010000010000000100010011;
ROM[8197] <= 32'b00000001010000000000001110010011;
ROM[8198] <= 32'b00000000010000111000001110010011;
ROM[8199] <= 32'b01000000011100010000001110110011;
ROM[8200] <= 32'b00000000011100000000001000110011;
ROM[8201] <= 32'b00000000001000000000000110110011;
ROM[8202] <= 32'b00000101010100001000000011101111;
ROM[8203] <= 32'b11111111110000010000000100010011;
ROM[8204] <= 32'b00000000000000010010001110000011;
ROM[8205] <= 32'b00000000011101100010000000100011;
ROM[8206] <= 32'b00001010010000000000000011101111;
ROM[8207] <= 32'b00000100000000011010001110000011;
ROM[8208] <= 32'b00000000011100010010000000100011;
ROM[8209] <= 32'b00000000010000010000000100010011;
ROM[8210] <= 32'b00000101110000011010001110000011;
ROM[8211] <= 32'b11111111110000010000000100010011;
ROM[8212] <= 32'b00000000000000010010010000000011;
ROM[8213] <= 32'b00000000011101000010010010110011;
ROM[8214] <= 32'b00000000100000111010010100110011;
ROM[8215] <= 32'b00000000101001001000001110110011;
ROM[8216] <= 32'b00000000000100111000001110010011;
ROM[8217] <= 32'b00000000000100111111001110010011;
ROM[8218] <= 32'b00000000000000111000101001100011;
ROM[8219] <= 32'b00000000000000001000001110110111;
ROM[8220] <= 32'b00001000000000111000001110010011;
ROM[8221] <= 32'b00000000111000111000001110110011;
ROM[8222] <= 32'b00000000000000111000000011100111;
ROM[8223] <= 32'b00000110000000000000000011101111;
ROM[8224] <= 32'b00000000000000001000001110110111;
ROM[8225] <= 32'b00001100110000111000001110010011;
ROM[8226] <= 32'b00000000111000111000001110110011;
ROM[8227] <= 32'b00000000011100010010000000100011;
ROM[8228] <= 32'b00000000010000010000000100010011;
ROM[8229] <= 32'b00000000001100010010000000100011;
ROM[8230] <= 32'b00000000010000010000000100010011;
ROM[8231] <= 32'b00000000010000010010000000100011;
ROM[8232] <= 32'b00000000010000010000000100010011;
ROM[8233] <= 32'b00000000010100010010000000100011;
ROM[8234] <= 32'b00000000010000010000000100010011;
ROM[8235] <= 32'b00000000011000010010000000100011;
ROM[8236] <= 32'b00000000010000010000000100010011;
ROM[8237] <= 32'b00000001010000000000001110010011;
ROM[8238] <= 32'b00000000000000111000001110010011;
ROM[8239] <= 32'b01000000011100010000001110110011;
ROM[8240] <= 32'b00000000011100000000001000110011;
ROM[8241] <= 32'b00000000001000000000000110110011;
ROM[8242] <= 32'b11001011010011111000000011101111;
ROM[8243] <= 32'b11111111110000010000000100010011;
ROM[8244] <= 32'b00000000000000010010001110000011;
ROM[8245] <= 32'b00000000011101100010000000100011;
ROM[8246] <= 32'b00000000010000000000000011101111;
ROM[8247] <= 32'b00000000000000001000001110110111;
ROM[8248] <= 32'b00010010100000111000001110010011;
ROM[8249] <= 32'b00000000111000111000001110110011;
ROM[8250] <= 32'b00000000011100010010000000100011;
ROM[8251] <= 32'b00000000010000010000000100010011;
ROM[8252] <= 32'b00000000001100010010000000100011;
ROM[8253] <= 32'b00000000010000010000000100010011;
ROM[8254] <= 32'b00000000010000010010000000100011;
ROM[8255] <= 32'b00000000010000010000000100010011;
ROM[8256] <= 32'b00000000010100010010000000100011;
ROM[8257] <= 32'b00000000010000010000000100010011;
ROM[8258] <= 32'b00000000011000010010000000100011;
ROM[8259] <= 32'b00000000010000010000000100010011;
ROM[8260] <= 32'b00000001010000000000001110010011;
ROM[8261] <= 32'b00000000000000111000001110010011;
ROM[8262] <= 32'b01000000011100010000001110110011;
ROM[8263] <= 32'b00000000011100000000001000110011;
ROM[8264] <= 32'b00000000001000000000000110110011;
ROM[8265] <= 32'b00010100000100001000000011101111;
ROM[8266] <= 32'b11111111110000010000000100010011;
ROM[8267] <= 32'b00000000000000010010001110000011;
ROM[8268] <= 32'b00000000011101100010000000100011;
ROM[8269] <= 32'b11011111100011111111000011101111;
ROM[8270] <= 32'b00000000000000000000001110010011;
ROM[8271] <= 32'b00000000011100010010000000100011;
ROM[8272] <= 32'b00000000010000010000000100010011;
ROM[8273] <= 32'b00000001010000000000001110010011;
ROM[8274] <= 32'b01000000011100011000001110110011;
ROM[8275] <= 32'b00000000000000111010000010000011;
ROM[8276] <= 32'b11111111110000010000000100010011;
ROM[8277] <= 32'b00000000000000010010001110000011;
ROM[8278] <= 32'b00000000011100100010000000100011;
ROM[8279] <= 32'b00000000010000100000000100010011;
ROM[8280] <= 32'b00000001010000000000001110010011;
ROM[8281] <= 32'b01000000011100011000001110110011;
ROM[8282] <= 32'b00000000010000111010000110000011;
ROM[8283] <= 32'b00000000100000111010001000000011;
ROM[8284] <= 32'b00000000110000111010001010000011;
ROM[8285] <= 32'b00000001000000111010001100000011;
ROM[8286] <= 32'b00000000000000001000000011100111;
ROM[8287] <= 32'b00000010000000000000001110010011;
ROM[8288] <= 32'b00000000011100010010000000100011;
ROM[8289] <= 32'b00000000010000010000000100010011;
ROM[8290] <= 32'b00000000000000001000001110110111;
ROM[8291] <= 32'b00011101010000111000001110010011;
ROM[8292] <= 32'b00000000111000111000001110110011;
ROM[8293] <= 32'b00000000011100010010000000100011;
ROM[8294] <= 32'b00000000010000010000000100010011;
ROM[8295] <= 32'b00000000001100010010000000100011;
ROM[8296] <= 32'b00000000010000010000000100010011;
ROM[8297] <= 32'b00000000010000010010000000100011;
ROM[8298] <= 32'b00000000010000010000000100010011;
ROM[8299] <= 32'b00000000010100010010000000100011;
ROM[8300] <= 32'b00000000010000010000000100010011;
ROM[8301] <= 32'b00000000011000010010000000100011;
ROM[8302] <= 32'b00000000010000010000000100010011;
ROM[8303] <= 32'b00000001010000000000001110010011;
ROM[8304] <= 32'b00000000010000111000001110010011;
ROM[8305] <= 32'b01000000011100010000001110110011;
ROM[8306] <= 32'b00000000011100000000001000110011;
ROM[8307] <= 32'b00000000001000000000000110110011;
ROM[8308] <= 32'b10100111000011111000000011101111;
ROM[8309] <= 32'b11111111110000010000000100010011;
ROM[8310] <= 32'b00000000000000010010001110000011;
ROM[8311] <= 32'b00000100011101101010010000100011;
ROM[8312] <= 32'b00000000000000000000001110010011;
ROM[8313] <= 32'b00000000011100010010000000100011;
ROM[8314] <= 32'b00000000010000010000000100010011;
ROM[8315] <= 32'b00000100100001101010001110000011;
ROM[8316] <= 32'b11111111110000010000000100010011;
ROM[8317] <= 32'b00000000000000010010010000000011;
ROM[8318] <= 32'b00000000011101000000001110110011;
ROM[8319] <= 32'b00000000011100010010000000100011;
ROM[8320] <= 32'b00000000010000010000000100010011;
ROM[8321] <= 32'b00000000000100000000001110010011;
ROM[8322] <= 32'b00000000011101100010000000100011;
ROM[8323] <= 32'b11111111110000010000000100010011;
ROM[8324] <= 32'b00000000000000010010001110000011;
ROM[8325] <= 32'b00000000000000111000001100010011;
ROM[8326] <= 32'b00000000000001100010001110000011;
ROM[8327] <= 32'b00000000110100110000010000110011;
ROM[8328] <= 32'b00000000011101000010000000100011;
ROM[8329] <= 32'b00000000010000000000001110010011;
ROM[8330] <= 32'b00000000011100010010000000100011;
ROM[8331] <= 32'b00000000010000010000000100010011;
ROM[8332] <= 32'b00000100100001101010001110000011;
ROM[8333] <= 32'b11111111110000010000000100010011;
ROM[8334] <= 32'b00000000000000010010010000000011;
ROM[8335] <= 32'b00000000011101000000001110110011;
ROM[8336] <= 32'b00000000011100010010000000100011;
ROM[8337] <= 32'b00000000010000010000000100010011;
ROM[8338] <= 32'b00000000001000000000001110010011;
ROM[8339] <= 32'b00000000011101100010000000100011;
ROM[8340] <= 32'b11111111110000010000000100010011;
ROM[8341] <= 32'b00000000000000010010001110000011;
ROM[8342] <= 32'b00000000000000111000001100010011;
ROM[8343] <= 32'b00000000000001100010001110000011;
ROM[8344] <= 32'b00000000110100110000010000110011;
ROM[8345] <= 32'b00000000011101000010000000100011;
ROM[8346] <= 32'b00000000100000000000001110010011;
ROM[8347] <= 32'b00000000011100010010000000100011;
ROM[8348] <= 32'b00000000010000010000000100010011;
ROM[8349] <= 32'b00000100100001101010001110000011;
ROM[8350] <= 32'b11111111110000010000000100010011;
ROM[8351] <= 32'b00000000000000010010010000000011;
ROM[8352] <= 32'b00000000011101000000001110110011;
ROM[8353] <= 32'b00000000011100010010000000100011;
ROM[8354] <= 32'b00000000010000010000000100010011;
ROM[8355] <= 32'b00000000010000000000001110010011;
ROM[8356] <= 32'b00000000011101100010000000100011;
ROM[8357] <= 32'b11111111110000010000000100010011;
ROM[8358] <= 32'b00000000000000010010001110000011;
ROM[8359] <= 32'b00000000000000111000001100010011;
ROM[8360] <= 32'b00000000000001100010001110000011;
ROM[8361] <= 32'b00000000110100110000010000110011;
ROM[8362] <= 32'b00000000011101000010000000100011;
ROM[8363] <= 32'b00000000110000000000001110010011;
ROM[8364] <= 32'b00000000011100010010000000100011;
ROM[8365] <= 32'b00000000010000010000000100010011;
ROM[8366] <= 32'b00000100100001101010001110000011;
ROM[8367] <= 32'b11111111110000010000000100010011;
ROM[8368] <= 32'b00000000000000010010010000000011;
ROM[8369] <= 32'b00000000011101000000001110110011;
ROM[8370] <= 32'b00000000011100010010000000100011;
ROM[8371] <= 32'b00000000010000010000000100010011;
ROM[8372] <= 32'b00000000100000000000001110010011;
ROM[8373] <= 32'b00000000011101100010000000100011;
ROM[8374] <= 32'b11111111110000010000000100010011;
ROM[8375] <= 32'b00000000000000010010001110000011;
ROM[8376] <= 32'b00000000000000111000001100010011;
ROM[8377] <= 32'b00000000000001100010001110000011;
ROM[8378] <= 32'b00000000110100110000010000110011;
ROM[8379] <= 32'b00000000011101000010000000100011;
ROM[8380] <= 32'b00000001000000000000001110010011;
ROM[8381] <= 32'b00000000011100010010000000100011;
ROM[8382] <= 32'b00000000010000010000000100010011;
ROM[8383] <= 32'b00000100100001101010001110000011;
ROM[8384] <= 32'b11111111110000010000000100010011;
ROM[8385] <= 32'b00000000000000010010010000000011;
ROM[8386] <= 32'b00000000011101000000001110110011;
ROM[8387] <= 32'b00000000011100010010000000100011;
ROM[8388] <= 32'b00000000010000010000000100010011;
ROM[8389] <= 32'b00000001000000000000001110010011;
ROM[8390] <= 32'b00000000011101100010000000100011;
ROM[8391] <= 32'b11111111110000010000000100010011;
ROM[8392] <= 32'b00000000000000010010001110000011;
ROM[8393] <= 32'b00000000000000111000001100010011;
ROM[8394] <= 32'b00000000000001100010001110000011;
ROM[8395] <= 32'b00000000110100110000010000110011;
ROM[8396] <= 32'b00000000011101000010000000100011;
ROM[8397] <= 32'b00000001010000000000001110010011;
ROM[8398] <= 32'b00000000011100010010000000100011;
ROM[8399] <= 32'b00000000010000010000000100010011;
ROM[8400] <= 32'b00000100100001101010001110000011;
ROM[8401] <= 32'b11111111110000010000000100010011;
ROM[8402] <= 32'b00000000000000010010010000000011;
ROM[8403] <= 32'b00000000011101000000001110110011;
ROM[8404] <= 32'b00000000011100010010000000100011;
ROM[8405] <= 32'b00000000010000010000000100010011;
ROM[8406] <= 32'b00000010000000000000001110010011;
ROM[8407] <= 32'b00000000011101100010000000100011;
ROM[8408] <= 32'b11111111110000010000000100010011;
ROM[8409] <= 32'b00000000000000010010001110000011;
ROM[8410] <= 32'b00000000000000111000001100010011;
ROM[8411] <= 32'b00000000000001100010001110000011;
ROM[8412] <= 32'b00000000110100110000010000110011;
ROM[8413] <= 32'b00000000011101000010000000100011;
ROM[8414] <= 32'b00000001100000000000001110010011;
ROM[8415] <= 32'b00000000011100010010000000100011;
ROM[8416] <= 32'b00000000010000010000000100010011;
ROM[8417] <= 32'b00000100100001101010001110000011;
ROM[8418] <= 32'b11111111110000010000000100010011;
ROM[8419] <= 32'b00000000000000010010010000000011;
ROM[8420] <= 32'b00000000011101000000001110110011;
ROM[8421] <= 32'b00000000011100010010000000100011;
ROM[8422] <= 32'b00000000010000010000000100010011;
ROM[8423] <= 32'b00000100000000000000001110010011;
ROM[8424] <= 32'b00000000011101100010000000100011;
ROM[8425] <= 32'b11111111110000010000000100010011;
ROM[8426] <= 32'b00000000000000010010001110000011;
ROM[8427] <= 32'b00000000000000111000001100010011;
ROM[8428] <= 32'b00000000000001100010001110000011;
ROM[8429] <= 32'b00000000110100110000010000110011;
ROM[8430] <= 32'b00000000011101000010000000100011;
ROM[8431] <= 32'b00000001110000000000001110010011;
ROM[8432] <= 32'b00000000011100010010000000100011;
ROM[8433] <= 32'b00000000010000010000000100010011;
ROM[8434] <= 32'b00000100100001101010001110000011;
ROM[8435] <= 32'b11111111110000010000000100010011;
ROM[8436] <= 32'b00000000000000010010010000000011;
ROM[8437] <= 32'b00000000011101000000001110110011;
ROM[8438] <= 32'b00000000011100010010000000100011;
ROM[8439] <= 32'b00000000010000010000000100010011;
ROM[8440] <= 32'b00001000000000000000001110010011;
ROM[8441] <= 32'b00000000011101100010000000100011;
ROM[8442] <= 32'b11111111110000010000000100010011;
ROM[8443] <= 32'b00000000000000010010001110000011;
ROM[8444] <= 32'b00000000000000111000001100010011;
ROM[8445] <= 32'b00000000000001100010001110000011;
ROM[8446] <= 32'b00000000110100110000010000110011;
ROM[8447] <= 32'b00000000011101000010000000100011;
ROM[8448] <= 32'b00000010000000000000001110010011;
ROM[8449] <= 32'b00000000011100010010000000100011;
ROM[8450] <= 32'b00000000010000010000000100010011;
ROM[8451] <= 32'b00000100100001101010001110000011;
ROM[8452] <= 32'b11111111110000010000000100010011;
ROM[8453] <= 32'b00000000000000010010010000000011;
ROM[8454] <= 32'b00000000011101000000001110110011;
ROM[8455] <= 32'b00000000011100010010000000100011;
ROM[8456] <= 32'b00000000010000010000000100010011;
ROM[8457] <= 32'b00010000000000000000001110010011;
ROM[8458] <= 32'b00000000011101100010000000100011;
ROM[8459] <= 32'b11111111110000010000000100010011;
ROM[8460] <= 32'b00000000000000010010001110000011;
ROM[8461] <= 32'b00000000000000111000001100010011;
ROM[8462] <= 32'b00000000000001100010001110000011;
ROM[8463] <= 32'b00000000110100110000010000110011;
ROM[8464] <= 32'b00000000011101000010000000100011;
ROM[8465] <= 32'b00000010010000000000001110010011;
ROM[8466] <= 32'b00000000011100010010000000100011;
ROM[8467] <= 32'b00000000010000010000000100010011;
ROM[8468] <= 32'b00000100100001101010001110000011;
ROM[8469] <= 32'b11111111110000010000000100010011;
ROM[8470] <= 32'b00000000000000010010010000000011;
ROM[8471] <= 32'b00000000011101000000001110110011;
ROM[8472] <= 32'b00000000011100010010000000100011;
ROM[8473] <= 32'b00000000010000010000000100010011;
ROM[8474] <= 32'b00100000000000000000001110010011;
ROM[8475] <= 32'b00000000011101100010000000100011;
ROM[8476] <= 32'b11111111110000010000000100010011;
ROM[8477] <= 32'b00000000000000010010001110000011;
ROM[8478] <= 32'b00000000000000111000001100010011;
ROM[8479] <= 32'b00000000000001100010001110000011;
ROM[8480] <= 32'b00000000110100110000010000110011;
ROM[8481] <= 32'b00000000011101000010000000100011;
ROM[8482] <= 32'b00000010100000000000001110010011;
ROM[8483] <= 32'b00000000011100010010000000100011;
ROM[8484] <= 32'b00000000010000010000000100010011;
ROM[8485] <= 32'b00000100100001101010001110000011;
ROM[8486] <= 32'b11111111110000010000000100010011;
ROM[8487] <= 32'b00000000000000010010010000000011;
ROM[8488] <= 32'b00000000011101000000001110110011;
ROM[8489] <= 32'b00000000011100010010000000100011;
ROM[8490] <= 32'b00000000010000010000000100010011;
ROM[8491] <= 32'b01000000000000000000001110010011;
ROM[8492] <= 32'b00000000011101100010000000100011;
ROM[8493] <= 32'b11111111110000010000000100010011;
ROM[8494] <= 32'b00000000000000010010001110000011;
ROM[8495] <= 32'b00000000000000111000001100010011;
ROM[8496] <= 32'b00000000000001100010001110000011;
ROM[8497] <= 32'b00000000110100110000010000110011;
ROM[8498] <= 32'b00000000011101000010000000100011;
ROM[8499] <= 32'b00000010110000000000001110010011;
ROM[8500] <= 32'b00000000011100010010000000100011;
ROM[8501] <= 32'b00000000010000010000000100010011;
ROM[8502] <= 32'b00000100100001101010001110000011;
ROM[8503] <= 32'b11111111110000010000000100010011;
ROM[8504] <= 32'b00000000000000010010010000000011;
ROM[8505] <= 32'b00000000011101000000001110110011;
ROM[8506] <= 32'b00000000011100010010000000100011;
ROM[8507] <= 32'b00000000010000010000000100010011;
ROM[8508] <= 32'b00000000000000000001001110110111;
ROM[8509] <= 32'b10000000000000111000001110010011;
ROM[8510] <= 32'b00000000011101100010000000100011;
ROM[8511] <= 32'b11111111110000010000000100010011;
ROM[8512] <= 32'b00000000000000010010001110000011;
ROM[8513] <= 32'b00000000000000111000001100010011;
ROM[8514] <= 32'b00000000000001100010001110000011;
ROM[8515] <= 32'b00000000110100110000010000110011;
ROM[8516] <= 32'b00000000011101000010000000100011;
ROM[8517] <= 32'b00000011000000000000001110010011;
ROM[8518] <= 32'b00000000011100010010000000100011;
ROM[8519] <= 32'b00000000010000010000000100010011;
ROM[8520] <= 32'b00000100100001101010001110000011;
ROM[8521] <= 32'b11111111110000010000000100010011;
ROM[8522] <= 32'b00000000000000010010010000000011;
ROM[8523] <= 32'b00000000011101000000001110110011;
ROM[8524] <= 32'b00000000011100010010000000100011;
ROM[8525] <= 32'b00000000010000010000000100010011;
ROM[8526] <= 32'b00000000000000000001001110110111;
ROM[8527] <= 32'b00000000000000111000001110010011;
ROM[8528] <= 32'b00000000011101100010000000100011;
ROM[8529] <= 32'b11111111110000010000000100010011;
ROM[8530] <= 32'b00000000000000010010001110000011;
ROM[8531] <= 32'b00000000000000111000001100010011;
ROM[8532] <= 32'b00000000000001100010001110000011;
ROM[8533] <= 32'b00000000110100110000010000110011;
ROM[8534] <= 32'b00000000011101000010000000100011;
ROM[8535] <= 32'b00000011010000000000001110010011;
ROM[8536] <= 32'b00000000011100010010000000100011;
ROM[8537] <= 32'b00000000010000010000000100010011;
ROM[8538] <= 32'b00000100100001101010001110000011;
ROM[8539] <= 32'b11111111110000010000000100010011;
ROM[8540] <= 32'b00000000000000010010010000000011;
ROM[8541] <= 32'b00000000011101000000001110110011;
ROM[8542] <= 32'b00000000011100010010000000100011;
ROM[8543] <= 32'b00000000010000010000000100010011;
ROM[8544] <= 32'b00000000000000000010001110110111;
ROM[8545] <= 32'b00000000000000111000001110010011;
ROM[8546] <= 32'b00000000011101100010000000100011;
ROM[8547] <= 32'b11111111110000010000000100010011;
ROM[8548] <= 32'b00000000000000010010001110000011;
ROM[8549] <= 32'b00000000000000111000001100010011;
ROM[8550] <= 32'b00000000000001100010001110000011;
ROM[8551] <= 32'b00000000110100110000010000110011;
ROM[8552] <= 32'b00000000011101000010000000100011;
ROM[8553] <= 32'b00000011100000000000001110010011;
ROM[8554] <= 32'b00000000011100010010000000100011;
ROM[8555] <= 32'b00000000010000010000000100010011;
ROM[8556] <= 32'b00000100100001101010001110000011;
ROM[8557] <= 32'b11111111110000010000000100010011;
ROM[8558] <= 32'b00000000000000010010010000000011;
ROM[8559] <= 32'b00000000011101000000001110110011;
ROM[8560] <= 32'b00000000011100010010000000100011;
ROM[8561] <= 32'b00000000010000010000000100010011;
ROM[8562] <= 32'b00000000000000000100001110110111;
ROM[8563] <= 32'b00000000000000111000001110010011;
ROM[8564] <= 32'b00000000011101100010000000100011;
ROM[8565] <= 32'b11111111110000010000000100010011;
ROM[8566] <= 32'b00000000000000010010001110000011;
ROM[8567] <= 32'b00000000000000111000001100010011;
ROM[8568] <= 32'b00000000000001100010001110000011;
ROM[8569] <= 32'b00000000110100110000010000110011;
ROM[8570] <= 32'b00000000011101000010000000100011;
ROM[8571] <= 32'b00000011110000000000001110010011;
ROM[8572] <= 32'b00000000011100010010000000100011;
ROM[8573] <= 32'b00000000010000010000000100010011;
ROM[8574] <= 32'b00000100100001101010001110000011;
ROM[8575] <= 32'b11111111110000010000000100010011;
ROM[8576] <= 32'b00000000000000010010010000000011;
ROM[8577] <= 32'b00000000011101000000001110110011;
ROM[8578] <= 32'b00000000011100010010000000100011;
ROM[8579] <= 32'b00000000010000010000000100010011;
ROM[8580] <= 32'b00000000000000000100001110110111;
ROM[8581] <= 32'b00000000000000111000001110010011;
ROM[8582] <= 32'b00000000011100010010000000100011;
ROM[8583] <= 32'b00000000010000010000000100010011;
ROM[8584] <= 32'b00000000000000000100001110110111;
ROM[8585] <= 32'b00000000000000111000001110010011;
ROM[8586] <= 32'b11111111110000010000000100010011;
ROM[8587] <= 32'b00000000000000010010010000000011;
ROM[8588] <= 32'b00000000011101000000001110110011;
ROM[8589] <= 32'b00000000011101100010000000100011;
ROM[8590] <= 32'b11111111110000010000000100010011;
ROM[8591] <= 32'b00000000000000010010001110000011;
ROM[8592] <= 32'b00000000000000111000001100010011;
ROM[8593] <= 32'b00000000000001100010001110000011;
ROM[8594] <= 32'b00000000110100110000010000110011;
ROM[8595] <= 32'b00000000011101000010000000100011;
ROM[8596] <= 32'b00000100000000000000001110010011;
ROM[8597] <= 32'b00000000011100010010000000100011;
ROM[8598] <= 32'b00000000010000010000000100010011;
ROM[8599] <= 32'b00000100100001101010001110000011;
ROM[8600] <= 32'b11111111110000010000000100010011;
ROM[8601] <= 32'b00000000000000010010010000000011;
ROM[8602] <= 32'b00000000011101000000001110110011;
ROM[8603] <= 32'b00000000011100010010000000100011;
ROM[8604] <= 32'b00000000010000010000000100010011;
ROM[8605] <= 32'b00000011110000000000001110010011;
ROM[8606] <= 32'b00000000011100010010000000100011;
ROM[8607] <= 32'b00000000010000010000000100010011;
ROM[8608] <= 32'b00000100100001101010001110000011;
ROM[8609] <= 32'b11111111110000010000000100010011;
ROM[8610] <= 32'b00000000000000010010010000000011;
ROM[8611] <= 32'b00000000011101000000001110110011;
ROM[8612] <= 32'b00000000000000111000001100010011;
ROM[8613] <= 32'b00000000110100110000010000110011;
ROM[8614] <= 32'b00000000000001000010001110000011;
ROM[8615] <= 32'b00000000011100010010000000100011;
ROM[8616] <= 32'b00000000010000010000000100010011;
ROM[8617] <= 32'b00000011110000000000001110010011;
ROM[8618] <= 32'b00000000011100010010000000100011;
ROM[8619] <= 32'b00000000010000010000000100010011;
ROM[8620] <= 32'b00000100100001101010001110000011;
ROM[8621] <= 32'b11111111110000010000000100010011;
ROM[8622] <= 32'b00000000000000010010010000000011;
ROM[8623] <= 32'b00000000011101000000001110110011;
ROM[8624] <= 32'b00000000000000111000001100010011;
ROM[8625] <= 32'b00000000110100110000010000110011;
ROM[8626] <= 32'b00000000000001000010001110000011;
ROM[8627] <= 32'b11111111110000010000000100010011;
ROM[8628] <= 32'b00000000000000010010010000000011;
ROM[8629] <= 32'b00000000011101000000001110110011;
ROM[8630] <= 32'b00000000011101100010000000100011;
ROM[8631] <= 32'b11111111110000010000000100010011;
ROM[8632] <= 32'b00000000000000010010001110000011;
ROM[8633] <= 32'b00000000000000111000001100010011;
ROM[8634] <= 32'b00000000000001100010001110000011;
ROM[8635] <= 32'b00000000110100110000010000110011;
ROM[8636] <= 32'b00000000011101000010000000100011;
ROM[8637] <= 32'b00000100010000000000001110010011;
ROM[8638] <= 32'b00000000011100010010000000100011;
ROM[8639] <= 32'b00000000010000010000000100010011;
ROM[8640] <= 32'b00000100100001101010001110000011;
ROM[8641] <= 32'b11111111110000010000000100010011;
ROM[8642] <= 32'b00000000000000010010010000000011;
ROM[8643] <= 32'b00000000011101000000001110110011;
ROM[8644] <= 32'b00000000011100010010000000100011;
ROM[8645] <= 32'b00000000010000010000000100010011;
ROM[8646] <= 32'b00000100000000000000001110010011;
ROM[8647] <= 32'b00000000011100010010000000100011;
ROM[8648] <= 32'b00000000010000010000000100010011;
ROM[8649] <= 32'b00000100100001101010001110000011;
ROM[8650] <= 32'b11111111110000010000000100010011;
ROM[8651] <= 32'b00000000000000010010010000000011;
ROM[8652] <= 32'b00000000011101000000001110110011;
ROM[8653] <= 32'b00000000000000111000001100010011;
ROM[8654] <= 32'b00000000110100110000010000110011;
ROM[8655] <= 32'b00000000000001000010001110000011;
ROM[8656] <= 32'b00000000011100010010000000100011;
ROM[8657] <= 32'b00000000010000010000000100010011;
ROM[8658] <= 32'b00000100000000000000001110010011;
ROM[8659] <= 32'b00000000011100010010000000100011;
ROM[8660] <= 32'b00000000010000010000000100010011;
ROM[8661] <= 32'b00000100100001101010001110000011;
ROM[8662] <= 32'b11111111110000010000000100010011;
ROM[8663] <= 32'b00000000000000010010010000000011;
ROM[8664] <= 32'b00000000011101000000001110110011;
ROM[8665] <= 32'b00000000000000111000001100010011;
ROM[8666] <= 32'b00000000110100110000010000110011;
ROM[8667] <= 32'b00000000000001000010001110000011;
ROM[8668] <= 32'b11111111110000010000000100010011;
ROM[8669] <= 32'b00000000000000010010010000000011;
ROM[8670] <= 32'b00000000011101000000001110110011;
ROM[8671] <= 32'b00000000011101100010000000100011;
ROM[8672] <= 32'b11111111110000010000000100010011;
ROM[8673] <= 32'b00000000000000010010001110000011;
ROM[8674] <= 32'b00000000000000111000001100010011;
ROM[8675] <= 32'b00000000000001100010001110000011;
ROM[8676] <= 32'b00000000110100110000010000110011;
ROM[8677] <= 32'b00000000011101000010000000100011;
ROM[8678] <= 32'b00000100100000000000001110010011;
ROM[8679] <= 32'b00000000011100010010000000100011;
ROM[8680] <= 32'b00000000010000010000000100010011;
ROM[8681] <= 32'b00000100100001101010001110000011;
ROM[8682] <= 32'b11111111110000010000000100010011;
ROM[8683] <= 32'b00000000000000010010010000000011;
ROM[8684] <= 32'b00000000011101000000001110110011;
ROM[8685] <= 32'b00000000011100010010000000100011;
ROM[8686] <= 32'b00000000010000010000000100010011;
ROM[8687] <= 32'b00000100010000000000001110010011;
ROM[8688] <= 32'b00000000011100010010000000100011;
ROM[8689] <= 32'b00000000010000010000000100010011;
ROM[8690] <= 32'b00000100100001101010001110000011;
ROM[8691] <= 32'b11111111110000010000000100010011;
ROM[8692] <= 32'b00000000000000010010010000000011;
ROM[8693] <= 32'b00000000011101000000001110110011;
ROM[8694] <= 32'b00000000000000111000001100010011;
ROM[8695] <= 32'b00000000110100110000010000110011;
ROM[8696] <= 32'b00000000000001000010001110000011;
ROM[8697] <= 32'b00000000011100010010000000100011;
ROM[8698] <= 32'b00000000010000010000000100010011;
ROM[8699] <= 32'b00000100010000000000001110010011;
ROM[8700] <= 32'b00000000011100010010000000100011;
ROM[8701] <= 32'b00000000010000010000000100010011;
ROM[8702] <= 32'b00000100100001101010001110000011;
ROM[8703] <= 32'b11111111110000010000000100010011;
ROM[8704] <= 32'b00000000000000010010010000000011;
ROM[8705] <= 32'b00000000011101000000001110110011;
ROM[8706] <= 32'b00000000000000111000001100010011;
ROM[8707] <= 32'b00000000110100110000010000110011;
ROM[8708] <= 32'b00000000000001000010001110000011;
ROM[8709] <= 32'b11111111110000010000000100010011;
ROM[8710] <= 32'b00000000000000010010010000000011;
ROM[8711] <= 32'b00000000011101000000001110110011;
ROM[8712] <= 32'b00000000011101100010000000100011;
ROM[8713] <= 32'b11111111110000010000000100010011;
ROM[8714] <= 32'b00000000000000010010001110000011;
ROM[8715] <= 32'b00000000000000111000001100010011;
ROM[8716] <= 32'b00000000000001100010001110000011;
ROM[8717] <= 32'b00000000110100110000010000110011;
ROM[8718] <= 32'b00000000011101000010000000100011;
ROM[8719] <= 32'b00000100110000000000001110010011;
ROM[8720] <= 32'b00000000011100010010000000100011;
ROM[8721] <= 32'b00000000010000010000000100010011;
ROM[8722] <= 32'b00000100100001101010001110000011;
ROM[8723] <= 32'b11111111110000010000000100010011;
ROM[8724] <= 32'b00000000000000010010010000000011;
ROM[8725] <= 32'b00000000011101000000001110110011;
ROM[8726] <= 32'b00000000011100010010000000100011;
ROM[8727] <= 32'b00000000010000010000000100010011;
ROM[8728] <= 32'b00000100100000000000001110010011;
ROM[8729] <= 32'b00000000011100010010000000100011;
ROM[8730] <= 32'b00000000010000010000000100010011;
ROM[8731] <= 32'b00000100100001101010001110000011;
ROM[8732] <= 32'b11111111110000010000000100010011;
ROM[8733] <= 32'b00000000000000010010010000000011;
ROM[8734] <= 32'b00000000011101000000001110110011;
ROM[8735] <= 32'b00000000000000111000001100010011;
ROM[8736] <= 32'b00000000110100110000010000110011;
ROM[8737] <= 32'b00000000000001000010001110000011;
ROM[8738] <= 32'b00000000011100010010000000100011;
ROM[8739] <= 32'b00000000010000010000000100010011;
ROM[8740] <= 32'b00000100100000000000001110010011;
ROM[8741] <= 32'b00000000011100010010000000100011;
ROM[8742] <= 32'b00000000010000010000000100010011;
ROM[8743] <= 32'b00000100100001101010001110000011;
ROM[8744] <= 32'b11111111110000010000000100010011;
ROM[8745] <= 32'b00000000000000010010010000000011;
ROM[8746] <= 32'b00000000011101000000001110110011;
ROM[8747] <= 32'b00000000000000111000001100010011;
ROM[8748] <= 32'b00000000110100110000010000110011;
ROM[8749] <= 32'b00000000000001000010001110000011;
ROM[8750] <= 32'b11111111110000010000000100010011;
ROM[8751] <= 32'b00000000000000010010010000000011;
ROM[8752] <= 32'b00000000011101000000001110110011;
ROM[8753] <= 32'b00000000011101100010000000100011;
ROM[8754] <= 32'b11111111110000010000000100010011;
ROM[8755] <= 32'b00000000000000010010001110000011;
ROM[8756] <= 32'b00000000000000111000001100010011;
ROM[8757] <= 32'b00000000000001100010001110000011;
ROM[8758] <= 32'b00000000110100110000010000110011;
ROM[8759] <= 32'b00000000011101000010000000100011;
ROM[8760] <= 32'b00000101000000000000001110010011;
ROM[8761] <= 32'b00000000011100010010000000100011;
ROM[8762] <= 32'b00000000010000010000000100010011;
ROM[8763] <= 32'b00000100100001101010001110000011;
ROM[8764] <= 32'b11111111110000010000000100010011;
ROM[8765] <= 32'b00000000000000010010010000000011;
ROM[8766] <= 32'b00000000011101000000001110110011;
ROM[8767] <= 32'b00000000011100010010000000100011;
ROM[8768] <= 32'b00000000010000010000000100010011;
ROM[8769] <= 32'b00000100110000000000001110010011;
ROM[8770] <= 32'b00000000011100010010000000100011;
ROM[8771] <= 32'b00000000010000010000000100010011;
ROM[8772] <= 32'b00000100100001101010001110000011;
ROM[8773] <= 32'b11111111110000010000000100010011;
ROM[8774] <= 32'b00000000000000010010010000000011;
ROM[8775] <= 32'b00000000011101000000001110110011;
ROM[8776] <= 32'b00000000000000111000001100010011;
ROM[8777] <= 32'b00000000110100110000010000110011;
ROM[8778] <= 32'b00000000000001000010001110000011;
ROM[8779] <= 32'b00000000011100010010000000100011;
ROM[8780] <= 32'b00000000010000010000000100010011;
ROM[8781] <= 32'b00000100110000000000001110010011;
ROM[8782] <= 32'b00000000011100010010000000100011;
ROM[8783] <= 32'b00000000010000010000000100010011;
ROM[8784] <= 32'b00000100100001101010001110000011;
ROM[8785] <= 32'b11111111110000010000000100010011;
ROM[8786] <= 32'b00000000000000010010010000000011;
ROM[8787] <= 32'b00000000011101000000001110110011;
ROM[8788] <= 32'b00000000000000111000001100010011;
ROM[8789] <= 32'b00000000110100110000010000110011;
ROM[8790] <= 32'b00000000000001000010001110000011;
ROM[8791] <= 32'b11111111110000010000000100010011;
ROM[8792] <= 32'b00000000000000010010010000000011;
ROM[8793] <= 32'b00000000011101000000001110110011;
ROM[8794] <= 32'b00000000011101100010000000100011;
ROM[8795] <= 32'b11111111110000010000000100010011;
ROM[8796] <= 32'b00000000000000010010001110000011;
ROM[8797] <= 32'b00000000000000111000001100010011;
ROM[8798] <= 32'b00000000000001100010001110000011;
ROM[8799] <= 32'b00000000110100110000010000110011;
ROM[8800] <= 32'b00000000011101000010000000100011;
ROM[8801] <= 32'b00000101010000000000001110010011;
ROM[8802] <= 32'b00000000011100010010000000100011;
ROM[8803] <= 32'b00000000010000010000000100010011;
ROM[8804] <= 32'b00000100100001101010001110000011;
ROM[8805] <= 32'b11111111110000010000000100010011;
ROM[8806] <= 32'b00000000000000010010010000000011;
ROM[8807] <= 32'b00000000011101000000001110110011;
ROM[8808] <= 32'b00000000011100010010000000100011;
ROM[8809] <= 32'b00000000010000010000000100010011;
ROM[8810] <= 32'b00000101000000000000001110010011;
ROM[8811] <= 32'b00000000011100010010000000100011;
ROM[8812] <= 32'b00000000010000010000000100010011;
ROM[8813] <= 32'b00000100100001101010001110000011;
ROM[8814] <= 32'b11111111110000010000000100010011;
ROM[8815] <= 32'b00000000000000010010010000000011;
ROM[8816] <= 32'b00000000011101000000001110110011;
ROM[8817] <= 32'b00000000000000111000001100010011;
ROM[8818] <= 32'b00000000110100110000010000110011;
ROM[8819] <= 32'b00000000000001000010001110000011;
ROM[8820] <= 32'b00000000011100010010000000100011;
ROM[8821] <= 32'b00000000010000010000000100010011;
ROM[8822] <= 32'b00000101000000000000001110010011;
ROM[8823] <= 32'b00000000011100010010000000100011;
ROM[8824] <= 32'b00000000010000010000000100010011;
ROM[8825] <= 32'b00000100100001101010001110000011;
ROM[8826] <= 32'b11111111110000010000000100010011;
ROM[8827] <= 32'b00000000000000010010010000000011;
ROM[8828] <= 32'b00000000011101000000001110110011;
ROM[8829] <= 32'b00000000000000111000001100010011;
ROM[8830] <= 32'b00000000110100110000010000110011;
ROM[8831] <= 32'b00000000000001000010001110000011;
ROM[8832] <= 32'b11111111110000010000000100010011;
ROM[8833] <= 32'b00000000000000010010010000000011;
ROM[8834] <= 32'b00000000011101000000001110110011;
ROM[8835] <= 32'b00000000011101100010000000100011;
ROM[8836] <= 32'b11111111110000010000000100010011;
ROM[8837] <= 32'b00000000000000010010001110000011;
ROM[8838] <= 32'b00000000000000111000001100010011;
ROM[8839] <= 32'b00000000000001100010001110000011;
ROM[8840] <= 32'b00000000110100110000010000110011;
ROM[8841] <= 32'b00000000011101000010000000100011;
ROM[8842] <= 32'b00000101100000000000001110010011;
ROM[8843] <= 32'b00000000011100010010000000100011;
ROM[8844] <= 32'b00000000010000010000000100010011;
ROM[8845] <= 32'b00000100100001101010001110000011;
ROM[8846] <= 32'b11111111110000010000000100010011;
ROM[8847] <= 32'b00000000000000010010010000000011;
ROM[8848] <= 32'b00000000011101000000001110110011;
ROM[8849] <= 32'b00000000011100010010000000100011;
ROM[8850] <= 32'b00000000010000010000000100010011;
ROM[8851] <= 32'b00000101010000000000001110010011;
ROM[8852] <= 32'b00000000011100010010000000100011;
ROM[8853] <= 32'b00000000010000010000000100010011;
ROM[8854] <= 32'b00000100100001101010001110000011;
ROM[8855] <= 32'b11111111110000010000000100010011;
ROM[8856] <= 32'b00000000000000010010010000000011;
ROM[8857] <= 32'b00000000011101000000001110110011;
ROM[8858] <= 32'b00000000000000111000001100010011;
ROM[8859] <= 32'b00000000110100110000010000110011;
ROM[8860] <= 32'b00000000000001000010001110000011;
ROM[8861] <= 32'b00000000011100010010000000100011;
ROM[8862] <= 32'b00000000010000010000000100010011;
ROM[8863] <= 32'b00000101010000000000001110010011;
ROM[8864] <= 32'b00000000011100010010000000100011;
ROM[8865] <= 32'b00000000010000010000000100010011;
ROM[8866] <= 32'b00000100100001101010001110000011;
ROM[8867] <= 32'b11111111110000010000000100010011;
ROM[8868] <= 32'b00000000000000010010010000000011;
ROM[8869] <= 32'b00000000011101000000001110110011;
ROM[8870] <= 32'b00000000000000111000001100010011;
ROM[8871] <= 32'b00000000110100110000010000110011;
ROM[8872] <= 32'b00000000000001000010001110000011;
ROM[8873] <= 32'b11111111110000010000000100010011;
ROM[8874] <= 32'b00000000000000010010010000000011;
ROM[8875] <= 32'b00000000011101000000001110110011;
ROM[8876] <= 32'b00000000011101100010000000100011;
ROM[8877] <= 32'b11111111110000010000000100010011;
ROM[8878] <= 32'b00000000000000010010001110000011;
ROM[8879] <= 32'b00000000000000111000001100010011;
ROM[8880] <= 32'b00000000000001100010001110000011;
ROM[8881] <= 32'b00000000110100110000010000110011;
ROM[8882] <= 32'b00000000011101000010000000100011;
ROM[8883] <= 32'b00000101110000000000001110010011;
ROM[8884] <= 32'b00000000011100010010000000100011;
ROM[8885] <= 32'b00000000010000010000000100010011;
ROM[8886] <= 32'b00000100100001101010001110000011;
ROM[8887] <= 32'b11111111110000010000000100010011;
ROM[8888] <= 32'b00000000000000010010010000000011;
ROM[8889] <= 32'b00000000011101000000001110110011;
ROM[8890] <= 32'b00000000011100010010000000100011;
ROM[8891] <= 32'b00000000010000010000000100010011;
ROM[8892] <= 32'b00000101100000000000001110010011;
ROM[8893] <= 32'b00000000011100010010000000100011;
ROM[8894] <= 32'b00000000010000010000000100010011;
ROM[8895] <= 32'b00000100100001101010001110000011;
ROM[8896] <= 32'b11111111110000010000000100010011;
ROM[8897] <= 32'b00000000000000010010010000000011;
ROM[8898] <= 32'b00000000011101000000001110110011;
ROM[8899] <= 32'b00000000000000111000001100010011;
ROM[8900] <= 32'b00000000110100110000010000110011;
ROM[8901] <= 32'b00000000000001000010001110000011;
ROM[8902] <= 32'b00000000011100010010000000100011;
ROM[8903] <= 32'b00000000010000010000000100010011;
ROM[8904] <= 32'b00000101100000000000001110010011;
ROM[8905] <= 32'b00000000011100010010000000100011;
ROM[8906] <= 32'b00000000010000010000000100010011;
ROM[8907] <= 32'b00000100100001101010001110000011;
ROM[8908] <= 32'b11111111110000010000000100010011;
ROM[8909] <= 32'b00000000000000010010010000000011;
ROM[8910] <= 32'b00000000011101000000001110110011;
ROM[8911] <= 32'b00000000000000111000001100010011;
ROM[8912] <= 32'b00000000110100110000010000110011;
ROM[8913] <= 32'b00000000000001000010001110000011;
ROM[8914] <= 32'b11111111110000010000000100010011;
ROM[8915] <= 32'b00000000000000010010010000000011;
ROM[8916] <= 32'b00000000011101000000001110110011;
ROM[8917] <= 32'b00000000011101100010000000100011;
ROM[8918] <= 32'b11111111110000010000000100010011;
ROM[8919] <= 32'b00000000000000010010001110000011;
ROM[8920] <= 32'b00000000000000111000001100010011;
ROM[8921] <= 32'b00000000000001100010001110000011;
ROM[8922] <= 32'b00000000110100110000010000110011;
ROM[8923] <= 32'b00000000011101000010000000100011;
ROM[8924] <= 32'b00000110000000000000001110010011;
ROM[8925] <= 32'b00000000011100010010000000100011;
ROM[8926] <= 32'b00000000010000010000000100010011;
ROM[8927] <= 32'b00000100100001101010001110000011;
ROM[8928] <= 32'b11111111110000010000000100010011;
ROM[8929] <= 32'b00000000000000010010010000000011;
ROM[8930] <= 32'b00000000011101000000001110110011;
ROM[8931] <= 32'b00000000011100010010000000100011;
ROM[8932] <= 32'b00000000010000010000000100010011;
ROM[8933] <= 32'b00000101110000000000001110010011;
ROM[8934] <= 32'b00000000011100010010000000100011;
ROM[8935] <= 32'b00000000010000010000000100010011;
ROM[8936] <= 32'b00000100100001101010001110000011;
ROM[8937] <= 32'b11111111110000010000000100010011;
ROM[8938] <= 32'b00000000000000010010010000000011;
ROM[8939] <= 32'b00000000011101000000001110110011;
ROM[8940] <= 32'b00000000000000111000001100010011;
ROM[8941] <= 32'b00000000110100110000010000110011;
ROM[8942] <= 32'b00000000000001000010001110000011;
ROM[8943] <= 32'b00000000011100010010000000100011;
ROM[8944] <= 32'b00000000010000010000000100010011;
ROM[8945] <= 32'b00000101110000000000001110010011;
ROM[8946] <= 32'b00000000011100010010000000100011;
ROM[8947] <= 32'b00000000010000010000000100010011;
ROM[8948] <= 32'b00000100100001101010001110000011;
ROM[8949] <= 32'b11111111110000010000000100010011;
ROM[8950] <= 32'b00000000000000010010010000000011;
ROM[8951] <= 32'b00000000011101000000001110110011;
ROM[8952] <= 32'b00000000000000111000001100010011;
ROM[8953] <= 32'b00000000110100110000010000110011;
ROM[8954] <= 32'b00000000000001000010001110000011;
ROM[8955] <= 32'b11111111110000010000000100010011;
ROM[8956] <= 32'b00000000000000010010010000000011;
ROM[8957] <= 32'b00000000011101000000001110110011;
ROM[8958] <= 32'b00000000011101100010000000100011;
ROM[8959] <= 32'b11111111110000010000000100010011;
ROM[8960] <= 32'b00000000000000010010001110000011;
ROM[8961] <= 32'b00000000000000111000001100010011;
ROM[8962] <= 32'b00000000000001100010001110000011;
ROM[8963] <= 32'b00000000110100110000010000110011;
ROM[8964] <= 32'b00000000011101000010000000100011;
ROM[8965] <= 32'b00000110010000000000001110010011;
ROM[8966] <= 32'b00000000011100010010000000100011;
ROM[8967] <= 32'b00000000010000010000000100010011;
ROM[8968] <= 32'b00000100100001101010001110000011;
ROM[8969] <= 32'b11111111110000010000000100010011;
ROM[8970] <= 32'b00000000000000010010010000000011;
ROM[8971] <= 32'b00000000011101000000001110110011;
ROM[8972] <= 32'b00000000011100010010000000100011;
ROM[8973] <= 32'b00000000010000010000000100010011;
ROM[8974] <= 32'b00000110000000000000001110010011;
ROM[8975] <= 32'b00000000011100010010000000100011;
ROM[8976] <= 32'b00000000010000010000000100010011;
ROM[8977] <= 32'b00000100100001101010001110000011;
ROM[8978] <= 32'b11111111110000010000000100010011;
ROM[8979] <= 32'b00000000000000010010010000000011;
ROM[8980] <= 32'b00000000011101000000001110110011;
ROM[8981] <= 32'b00000000000000111000001100010011;
ROM[8982] <= 32'b00000000110100110000010000110011;
ROM[8983] <= 32'b00000000000001000010001110000011;
ROM[8984] <= 32'b00000000011100010010000000100011;
ROM[8985] <= 32'b00000000010000010000000100010011;
ROM[8986] <= 32'b00000110000000000000001110010011;
ROM[8987] <= 32'b00000000011100010010000000100011;
ROM[8988] <= 32'b00000000010000010000000100010011;
ROM[8989] <= 32'b00000100100001101010001110000011;
ROM[8990] <= 32'b11111111110000010000000100010011;
ROM[8991] <= 32'b00000000000000010010010000000011;
ROM[8992] <= 32'b00000000011101000000001110110011;
ROM[8993] <= 32'b00000000000000111000001100010011;
ROM[8994] <= 32'b00000000110100110000010000110011;
ROM[8995] <= 32'b00000000000001000010001110000011;
ROM[8996] <= 32'b11111111110000010000000100010011;
ROM[8997] <= 32'b00000000000000010010010000000011;
ROM[8998] <= 32'b00000000011101000000001110110011;
ROM[8999] <= 32'b00000000011101100010000000100011;
ROM[9000] <= 32'b11111111110000010000000100010011;
ROM[9001] <= 32'b00000000000000010010001110000011;
ROM[9002] <= 32'b00000000000000111000001100010011;
ROM[9003] <= 32'b00000000000001100010001110000011;
ROM[9004] <= 32'b00000000110100110000010000110011;
ROM[9005] <= 32'b00000000011101000010000000100011;
ROM[9006] <= 32'b00000110100000000000001110010011;
ROM[9007] <= 32'b00000000011100010010000000100011;
ROM[9008] <= 32'b00000000010000010000000100010011;
ROM[9009] <= 32'b00000100100001101010001110000011;
ROM[9010] <= 32'b11111111110000010000000100010011;
ROM[9011] <= 32'b00000000000000010010010000000011;
ROM[9012] <= 32'b00000000011101000000001110110011;
ROM[9013] <= 32'b00000000011100010010000000100011;
ROM[9014] <= 32'b00000000010000010000000100010011;
ROM[9015] <= 32'b00000110010000000000001110010011;
ROM[9016] <= 32'b00000000011100010010000000100011;
ROM[9017] <= 32'b00000000010000010000000100010011;
ROM[9018] <= 32'b00000100100001101010001110000011;
ROM[9019] <= 32'b11111111110000010000000100010011;
ROM[9020] <= 32'b00000000000000010010010000000011;
ROM[9021] <= 32'b00000000011101000000001110110011;
ROM[9022] <= 32'b00000000000000111000001100010011;
ROM[9023] <= 32'b00000000110100110000010000110011;
ROM[9024] <= 32'b00000000000001000010001110000011;
ROM[9025] <= 32'b00000000011100010010000000100011;
ROM[9026] <= 32'b00000000010000010000000100010011;
ROM[9027] <= 32'b00000110010000000000001110010011;
ROM[9028] <= 32'b00000000011100010010000000100011;
ROM[9029] <= 32'b00000000010000010000000100010011;
ROM[9030] <= 32'b00000100100001101010001110000011;
ROM[9031] <= 32'b11111111110000010000000100010011;
ROM[9032] <= 32'b00000000000000010010010000000011;
ROM[9033] <= 32'b00000000011101000000001110110011;
ROM[9034] <= 32'b00000000000000111000001100010011;
ROM[9035] <= 32'b00000000110100110000010000110011;
ROM[9036] <= 32'b00000000000001000010001110000011;
ROM[9037] <= 32'b11111111110000010000000100010011;
ROM[9038] <= 32'b00000000000000010010010000000011;
ROM[9039] <= 32'b00000000011101000000001110110011;
ROM[9040] <= 32'b00000000011101100010000000100011;
ROM[9041] <= 32'b11111111110000010000000100010011;
ROM[9042] <= 32'b00000000000000010010001110000011;
ROM[9043] <= 32'b00000000000000111000001100010011;
ROM[9044] <= 32'b00000000000001100010001110000011;
ROM[9045] <= 32'b00000000110100110000010000110011;
ROM[9046] <= 32'b00000000011101000010000000100011;
ROM[9047] <= 32'b00000110110000000000001110010011;
ROM[9048] <= 32'b00000000011100010010000000100011;
ROM[9049] <= 32'b00000000010000010000000100010011;
ROM[9050] <= 32'b00000100100001101010001110000011;
ROM[9051] <= 32'b11111111110000010000000100010011;
ROM[9052] <= 32'b00000000000000010010010000000011;
ROM[9053] <= 32'b00000000011101000000001110110011;
ROM[9054] <= 32'b00000000011100010010000000100011;
ROM[9055] <= 32'b00000000010000010000000100010011;
ROM[9056] <= 32'b00000110100000000000001110010011;
ROM[9057] <= 32'b00000000011100010010000000100011;
ROM[9058] <= 32'b00000000010000010000000100010011;
ROM[9059] <= 32'b00000100100001101010001110000011;
ROM[9060] <= 32'b11111111110000010000000100010011;
ROM[9061] <= 32'b00000000000000010010010000000011;
ROM[9062] <= 32'b00000000011101000000001110110011;
ROM[9063] <= 32'b00000000000000111000001100010011;
ROM[9064] <= 32'b00000000110100110000010000110011;
ROM[9065] <= 32'b00000000000001000010001110000011;
ROM[9066] <= 32'b00000000011100010010000000100011;
ROM[9067] <= 32'b00000000010000010000000100010011;
ROM[9068] <= 32'b00000110100000000000001110010011;
ROM[9069] <= 32'b00000000011100010010000000100011;
ROM[9070] <= 32'b00000000010000010000000100010011;
ROM[9071] <= 32'b00000100100001101010001110000011;
ROM[9072] <= 32'b11111111110000010000000100010011;
ROM[9073] <= 32'b00000000000000010010010000000011;
ROM[9074] <= 32'b00000000011101000000001110110011;
ROM[9075] <= 32'b00000000000000111000001100010011;
ROM[9076] <= 32'b00000000110100110000010000110011;
ROM[9077] <= 32'b00000000000001000010001110000011;
ROM[9078] <= 32'b11111111110000010000000100010011;
ROM[9079] <= 32'b00000000000000010010010000000011;
ROM[9080] <= 32'b00000000011101000000001110110011;
ROM[9081] <= 32'b00000000011101100010000000100011;
ROM[9082] <= 32'b11111111110000010000000100010011;
ROM[9083] <= 32'b00000000000000010010001110000011;
ROM[9084] <= 32'b00000000000000111000001100010011;
ROM[9085] <= 32'b00000000000001100010001110000011;
ROM[9086] <= 32'b00000000110100110000010000110011;
ROM[9087] <= 32'b00000000011101000010000000100011;
ROM[9088] <= 32'b00000111000000000000001110010011;
ROM[9089] <= 32'b00000000011100010010000000100011;
ROM[9090] <= 32'b00000000010000010000000100010011;
ROM[9091] <= 32'b00000100100001101010001110000011;
ROM[9092] <= 32'b11111111110000010000000100010011;
ROM[9093] <= 32'b00000000000000010010010000000011;
ROM[9094] <= 32'b00000000011101000000001110110011;
ROM[9095] <= 32'b00000000011100010010000000100011;
ROM[9096] <= 32'b00000000010000010000000100010011;
ROM[9097] <= 32'b00000110110000000000001110010011;
ROM[9098] <= 32'b00000000011100010010000000100011;
ROM[9099] <= 32'b00000000010000010000000100010011;
ROM[9100] <= 32'b00000100100001101010001110000011;
ROM[9101] <= 32'b11111111110000010000000100010011;
ROM[9102] <= 32'b00000000000000010010010000000011;
ROM[9103] <= 32'b00000000011101000000001110110011;
ROM[9104] <= 32'b00000000000000111000001100010011;
ROM[9105] <= 32'b00000000110100110000010000110011;
ROM[9106] <= 32'b00000000000001000010001110000011;
ROM[9107] <= 32'b00000000011100010010000000100011;
ROM[9108] <= 32'b00000000010000010000000100010011;
ROM[9109] <= 32'b00000110110000000000001110010011;
ROM[9110] <= 32'b00000000011100010010000000100011;
ROM[9111] <= 32'b00000000010000010000000100010011;
ROM[9112] <= 32'b00000100100001101010001110000011;
ROM[9113] <= 32'b11111111110000010000000100010011;
ROM[9114] <= 32'b00000000000000010010010000000011;
ROM[9115] <= 32'b00000000011101000000001110110011;
ROM[9116] <= 32'b00000000000000111000001100010011;
ROM[9117] <= 32'b00000000110100110000010000110011;
ROM[9118] <= 32'b00000000000001000010001110000011;
ROM[9119] <= 32'b11111111110000010000000100010011;
ROM[9120] <= 32'b00000000000000010010010000000011;
ROM[9121] <= 32'b00000000011101000000001110110011;
ROM[9122] <= 32'b00000000011101100010000000100011;
ROM[9123] <= 32'b11111111110000010000000100010011;
ROM[9124] <= 32'b00000000000000010010001110000011;
ROM[9125] <= 32'b00000000000000111000001100010011;
ROM[9126] <= 32'b00000000000001100010001110000011;
ROM[9127] <= 32'b00000000110100110000010000110011;
ROM[9128] <= 32'b00000000011101000010000000100011;
ROM[9129] <= 32'b00000111010000000000001110010011;
ROM[9130] <= 32'b00000000011100010010000000100011;
ROM[9131] <= 32'b00000000010000010000000100010011;
ROM[9132] <= 32'b00000100100001101010001110000011;
ROM[9133] <= 32'b11111111110000010000000100010011;
ROM[9134] <= 32'b00000000000000010010010000000011;
ROM[9135] <= 32'b00000000011101000000001110110011;
ROM[9136] <= 32'b00000000011100010010000000100011;
ROM[9137] <= 32'b00000000010000010000000100010011;
ROM[9138] <= 32'b00000111000000000000001110010011;
ROM[9139] <= 32'b00000000011100010010000000100011;
ROM[9140] <= 32'b00000000010000010000000100010011;
ROM[9141] <= 32'b00000100100001101010001110000011;
ROM[9142] <= 32'b11111111110000010000000100010011;
ROM[9143] <= 32'b00000000000000010010010000000011;
ROM[9144] <= 32'b00000000011101000000001110110011;
ROM[9145] <= 32'b00000000000000111000001100010011;
ROM[9146] <= 32'b00000000110100110000010000110011;
ROM[9147] <= 32'b00000000000001000010001110000011;
ROM[9148] <= 32'b00000000011100010010000000100011;
ROM[9149] <= 32'b00000000010000010000000100010011;
ROM[9150] <= 32'b00000111000000000000001110010011;
ROM[9151] <= 32'b00000000011100010010000000100011;
ROM[9152] <= 32'b00000000010000010000000100010011;
ROM[9153] <= 32'b00000100100001101010001110000011;
ROM[9154] <= 32'b11111111110000010000000100010011;
ROM[9155] <= 32'b00000000000000010010010000000011;
ROM[9156] <= 32'b00000000011101000000001110110011;
ROM[9157] <= 32'b00000000000000111000001100010011;
ROM[9158] <= 32'b00000000110100110000010000110011;
ROM[9159] <= 32'b00000000000001000010001110000011;
ROM[9160] <= 32'b11111111110000010000000100010011;
ROM[9161] <= 32'b00000000000000010010010000000011;
ROM[9162] <= 32'b00000000011101000000001110110011;
ROM[9163] <= 32'b00000000011101100010000000100011;
ROM[9164] <= 32'b11111111110000010000000100010011;
ROM[9165] <= 32'b00000000000000010010001110000011;
ROM[9166] <= 32'b00000000000000111000001100010011;
ROM[9167] <= 32'b00000000000001100010001110000011;
ROM[9168] <= 32'b00000000110100110000010000110011;
ROM[9169] <= 32'b00000000011101000010000000100011;
ROM[9170] <= 32'b00000111100000000000001110010011;
ROM[9171] <= 32'b00000000011100010010000000100011;
ROM[9172] <= 32'b00000000010000010000000100010011;
ROM[9173] <= 32'b00000100100001101010001110000011;
ROM[9174] <= 32'b11111111110000010000000100010011;
ROM[9175] <= 32'b00000000000000010010010000000011;
ROM[9176] <= 32'b00000000011101000000001110110011;
ROM[9177] <= 32'b00000000011100010010000000100011;
ROM[9178] <= 32'b00000000010000010000000100010011;
ROM[9179] <= 32'b00000111010000000000001110010011;
ROM[9180] <= 32'b00000000011100010010000000100011;
ROM[9181] <= 32'b00000000010000010000000100010011;
ROM[9182] <= 32'b00000100100001101010001110000011;
ROM[9183] <= 32'b11111111110000010000000100010011;
ROM[9184] <= 32'b00000000000000010010010000000011;
ROM[9185] <= 32'b00000000011101000000001110110011;
ROM[9186] <= 32'b00000000000000111000001100010011;
ROM[9187] <= 32'b00000000110100110000010000110011;
ROM[9188] <= 32'b00000000000001000010001110000011;
ROM[9189] <= 32'b00000000011100010010000000100011;
ROM[9190] <= 32'b00000000010000010000000100010011;
ROM[9191] <= 32'b00000111010000000000001110010011;
ROM[9192] <= 32'b00000000011100010010000000100011;
ROM[9193] <= 32'b00000000010000010000000100010011;
ROM[9194] <= 32'b00000100100001101010001110000011;
ROM[9195] <= 32'b11111111110000010000000100010011;
ROM[9196] <= 32'b00000000000000010010010000000011;
ROM[9197] <= 32'b00000000011101000000001110110011;
ROM[9198] <= 32'b00000000000000111000001100010011;
ROM[9199] <= 32'b00000000110100110000010000110011;
ROM[9200] <= 32'b00000000000001000010001110000011;
ROM[9201] <= 32'b11111111110000010000000100010011;
ROM[9202] <= 32'b00000000000000010010010000000011;
ROM[9203] <= 32'b00000000011101000000001110110011;
ROM[9204] <= 32'b00000000011101100010000000100011;
ROM[9205] <= 32'b11111111110000010000000100010011;
ROM[9206] <= 32'b00000000000000010010001110000011;
ROM[9207] <= 32'b00000000000000111000001100010011;
ROM[9208] <= 32'b00000000000001100010001110000011;
ROM[9209] <= 32'b00000000110100110000010000110011;
ROM[9210] <= 32'b00000000011101000010000000100011;
ROM[9211] <= 32'b00000111110000000000001110010011;
ROM[9212] <= 32'b00000000011100010010000000100011;
ROM[9213] <= 32'b00000000010000010000000100010011;
ROM[9214] <= 32'b00000100100001101010001110000011;
ROM[9215] <= 32'b11111111110000010000000100010011;
ROM[9216] <= 32'b00000000000000010010010000000011;
ROM[9217] <= 32'b00000000011101000000001110110011;
ROM[9218] <= 32'b00000000011100010010000000100011;
ROM[9219] <= 32'b00000000010000010000000100010011;
ROM[9220] <= 32'b00000111100000000000001110010011;
ROM[9221] <= 32'b00000000011100010010000000100011;
ROM[9222] <= 32'b00000000010000010000000100010011;
ROM[9223] <= 32'b00000100100001101010001110000011;
ROM[9224] <= 32'b11111111110000010000000100010011;
ROM[9225] <= 32'b00000000000000010010010000000011;
ROM[9226] <= 32'b00000000011101000000001110110011;
ROM[9227] <= 32'b00000000000000111000001100010011;
ROM[9228] <= 32'b00000000110100110000010000110011;
ROM[9229] <= 32'b00000000000001000010001110000011;
ROM[9230] <= 32'b00000000011100010010000000100011;
ROM[9231] <= 32'b00000000010000010000000100010011;
ROM[9232] <= 32'b00000111100000000000001110010011;
ROM[9233] <= 32'b00000000011100010010000000100011;
ROM[9234] <= 32'b00000000010000010000000100010011;
ROM[9235] <= 32'b00000100100001101010001110000011;
ROM[9236] <= 32'b11111111110000010000000100010011;
ROM[9237] <= 32'b00000000000000010010010000000011;
ROM[9238] <= 32'b00000000011101000000001110110011;
ROM[9239] <= 32'b00000000000000111000001100010011;
ROM[9240] <= 32'b00000000110100110000010000110011;
ROM[9241] <= 32'b00000000000001000010001110000011;
ROM[9242] <= 32'b11111111110000010000000100010011;
ROM[9243] <= 32'b00000000000000010010010000000011;
ROM[9244] <= 32'b00000000011101000000001110110011;
ROM[9245] <= 32'b00000000011101100010000000100011;
ROM[9246] <= 32'b11111111110000010000000100010011;
ROM[9247] <= 32'b00000000000000010010001110000011;
ROM[9248] <= 32'b00000000000000111000001100010011;
ROM[9249] <= 32'b00000000000001100010001110000011;
ROM[9250] <= 32'b00000000110100110000010000110011;
ROM[9251] <= 32'b00000000011101000010000000100011;
ROM[9252] <= 32'b00000000000000000000001110010011;
ROM[9253] <= 32'b00000000011100010010000000100011;
ROM[9254] <= 32'b00000000010000010000000100010011;
ROM[9255] <= 32'b00000001010000000000001110010011;
ROM[9256] <= 32'b01000000011100011000001110110011;
ROM[9257] <= 32'b00000000000000111010000010000011;
ROM[9258] <= 32'b11111111110000010000000100010011;
ROM[9259] <= 32'b00000000000000010010001110000011;
ROM[9260] <= 32'b00000000011100100010000000100011;
ROM[9261] <= 32'b00000000010000100000000100010011;
ROM[9262] <= 32'b00000001010000000000001110010011;
ROM[9263] <= 32'b01000000011100011000001110110011;
ROM[9264] <= 32'b00000000010000111010000110000011;
ROM[9265] <= 32'b00000000100000111010001000000011;
ROM[9266] <= 32'b00000000110000111010001010000011;
ROM[9267] <= 32'b00000001000000111010001100000011;
ROM[9268] <= 32'b00000000000000001000000011100111;
ROM[9269] <= 32'b00000000000000010010000000100011;
ROM[9270] <= 32'b00000000010000010000000100010011;
ROM[9271] <= 32'b00000000000000010010000000100011;
ROM[9272] <= 32'b00000000010000010000000100010011;
ROM[9273] <= 32'b00000000000000010010000000100011;
ROM[9274] <= 32'b00000000010000010000000100010011;
ROM[9275] <= 32'b00000000000000000000001110010011;
ROM[9276] <= 32'b00000000011100011010000000100011;
ROM[9277] <= 32'b00000000000000100010001110000011;
ROM[9278] <= 32'b00000000011100011010001000100011;
ROM[9279] <= 32'b00000000000000000000001110010011;
ROM[9280] <= 32'b00000000011100011010010000100011;
ROM[9281] <= 32'b00000000100000011010001110000011;
ROM[9282] <= 32'b00000000011100010010000000100011;
ROM[9283] <= 32'b00000000010000010000000100010011;
ROM[9284] <= 32'b00001000000000000000001110010011;
ROM[9285] <= 32'b11111111110000010000000100010011;
ROM[9286] <= 32'b00000000000000010010010000000011;
ROM[9287] <= 32'b00000000011101000010001110110011;
ROM[9288] <= 32'b01000000011100000000001110110011;
ROM[9289] <= 32'b00000000000100111000001110010011;
ROM[9290] <= 32'b00000000000000111000101001100011;
ROM[9291] <= 32'b00000000000000001001001110110111;
ROM[9292] <= 32'b00100010110000111000001110010011;
ROM[9293] <= 32'b00000000111000111000001110110011;
ROM[9294] <= 32'b00000000000000111000000011100111;
ROM[9295] <= 32'b00000000010000100010001110000011;
ROM[9296] <= 32'b00000000011100010010000000100011;
ROM[9297] <= 32'b00000000010000010000000100010011;
ROM[9298] <= 32'b00000000100000011010001110000011;
ROM[9299] <= 32'b00000000011100010010000000100011;
ROM[9300] <= 32'b00000000010000010000000100010011;
ROM[9301] <= 32'b00000100100001101010001110000011;
ROM[9302] <= 32'b11111111110000010000000100010011;
ROM[9303] <= 32'b00000000000000010010010000000011;
ROM[9304] <= 32'b00000000011101000000001110110011;
ROM[9305] <= 32'b00000000000000111000001100010011;
ROM[9306] <= 32'b00000000110100110000010000110011;
ROM[9307] <= 32'b00000000000001000010001110000011;
ROM[9308] <= 32'b11111111110000010000000100010011;
ROM[9309] <= 32'b00000000000000010010010000000011;
ROM[9310] <= 32'b00000000011101000111001110110011;
ROM[9311] <= 32'b00000000011100010010000000100011;
ROM[9312] <= 32'b00000000010000010000000100010011;
ROM[9313] <= 32'b00000000000000000000001110010011;
ROM[9314] <= 32'b11111111110000010000000100010011;
ROM[9315] <= 32'b00000000000000010010010000000011;
ROM[9316] <= 32'b00000000011101000010010010110011;
ROM[9317] <= 32'b00000000100000111010010100110011;
ROM[9318] <= 32'b00000000101001001000001110110011;
ROM[9319] <= 32'b00000000000100111000001110010011;
ROM[9320] <= 32'b00000000000100111111001110010011;
ROM[9321] <= 32'b01000000011100000000001110110011;
ROM[9322] <= 32'b00000000000100111000001110010011;
ROM[9323] <= 32'b00000000000000111000101001100011;
ROM[9324] <= 32'b00000000000000001001001110110111;
ROM[9325] <= 32'b00011100010000111000001110010011;
ROM[9326] <= 32'b00000000111000111000001110110011;
ROM[9327] <= 32'b00000000000000111000000011100111;
ROM[9328] <= 32'b00000010100000000000000011101111;
ROM[9329] <= 32'b00000000000000011010001110000011;
ROM[9330] <= 32'b00000000011100010010000000100011;
ROM[9331] <= 32'b00000000010000010000000100010011;
ROM[9332] <= 32'b00000000010000011010001110000011;
ROM[9333] <= 32'b11111111110000010000000100010011;
ROM[9334] <= 32'b00000000000000010010010000000011;
ROM[9335] <= 32'b00000000011101000000001110110011;
ROM[9336] <= 32'b00000000011100011010000000100011;
ROM[9337] <= 32'b00000000010000000000000011101111;
ROM[9338] <= 32'b00000000010000011010001110000011;
ROM[9339] <= 32'b00000000011100010010000000100011;
ROM[9340] <= 32'b00000000010000010000000100010011;
ROM[9341] <= 32'b00000000010000011010001110000011;
ROM[9342] <= 32'b11111111110000010000000100010011;
ROM[9343] <= 32'b00000000000000010010010000000011;
ROM[9344] <= 32'b00000000011101000000001110110011;
ROM[9345] <= 32'b00000000011100011010001000100011;
ROM[9346] <= 32'b00000000100000011010001110000011;
ROM[9347] <= 32'b00000000011100010010000000100011;
ROM[9348] <= 32'b00000000010000010000000100010011;
ROM[9349] <= 32'b00000000010000000000001110010011;
ROM[9350] <= 32'b11111111110000010000000100010011;
ROM[9351] <= 32'b00000000000000010010010000000011;
ROM[9352] <= 32'b00000000011101000000001110110011;
ROM[9353] <= 32'b00000000011100011010010000100011;
ROM[9354] <= 32'b11101101110111111111000011101111;
ROM[9355] <= 32'b00000000000000011010001110000011;
ROM[9356] <= 32'b00000000011100010010000000100011;
ROM[9357] <= 32'b00000000010000010000000100010011;
ROM[9358] <= 32'b00000001010000000000001110010011;
ROM[9359] <= 32'b01000000011100011000001110110011;
ROM[9360] <= 32'b00000000000000111010000010000011;
ROM[9361] <= 32'b11111111110000010000000100010011;
ROM[9362] <= 32'b00000000000000010010001110000011;
ROM[9363] <= 32'b00000000011100100010000000100011;
ROM[9364] <= 32'b00000000010000100000000100010011;
ROM[9365] <= 32'b00000001010000000000001110010011;
ROM[9366] <= 32'b01000000011100011000001110110011;
ROM[9367] <= 32'b00000000010000111010000110000011;
ROM[9368] <= 32'b00000000100000111010001000000011;
ROM[9369] <= 32'b00000000110000111010001010000011;
ROM[9370] <= 32'b00000001000000111010001100000011;
ROM[9371] <= 32'b00000000000000001000000011100111;
ROM[9372] <= 32'b00000000000000100010001110000011;
ROM[9373] <= 32'b00000000011100010010000000100011;
ROM[9374] <= 32'b00000000010000010000000100010011;
ROM[9375] <= 32'b00000000000000000000001110010011;
ROM[9376] <= 32'b11111111110000010000000100010011;
ROM[9377] <= 32'b00000000000000010010010000000011;
ROM[9378] <= 32'b00000000011101000010001110110011;
ROM[9379] <= 32'b00000000000000111000101001100011;
ROM[9380] <= 32'b00000000000000001001001110110111;
ROM[9381] <= 32'b00101010010000111000001110010011;
ROM[9382] <= 32'b00000000111000111000001110110011;
ROM[9383] <= 32'b00000000000000111000000011100111;
ROM[9384] <= 32'b00000001010000000000000011101111;
ROM[9385] <= 32'b00000000000000100010001110000011;
ROM[9386] <= 32'b01000000011100000000001110110011;
ROM[9387] <= 32'b00000000011100100010000000100011;
ROM[9388] <= 32'b00000000010000000000000011101111;
ROM[9389] <= 32'b00000000000000100010001110000011;
ROM[9390] <= 32'b00000000011100010010000000100011;
ROM[9391] <= 32'b00000000010000010000000100010011;
ROM[9392] <= 32'b00000001010000000000001110010011;
ROM[9393] <= 32'b01000000011100011000001110110011;
ROM[9394] <= 32'b00000000000000111010000010000011;
ROM[9395] <= 32'b11111111110000010000000100010011;
ROM[9396] <= 32'b00000000000000010010001110000011;
ROM[9397] <= 32'b00000000011100100010000000100011;
ROM[9398] <= 32'b00000000010000100000000100010011;
ROM[9399] <= 32'b00000001010000000000001110010011;
ROM[9400] <= 32'b01000000011100011000001110110011;
ROM[9401] <= 32'b00000000010000111010000110000011;
ROM[9402] <= 32'b00000000100000111010001000000011;
ROM[9403] <= 32'b00000000110000111010001010000011;
ROM[9404] <= 32'b00000001000000111010001100000011;
ROM[9405] <= 32'b00000000000000001000000011100111;
ROM[9406] <= 32'b00000000000000010010000000100011;
ROM[9407] <= 32'b00000000010000010000000100010011;
ROM[9408] <= 32'b00000000000000010010000000100011;
ROM[9409] <= 32'b00000000010000010000000100010011;
ROM[9410] <= 32'b00000000000000010010000000100011;
ROM[9411] <= 32'b00000000010000010000000100010011;
ROM[9412] <= 32'b00000000010000100010001110000011;
ROM[9413] <= 32'b00000000011100010010000000100011;
ROM[9414] <= 32'b00000000010000010000000100010011;
ROM[9415] <= 32'b00000000000000000000001110010011;
ROM[9416] <= 32'b11111111110000010000000100010011;
ROM[9417] <= 32'b00000000000000010010010000000011;
ROM[9418] <= 32'b00000000011101000010010010110011;
ROM[9419] <= 32'b00000000100000111010010100110011;
ROM[9420] <= 32'b00000000101001001000001110110011;
ROM[9421] <= 32'b00000000000100111000001110010011;
ROM[9422] <= 32'b00000000000100111111001110010011;
ROM[9423] <= 32'b00000000000000111000101001100011;
ROM[9424] <= 32'b00000000000000001001001110110111;
ROM[9425] <= 32'b00110101010000111000001110010011;
ROM[9426] <= 32'b00000000111000111000001110110011;
ROM[9427] <= 32'b00000000000000111000000011100111;
ROM[9428] <= 32'b00000101000000000000000011101111;
ROM[9429] <= 32'b00000000000100000000001110010011;
ROM[9430] <= 32'b01000000011100000000001110110011;
ROM[9431] <= 32'b00000000011100010010000000100011;
ROM[9432] <= 32'b00000000010000010000000100010011;
ROM[9433] <= 32'b00000001010000000000001110010011;
ROM[9434] <= 32'b01000000011100011000001110110011;
ROM[9435] <= 32'b00000000000000111010000010000011;
ROM[9436] <= 32'b11111111110000010000000100010011;
ROM[9437] <= 32'b00000000000000010010001110000011;
ROM[9438] <= 32'b00000000011100100010000000100011;
ROM[9439] <= 32'b00000000010000100000000100010011;
ROM[9440] <= 32'b00000001010000000000001110010011;
ROM[9441] <= 32'b01000000011100011000001110110011;
ROM[9442] <= 32'b00000000010000111010000110000011;
ROM[9443] <= 32'b00000000100000111010001000000011;
ROM[9444] <= 32'b00000000110000111010001010000011;
ROM[9445] <= 32'b00000001000000111010001100000011;
ROM[9446] <= 32'b00000000000000001000000011100111;
ROM[9447] <= 32'b00000000010000000000000011101111;
ROM[9448] <= 32'b00000000000000100010001110000011;
ROM[9449] <= 32'b00000000011100010010000000100011;
ROM[9450] <= 32'b00000000010000010000000100010011;
ROM[9451] <= 32'b00000000000000000000001110010011;
ROM[9452] <= 32'b11111111110000010000000100010011;
ROM[9453] <= 32'b00000000000000010010010000000011;
ROM[9454] <= 32'b00000000011101000010001110110011;
ROM[9455] <= 32'b00000000011100010010000000100011;
ROM[9456] <= 32'b00000000010000010000000100010011;
ROM[9457] <= 32'b00000000010000100010001110000011;
ROM[9458] <= 32'b00000000011100010010000000100011;
ROM[9459] <= 32'b00000000010000010000000100010011;
ROM[9460] <= 32'b00000000000000000000001110010011;
ROM[9461] <= 32'b11111111110000010000000100010011;
ROM[9462] <= 32'b00000000000000010010010000000011;
ROM[9463] <= 32'b00000000011101000010001110110011;
ROM[9464] <= 32'b11111111110000010000000100010011;
ROM[9465] <= 32'b00000000000000010010010000000011;
ROM[9466] <= 32'b00000000011101000010010010110011;
ROM[9467] <= 32'b00000000100000111010010100110011;
ROM[9468] <= 32'b00000000101001001000001110110011;
ROM[9469] <= 32'b00000000000100111000001110010011;
ROM[9470] <= 32'b00000000000100111111001110010011;
ROM[9471] <= 32'b01000000011100000000001110110011;
ROM[9472] <= 32'b00000000000100111000001110010011;
ROM[9473] <= 32'b00000000011100011010001000100011;
ROM[9474] <= 32'b00000000000000100010001110000011;
ROM[9475] <= 32'b00000000011100010010000000100011;
ROM[9476] <= 32'b00000000010000010000000100010011;
ROM[9477] <= 32'b00000000000000001001001110110111;
ROM[9478] <= 32'b01000110000000111000001110010011;
ROM[9479] <= 32'b00000000111000111000001110110011;
ROM[9480] <= 32'b00000000011100010010000000100011;
ROM[9481] <= 32'b00000000010000010000000100010011;
ROM[9482] <= 32'b00000000001100010010000000100011;
ROM[9483] <= 32'b00000000010000010000000100010011;
ROM[9484] <= 32'b00000000010000010010000000100011;
ROM[9485] <= 32'b00000000010000010000000100010011;
ROM[9486] <= 32'b00000000010100010010000000100011;
ROM[9487] <= 32'b00000000010000010000000100010011;
ROM[9488] <= 32'b00000000011000010010000000100011;
ROM[9489] <= 32'b00000000010000010000000100010011;
ROM[9490] <= 32'b00000001010000000000001110010011;
ROM[9491] <= 32'b00000000010000111000001110010011;
ROM[9492] <= 32'b01000000011100010000001110110011;
ROM[9493] <= 32'b00000000011100000000001000110011;
ROM[9494] <= 32'b00000000001000000000000110110011;
ROM[9495] <= 32'b11100001010111111111000011101111;
ROM[9496] <= 32'b11111111110000010000000100010011;
ROM[9497] <= 32'b00000000000000010010001110000011;
ROM[9498] <= 32'b00000000011100100010000000100011;
ROM[9499] <= 32'b00000000010000100010001110000011;
ROM[9500] <= 32'b00000000011100010010000000100011;
ROM[9501] <= 32'b00000000010000010000000100010011;
ROM[9502] <= 32'b00000000000000001001001110110111;
ROM[9503] <= 32'b01001100010000111000001110010011;
ROM[9504] <= 32'b00000000111000111000001110110011;
ROM[9505] <= 32'b00000000011100010010000000100011;
ROM[9506] <= 32'b00000000010000010000000100010011;
ROM[9507] <= 32'b00000000001100010010000000100011;
ROM[9508] <= 32'b00000000010000010000000100010011;
ROM[9509] <= 32'b00000000010000010010000000100011;
ROM[9510] <= 32'b00000000010000010000000100010011;
ROM[9511] <= 32'b00000000010100010010000000100011;
ROM[9512] <= 32'b00000000010000010000000100010011;
ROM[9513] <= 32'b00000000011000010010000000100011;
ROM[9514] <= 32'b00000000010000010000000100010011;
ROM[9515] <= 32'b00000001010000000000001110010011;
ROM[9516] <= 32'b00000000010000111000001110010011;
ROM[9517] <= 32'b01000000011100010000001110110011;
ROM[9518] <= 32'b00000000011100000000001000110011;
ROM[9519] <= 32'b00000000001000000000000110110011;
ROM[9520] <= 32'b11011011000111111111000011101111;
ROM[9521] <= 32'b11111111110000010000000100010011;
ROM[9522] <= 32'b00000000000000010010001110000011;
ROM[9523] <= 32'b00000000011100100010001000100011;
ROM[9524] <= 32'b00000000000000000000001110010011;
ROM[9525] <= 32'b00000000011100011010000000100011;
ROM[9526] <= 32'b00000000010000100010001110000011;
ROM[9527] <= 32'b00000000011100010010000000100011;
ROM[9528] <= 32'b00000000010000010000000100010011;
ROM[9529] <= 32'b00000000000000100010001110000011;
ROM[9530] <= 32'b11111111110000010000000100010011;
ROM[9531] <= 32'b00000000000000010010010000000011;
ROM[9532] <= 32'b00000000100000111010001110110011;
ROM[9533] <= 32'b01000000011100000000001110110011;
ROM[9534] <= 32'b00000000000100111000001110010011;
ROM[9535] <= 32'b00000000011100011010010000100011;
ROM[9536] <= 32'b00000000100000011010001110000011;
ROM[9537] <= 32'b01000000011100000000001110110011;
ROM[9538] <= 32'b00000000000100111000001110010011;
ROM[9539] <= 32'b00000000000000111000101001100011;
ROM[9540] <= 32'b00000000000000001001001110110111;
ROM[9541] <= 32'b01011000110000111000001110010011;
ROM[9542] <= 32'b00000000111000111000001110110011;
ROM[9543] <= 32'b00000000000000111000000011100111;
ROM[9544] <= 32'b00000000000000100010001110000011;
ROM[9545] <= 32'b00000000011100010010000000100011;
ROM[9546] <= 32'b00000000010000010000000100010011;
ROM[9547] <= 32'b00000000010000100010001110000011;
ROM[9548] <= 32'b11111111110000010000000100010011;
ROM[9549] <= 32'b00000000000000010010010000000011;
ROM[9550] <= 32'b01000000011101000000001110110011;
ROM[9551] <= 32'b00000000011100100010000000100011;
ROM[9552] <= 32'b00000000000000011010001110000011;
ROM[9553] <= 32'b00000000011100010010000000100011;
ROM[9554] <= 32'b00000000010000010000000100010011;
ROM[9555] <= 32'b00000000000100000000001110010011;
ROM[9556] <= 32'b11111111110000010000000100010011;
ROM[9557] <= 32'b00000000000000010010010000000011;
ROM[9558] <= 32'b00000000011101000000001110110011;
ROM[9559] <= 32'b00000000011100011010000000100011;
ROM[9560] <= 32'b00000000010000100010001110000011;
ROM[9561] <= 32'b00000000011100010010000000100011;
ROM[9562] <= 32'b00000000010000010000000100010011;
ROM[9563] <= 32'b00000000000000100010001110000011;
ROM[9564] <= 32'b11111111110000010000000100010011;
ROM[9565] <= 32'b00000000000000010010010000000011;
ROM[9566] <= 32'b00000000100000111010001110110011;
ROM[9567] <= 32'b01000000011100000000001110110011;
ROM[9568] <= 32'b00000000000100111000001110010011;
ROM[9569] <= 32'b00000000011100011010010000100011;
ROM[9570] <= 32'b11110111100111111111000011101111;
ROM[9571] <= 32'b00000000010000011010001110000011;
ROM[9572] <= 32'b00000000000000111000101001100011;
ROM[9573] <= 32'b00000000000000001001001110110111;
ROM[9574] <= 32'b01011010100000111000001110010011;
ROM[9575] <= 32'b00000000111000111000001110110011;
ROM[9576] <= 32'b00000000000000111000000011100111;
ROM[9577] <= 32'b00000001010000000000000011101111;
ROM[9578] <= 32'b00000000000000011010001110000011;
ROM[9579] <= 32'b01000000011100000000001110110011;
ROM[9580] <= 32'b00000000011100011010000000100011;
ROM[9581] <= 32'b00000000010000000000000011101111;
ROM[9582] <= 32'b00000000000000011010001110000011;
ROM[9583] <= 32'b00000000011100010010000000100011;
ROM[9584] <= 32'b00000000010000010000000100010011;
ROM[9585] <= 32'b00000001010000000000001110010011;
ROM[9586] <= 32'b01000000011100011000001110110011;
ROM[9587] <= 32'b00000000000000111010000010000011;
ROM[9588] <= 32'b11111111110000010000000100010011;
ROM[9589] <= 32'b00000000000000010010001110000011;
ROM[9590] <= 32'b00000000011100100010000000100011;
ROM[9591] <= 32'b00000000010000100000000100010011;
ROM[9592] <= 32'b00000001010000000000001110010011;
ROM[9593] <= 32'b01000000011100011000001110110011;
ROM[9594] <= 32'b00000000010000111010000110000011;
ROM[9595] <= 32'b00000000100000111010001000000011;
ROM[9596] <= 32'b00000000110000111010001010000011;
ROM[9597] <= 32'b00000001000000111010001100000011;
ROM[9598] <= 32'b00000000000000001000000011100111;
ROM[9599] <= 32'b00000000000000100010001110000011;
ROM[9600] <= 32'b00000000011100010010000000100011;
ROM[9601] <= 32'b00000000010000010000000100010011;
ROM[9602] <= 32'b00000000010000000000001110010011;
ROM[9603] <= 32'b00000000011100010010000000100011;
ROM[9604] <= 32'b00000000010000010000000100010011;
ROM[9605] <= 32'b00000000000000001001001110110111;
ROM[9606] <= 32'b01100110000000111000001110010011;
ROM[9607] <= 32'b00000000111000111000001110110011;
ROM[9608] <= 32'b00000000011100010010000000100011;
ROM[9609] <= 32'b00000000010000010000000100010011;
ROM[9610] <= 32'b00000000001100010010000000100011;
ROM[9611] <= 32'b00000000010000010000000100010011;
ROM[9612] <= 32'b00000000010000010010000000100011;
ROM[9613] <= 32'b00000000010000010000000100010011;
ROM[9614] <= 32'b00000000010100010010000000100011;
ROM[9615] <= 32'b00000000010000010000000100010011;
ROM[9616] <= 32'b00000000011000010010000000100011;
ROM[9617] <= 32'b00000000010000010000000100010011;
ROM[9618] <= 32'b00000001010000000000001110010011;
ROM[9619] <= 32'b00000000100000111000001110010011;
ROM[9620] <= 32'b01000000011100010000001110110011;
ROM[9621] <= 32'b00000000011100000000001000110011;
ROM[9622] <= 32'b00000000001000000000000110110011;
ROM[9623] <= 32'b10100111100111111111000011101111;
ROM[9624] <= 32'b11111111110000010000000100010011;
ROM[9625] <= 32'b00000000000000010010001110000011;
ROM[9626] <= 32'b00000000011100100010000000100011;
ROM[9627] <= 32'b00000000000000100010001110000011;
ROM[9628] <= 32'b00000000011100010010000000100011;
ROM[9629] <= 32'b00000000010000010000000100010011;
ROM[9630] <= 32'b00000100100001101010001110000011;
ROM[9631] <= 32'b11111111110000010000000100010011;
ROM[9632] <= 32'b00000000000000010010010000000011;
ROM[9633] <= 32'b00000000011101000000001110110011;
ROM[9634] <= 32'b00000000000000111000001100010011;
ROM[9635] <= 32'b00000000110100110000010000110011;
ROM[9636] <= 32'b00000000000001000010001110000011;
ROM[9637] <= 32'b00000000011100010010000000100011;
ROM[9638] <= 32'b00000000010000010000000100010011;
ROM[9639] <= 32'b00000001010000000000001110010011;
ROM[9640] <= 32'b01000000011100011000001110110011;
ROM[9641] <= 32'b00000000000000111010000010000011;
ROM[9642] <= 32'b11111111110000010000000100010011;
ROM[9643] <= 32'b00000000000000010010001110000011;
ROM[9644] <= 32'b00000000011100100010000000100011;
ROM[9645] <= 32'b00000000010000100000000100010011;
ROM[9646] <= 32'b00000001010000000000001110010011;
ROM[9647] <= 32'b01000000011100011000001110110011;
ROM[9648] <= 32'b00000000010000111010000110000011;
ROM[9649] <= 32'b00000000100000111010001000000011;
ROM[9650] <= 32'b00000000110000111010001010000011;
ROM[9651] <= 32'b00000001000000111010001100000011;
ROM[9652] <= 32'b00000000000000001000000011100111;
ROM[9653] <= 32'b00000000000000000010001110110111;
ROM[9654] <= 32'b00000000000000111000001110010011;
ROM[9655] <= 32'b00000100011101101010011000100011;
ROM[9656] <= 32'b00000000000000000100001110110111;
ROM[9657] <= 32'b00000000000000111000001110010011;
ROM[9658] <= 32'b00000100011101101010100000100011;
ROM[9659] <= 32'b00000101000001101010001110000011;
ROM[9660] <= 32'b00000000011100010010000000100011;
ROM[9661] <= 32'b00000000010000010000000100010011;
ROM[9662] <= 32'b00000000010000000000001110010011;
ROM[9663] <= 32'b00000000011100010010000000100011;
ROM[9664] <= 32'b00000000010000010000000100010011;
ROM[9665] <= 32'b00000000000000001001001110110111;
ROM[9666] <= 32'b01110101000000111000001110010011;
ROM[9667] <= 32'b00000000111000111000001110110011;
ROM[9668] <= 32'b00000000011100010010000000100011;
ROM[9669] <= 32'b00000000010000010000000100010011;
ROM[9670] <= 32'b00000000001100010010000000100011;
ROM[9671] <= 32'b00000000010000010000000100010011;
ROM[9672] <= 32'b00000000010000010010000000100011;
ROM[9673] <= 32'b00000000010000010000000100010011;
ROM[9674] <= 32'b00000000010100010010000000100011;
ROM[9675] <= 32'b00000000010000010000000100010011;
ROM[9676] <= 32'b00000000011000010010000000100011;
ROM[9677] <= 32'b00000000010000010000000100010011;
ROM[9678] <= 32'b00000001010000000000001110010011;
ROM[9679] <= 32'b00000000100000111000001110010011;
ROM[9680] <= 32'b01000000011100010000001110110011;
ROM[9681] <= 32'b00000000011100000000001000110011;
ROM[9682] <= 32'b00000000001000000000000110110011;
ROM[9683] <= 32'b10011000100111111111000011101111;
ROM[9684] <= 32'b11111111110000010000000100010011;
ROM[9685] <= 32'b00000000000000010010001110000011;
ROM[9686] <= 32'b00000100011101101010100000100011;
ROM[9687] <= 32'b00000000000000000001001110110111;
ROM[9688] <= 32'b10000000000000111000001110010011;
ROM[9689] <= 32'b00000100011101101010101000100011;
ROM[9690] <= 32'b00000000000000000100001110110111;
ROM[9691] <= 32'b00000000000000111000001110010011;
ROM[9692] <= 32'b00000100011101101010110000100011;
ROM[9693] <= 32'b00000000000000000000001110010011;
ROM[9694] <= 32'b00000100011101101010111000100011;
ROM[9695] <= 32'b00000100110001101010001110000011;
ROM[9696] <= 32'b00000110011101101010000000100011;
ROM[9697] <= 32'b00000000000000000000001110010011;
ROM[9698] <= 32'b00000110011101101010001000100011;
ROM[9699] <= 32'b00000000010000000000001110010011;
ROM[9700] <= 32'b00000110011101101010010000100011;
ROM[9701] <= 32'b00000110010001101010001110000011;
ROM[9702] <= 32'b00000000011100010010000000100011;
ROM[9703] <= 32'b00000000010000010000000100010011;
ROM[9704] <= 32'b00000110000001101010001110000011;
ROM[9705] <= 32'b11111111110000010000000100010011;
ROM[9706] <= 32'b00000000000000010010010000000011;
ROM[9707] <= 32'b00000000011101000000001110110011;
ROM[9708] <= 32'b00000000011100010010000000100011;
ROM[9709] <= 32'b00000000010000010000000100010011;
ROM[9710] <= 32'b00000101100001101010001110000011;
ROM[9711] <= 32'b00000000011100010010000000100011;
ROM[9712] <= 32'b00000000010000010000000100010011;
ROM[9713] <= 32'b00000101010001101010001110000011;
ROM[9714] <= 32'b11111111110000010000000100010011;
ROM[9715] <= 32'b00000000000000010010010000000011;
ROM[9716] <= 32'b01000000011101000000001110110011;
ROM[9717] <= 32'b00000000011101100010000000100011;
ROM[9718] <= 32'b11111111110000010000000100010011;
ROM[9719] <= 32'b00000000000000010010001110000011;
ROM[9720] <= 32'b00000000000000111000001100010011;
ROM[9721] <= 32'b00000000000001100010001110000011;
ROM[9722] <= 32'b00000000110100110000010000110011;
ROM[9723] <= 32'b00000000011101000010000000100011;
ROM[9724] <= 32'b00000110100001101010001110000011;
ROM[9725] <= 32'b00000000011100010010000000100011;
ROM[9726] <= 32'b00000000010000010000000100010011;
ROM[9727] <= 32'b00000110000001101010001110000011;
ROM[9728] <= 32'b11111111110000010000000100010011;
ROM[9729] <= 32'b00000000000000010010010000000011;
ROM[9730] <= 32'b00000000011101000000001110110011;
ROM[9731] <= 32'b00000000011100010010000000100011;
ROM[9732] <= 32'b00000000010000010000000100010011;
ROM[9733] <= 32'b00000000000000000000001110010011;
ROM[9734] <= 32'b00000000011101100010000000100011;
ROM[9735] <= 32'b11111111110000010000000100010011;
ROM[9736] <= 32'b00000000000000010010001110000011;
ROM[9737] <= 32'b00000000000000111000001100010011;
ROM[9738] <= 32'b00000000000001100010001110000011;
ROM[9739] <= 32'b00000000110100110000010000110011;
ROM[9740] <= 32'b00000000011101000010000000100011;
ROM[9741] <= 32'b00000000010000000000001110010011;
ROM[9742] <= 32'b01000000011100000000001110110011;
ROM[9743] <= 32'b00000110011101101010011000100011;
ROM[9744] <= 32'b00000000000000000000001110010011;
ROM[9745] <= 32'b00000000011100010010000000100011;
ROM[9746] <= 32'b00000000010000010000000100010011;
ROM[9747] <= 32'b00000001010000000000001110010011;
ROM[9748] <= 32'b01000000011100011000001110110011;
ROM[9749] <= 32'b00000000000000111010000010000011;
ROM[9750] <= 32'b11111111110000010000000100010011;
ROM[9751] <= 32'b00000000000000010010001110000011;
ROM[9752] <= 32'b00000000011100100010000000100011;
ROM[9753] <= 32'b00000000010000100000000100010011;
ROM[9754] <= 32'b00000001010000000000001110010011;
ROM[9755] <= 32'b01000000011100011000001110110011;
ROM[9756] <= 32'b00000000010000111010000110000011;
ROM[9757] <= 32'b00000000100000111010001000000011;
ROM[9758] <= 32'b00000000110000111010001010000011;
ROM[9759] <= 32'b00000001000000111010001100000011;
ROM[9760] <= 32'b00000000000000001000000011100111;
ROM[9761] <= 32'b00000000000000100010001110000011;
ROM[9762] <= 32'b00000000011100010010000000100011;
ROM[9763] <= 32'b00000000010000010000000100010011;
ROM[9764] <= 32'b00000000000000100010001110000011;
ROM[9765] <= 32'b11111111110000010000000100010011;
ROM[9766] <= 32'b00000000000000010010010000000011;
ROM[9767] <= 32'b00000000011101000000001110110011;
ROM[9768] <= 32'b00000000011100100010000000100011;
ROM[9769] <= 32'b00000000000000100010001110000011;
ROM[9770] <= 32'b00000000011100010010000000100011;
ROM[9771] <= 32'b00000000010000010000000100010011;
ROM[9772] <= 32'b00000000000000100010001110000011;
ROM[9773] <= 32'b11111111110000010000000100010011;
ROM[9774] <= 32'b00000000000000010010010000000011;
ROM[9775] <= 32'b00000000011101000000001110110011;
ROM[9776] <= 32'b00000000011100100010000000100011;
ROM[9777] <= 32'b00000000000000100010001110000011;
ROM[9778] <= 32'b00000000011100010010000000100011;
ROM[9779] <= 32'b00000000010000010000000100010011;
ROM[9780] <= 32'b00000101110001101010001110000011;
ROM[9781] <= 32'b11111111110000010000000100010011;
ROM[9782] <= 32'b00000000000000010010010000000011;
ROM[9783] <= 32'b00000000011101000000001110110011;
ROM[9784] <= 32'b00000000000000111000001100010011;
ROM[9785] <= 32'b00000000110100110000010000110011;
ROM[9786] <= 32'b00000000000001000010001110000011;
ROM[9787] <= 32'b00000000011100010010000000100011;
ROM[9788] <= 32'b00000000010000010000000100010011;
ROM[9789] <= 32'b00000001010000000000001110010011;
ROM[9790] <= 32'b01000000011100011000001110110011;
ROM[9791] <= 32'b00000000000000111010000010000011;
ROM[9792] <= 32'b11111111110000010000000100010011;
ROM[9793] <= 32'b00000000000000010010001110000011;
ROM[9794] <= 32'b00000000011100100010000000100011;
ROM[9795] <= 32'b00000000010000100000000100010011;
ROM[9796] <= 32'b00000001010000000000001110010011;
ROM[9797] <= 32'b01000000011100011000001110110011;
ROM[9798] <= 32'b00000000010000111010000110000011;
ROM[9799] <= 32'b00000000100000111010001000000011;
ROM[9800] <= 32'b00000000110000111010001010000011;
ROM[9801] <= 32'b00000001000000111010001100000011;
ROM[9802] <= 32'b00000000000000001000000011100111;
ROM[9803] <= 32'b00000000000000100010001110000011;
ROM[9804] <= 32'b00000000011100010010000000100011;
ROM[9805] <= 32'b00000000010000010000000100010011;
ROM[9806] <= 32'b00000000000000100010001110000011;
ROM[9807] <= 32'b11111111110000010000000100010011;
ROM[9808] <= 32'b00000000000000010010010000000011;
ROM[9809] <= 32'b00000000011101000000001110110011;
ROM[9810] <= 32'b00000000011100100010000000100011;
ROM[9811] <= 32'b00000000000000100010001110000011;
ROM[9812] <= 32'b00000000011100010010000000100011;
ROM[9813] <= 32'b00000000010000010000000100010011;
ROM[9814] <= 32'b00000000000000100010001110000011;
ROM[9815] <= 32'b11111111110000010000000100010011;
ROM[9816] <= 32'b00000000000000010010010000000011;
ROM[9817] <= 32'b00000000011101000000001110110011;
ROM[9818] <= 32'b00000000011100100010000000100011;
ROM[9819] <= 32'b00000000000000100010001110000011;
ROM[9820] <= 32'b00000000011100010010000000100011;
ROM[9821] <= 32'b00000000010000010000000100010011;
ROM[9822] <= 32'b00000101110001101010001110000011;
ROM[9823] <= 32'b11111111110000010000000100010011;
ROM[9824] <= 32'b00000000000000010010010000000011;
ROM[9825] <= 32'b00000000011101000000001110110011;
ROM[9826] <= 32'b00000000011100010010000000100011;
ROM[9827] <= 32'b00000000010000010000000100010011;
ROM[9828] <= 32'b00000000010000100010001110000011;
ROM[9829] <= 32'b00000000011101100010000000100011;
ROM[9830] <= 32'b11111111110000010000000100010011;
ROM[9831] <= 32'b00000000000000010010001110000011;
ROM[9832] <= 32'b00000000000000111000001100010011;
ROM[9833] <= 32'b00000000000001100010001110000011;
ROM[9834] <= 32'b00000000110100110000010000110011;
ROM[9835] <= 32'b00000000011101000010000000100011;
ROM[9836] <= 32'b00000000000000000000001110010011;
ROM[9837] <= 32'b00000000011100010010000000100011;
ROM[9838] <= 32'b00000000010000010000000100010011;
ROM[9839] <= 32'b00000001010000000000001110010011;
ROM[9840] <= 32'b01000000011100011000001110110011;
ROM[9841] <= 32'b00000000000000111010000010000011;
ROM[9842] <= 32'b11111111110000010000000100010011;
ROM[9843] <= 32'b00000000000000010010001110000011;
ROM[9844] <= 32'b00000000011100100010000000100011;
ROM[9845] <= 32'b00000000010000100000000100010011;
ROM[9846] <= 32'b00000001010000000000001110010011;
ROM[9847] <= 32'b01000000011100011000001110110011;
ROM[9848] <= 32'b00000000010000111010000110000011;
ROM[9849] <= 32'b00000000100000111010001000000011;
ROM[9850] <= 32'b00000000110000111010001010000011;
ROM[9851] <= 32'b00000001000000111010001100000011;
ROM[9852] <= 32'b00000000000000001000000011100111;
ROM[9853] <= 32'b00000000000000010010000000100011;
ROM[9854] <= 32'b00000000010000010000000100010011;
ROM[9855] <= 32'b00000000000000010010000000100011;
ROM[9856] <= 32'b00000000010000010000000100010011;
ROM[9857] <= 32'b00000000000000010010000000100011;
ROM[9858] <= 32'b00000000010000010000000100010011;
ROM[9859] <= 32'b00000000000000010010000000100011;
ROM[9860] <= 32'b00000000010000010000000100010011;
ROM[9861] <= 32'b00000000000000000000001110010011;
ROM[9862] <= 32'b00000000011100011010001000100011;
ROM[9863] <= 32'b00000101100001101010001110000011;
ROM[9864] <= 32'b00000000011100010010000000100011;
ROM[9865] <= 32'b00000000010000010000000100010011;
ROM[9866] <= 32'b00000101010001101010001110000011;
ROM[9867] <= 32'b11111111110000010000000100010011;
ROM[9868] <= 32'b00000000000000010010010000000011;
ROM[9869] <= 32'b01000000011101000000001110110011;
ROM[9870] <= 32'b00000000011100011010010000100011;
ROM[9871] <= 32'b00000110000001101010001110000011;
ROM[9872] <= 32'b00000000011100011010000000100011;
ROM[9873] <= 32'b00000110100001101010001110000011;
ROM[9874] <= 32'b00000000011100010010000000100011;
ROM[9875] <= 32'b00000000010000010000000100010011;
ROM[9876] <= 32'b00000000000000011010001110000011;
ROM[9877] <= 32'b11111111110000010000000100010011;
ROM[9878] <= 32'b00000000000000010010010000000011;
ROM[9879] <= 32'b00000000011101000000001110110011;
ROM[9880] <= 32'b00000000000000111000001100010011;
ROM[9881] <= 32'b00000000110100110000010000110011;
ROM[9882] <= 32'b00000000000001000010001110000011;
ROM[9883] <= 32'b00000000011100010010000000100011;
ROM[9884] <= 32'b00000000010000010000000100010011;
ROM[9885] <= 32'b00000000000000000000001110010011;
ROM[9886] <= 32'b11111111110000010000000100010011;
ROM[9887] <= 32'b00000000000000010010010000000011;
ROM[9888] <= 32'b00000000011101000010010010110011;
ROM[9889] <= 32'b00000000100000111010010100110011;
ROM[9890] <= 32'b00000000101001001000001110110011;
ROM[9891] <= 32'b00000000000100111000001110010011;
ROM[9892] <= 32'b00000000000100111111001110010011;
ROM[9893] <= 32'b00000000000000111000101001100011;
ROM[9894] <= 32'b00000000000000001010001110110111;
ROM[9895] <= 32'b10101010110000111000001110010011;
ROM[9896] <= 32'b00000000111000111000001110110011;
ROM[9897] <= 32'b00000000000000111000000011100111;
ROM[9898] <= 32'b00000100110000000000000011101111;
ROM[9899] <= 32'b00000000000000011010001110000011;
ROM[9900] <= 32'b00000000011100010010000000100011;
ROM[9901] <= 32'b00000000010000010000000100010011;
ROM[9902] <= 32'b00000001010000000000001110010011;
ROM[9903] <= 32'b01000000011100011000001110110011;
ROM[9904] <= 32'b00000000000000111010000010000011;
ROM[9905] <= 32'b11111111110000010000000100010011;
ROM[9906] <= 32'b00000000000000010010001110000011;
ROM[9907] <= 32'b00000000011100100010000000100011;
ROM[9908] <= 32'b00000000010000100000000100010011;
ROM[9909] <= 32'b00000001010000000000001110010011;
ROM[9910] <= 32'b01000000011100011000001110110011;
ROM[9911] <= 32'b00000000010000111010000110000011;
ROM[9912] <= 32'b00000000100000111010001000000011;
ROM[9913] <= 32'b00000000110000111010001010000011;
ROM[9914] <= 32'b00000001000000111010001100000011;
ROM[9915] <= 32'b00000000000000001000000011100111;
ROM[9916] <= 32'b00000000010000000000000011101111;
ROM[9917] <= 32'b00000000000000011010001110000011;
ROM[9918] <= 32'b00000000011100010010000000100011;
ROM[9919] <= 32'b00000000010000010000000100010011;
ROM[9920] <= 32'b00000000000000000000001110010011;
ROM[9921] <= 32'b11111111110000010000000100010011;
ROM[9922] <= 32'b00000000000000010010010000000011;
ROM[9923] <= 32'b00000000011101000010010010110011;
ROM[9924] <= 32'b00000000100000111010010100110011;
ROM[9925] <= 32'b00000000101001001000001110110011;
ROM[9926] <= 32'b00000000000100111000001110010011;
ROM[9927] <= 32'b00000000000100111111001110010011;
ROM[9928] <= 32'b01000000011100000000001110110011;
ROM[9929] <= 32'b00000000000100111000001110010011;
ROM[9930] <= 32'b01000000011100000000001110110011;
ROM[9931] <= 32'b00000000000100111000001110010011;
ROM[9932] <= 32'b00000000000000111000101001100011;
ROM[9933] <= 32'b00000000000000001010001110110111;
ROM[9934] <= 32'b11000011100000111000001110010011;
ROM[9935] <= 32'b00000000111000111000001110110011;
ROM[9936] <= 32'b00000000000000111000000011100111;
ROM[9937] <= 32'b00000110010001101010001110000011;
ROM[9938] <= 32'b00000000011100010010000000100011;
ROM[9939] <= 32'b00000000010000010000000100010011;
ROM[9940] <= 32'b00000000000000011010001110000011;
ROM[9941] <= 32'b11111111110000010000000100010011;
ROM[9942] <= 32'b00000000000000010010010000000011;
ROM[9943] <= 32'b00000000011101000000001110110011;
ROM[9944] <= 32'b00000000000000111000001100010011;
ROM[9945] <= 32'b00000000110100110000010000110011;
ROM[9946] <= 32'b00000000000001000010001110000011;
ROM[9947] <= 32'b00000000011100010010000000100011;
ROM[9948] <= 32'b00000000010000010000000100010011;
ROM[9949] <= 32'b00000000000100000000001110010011;
ROM[9950] <= 32'b11111111110000010000000100010011;
ROM[9951] <= 32'b00000000000000010010010000000011;
ROM[9952] <= 32'b01000000011101000000001110110011;
ROM[9953] <= 32'b00000000011100011010011000100011;
ROM[9954] <= 32'b00000000110000011010001110000011;
ROM[9955] <= 32'b00000000011100010010000000100011;
ROM[9956] <= 32'b00000000010000010000000100010011;
ROM[9957] <= 32'b00000000000000100010001110000011;
ROM[9958] <= 32'b11111111110000010000000100010011;
ROM[9959] <= 32'b00000000000000010010010000000011;
ROM[9960] <= 32'b00000000011101000010001110110011;
ROM[9961] <= 32'b01000000011100000000001110110011;
ROM[9962] <= 32'b00000000000100111000001110010011;
ROM[9963] <= 32'b00000000011100010010000000100011;
ROM[9964] <= 32'b00000000010000010000000100010011;
ROM[9965] <= 32'b00000000110000011010001110000011;
ROM[9966] <= 32'b00000000011100010010000000100011;
ROM[9967] <= 32'b00000000010000010000000100010011;
ROM[9968] <= 32'b00000000100000011010001110000011;
ROM[9969] <= 32'b11111111110000010000000100010011;
ROM[9970] <= 32'b00000000000000010010010000000011;
ROM[9971] <= 32'b00000000011101000010001110110011;
ROM[9972] <= 32'b11111111110000010000000100010011;
ROM[9973] <= 32'b00000000000000010010010000000011;
ROM[9974] <= 32'b00000000011101000111001110110011;
ROM[9975] <= 32'b00000000000000111000101001100011;
ROM[9976] <= 32'b00000000000000001010001110110111;
ROM[9977] <= 32'b10111111010000111000001110010011;
ROM[9978] <= 32'b00000000111000111000001110110011;
ROM[9979] <= 32'b00000000000000111000000011100111;
ROM[9980] <= 32'b00000001100000000000000011101111;
ROM[9981] <= 32'b00000000000000011010001110000011;
ROM[9982] <= 32'b00000000011100011010001000100011;
ROM[9983] <= 32'b00000000110000011010001110000011;
ROM[9984] <= 32'b00000000011100011010010000100011;
ROM[9985] <= 32'b00000000010000000000000011101111;
ROM[9986] <= 32'b00000110100001101010001110000011;
ROM[9987] <= 32'b00000000011100010010000000100011;
ROM[9988] <= 32'b00000000010000010000000100010011;
ROM[9989] <= 32'b00000000000000011010001110000011;
ROM[9990] <= 32'b11111111110000010000000100010011;
ROM[9991] <= 32'b00000000000000010010010000000011;
ROM[9992] <= 32'b00000000011101000000001110110011;
ROM[9993] <= 32'b00000000000000111000001100010011;
ROM[9994] <= 32'b00000000110100110000010000110011;
ROM[9995] <= 32'b00000000000001000010001110000011;
ROM[9996] <= 32'b00000000011100011010000000100011;
ROM[9997] <= 32'b11101100000111111111000011101111;
ROM[9998] <= 32'b00000000010000011010001110000011;
ROM[9999] <= 32'b00000000011100010010000000100011;
ROM[10000] <= 32'b00000000010000010000000100010011;
ROM[10001] <= 32'b00000001010000000000001110010011;
ROM[10002] <= 32'b01000000011100011000001110110011;
ROM[10003] <= 32'b00000000000000111010000010000011;
ROM[10004] <= 32'b11111111110000010000000100010011;
ROM[10005] <= 32'b00000000000000010010001110000011;
ROM[10006] <= 32'b00000000011100100010000000100011;
ROM[10007] <= 32'b00000000010000100000000100010011;
ROM[10008] <= 32'b00000001010000000000001110010011;
ROM[10009] <= 32'b01000000011100011000001110110011;
ROM[10010] <= 32'b00000000010000111010000110000011;
ROM[10011] <= 32'b00000000100000111010001000000011;
ROM[10012] <= 32'b00000000110000111010001010000011;
ROM[10013] <= 32'b00000001000000111010001100000011;
ROM[10014] <= 32'b00000000000000001000000011100111;
ROM[10015] <= 32'b00000000000000010010000000100011;
ROM[10016] <= 32'b00000000010000010000000100010011;
ROM[10017] <= 32'b00000000000000010010000000100011;
ROM[10018] <= 32'b00000000010000010000000100010011;
ROM[10019] <= 32'b00000000000000010010000000100011;
ROM[10020] <= 32'b00000000010000010000000100010011;
ROM[10021] <= 32'b00000110110001101010001110000011;
ROM[10022] <= 32'b00000000011100010010000000100011;
ROM[10023] <= 32'b00000000010000010000000100010011;
ROM[10024] <= 32'b00000000000000100010001110000011;
ROM[10025] <= 32'b11111111110000010000000100010011;
ROM[10026] <= 32'b00000000000000010010010000000011;
ROM[10027] <= 32'b00000000011101000000001110110011;
ROM[10028] <= 32'b00000000000000111000001100010011;
ROM[10029] <= 32'b00000000110100110000010000110011;
ROM[10030] <= 32'b00000000000001000010001110000011;
ROM[10031] <= 32'b00000000011100011010010000100011;
ROM[10032] <= 32'b00000000000000100010001110000011;
ROM[10033] <= 32'b00000000011100010010000000100011;
ROM[10034] <= 32'b00000000010000010000000100010011;
ROM[10035] <= 32'b00000000000100000000001110010011;
ROM[10036] <= 32'b11111111110000010000000100010011;
ROM[10037] <= 32'b00000000000000010010010000000011;
ROM[10038] <= 32'b00000000011101000000001110110011;
ROM[10039] <= 32'b00000000011100100010000000100011;
ROM[10040] <= 32'b00000000000000100010001110000011;
ROM[10041] <= 32'b00000000011100010010000000100011;
ROM[10042] <= 32'b00000000010000010000000100010011;
ROM[10043] <= 32'b00000000000000001010001110110111;
ROM[10044] <= 32'b11010011100000111000001110010011;
ROM[10045] <= 32'b00000000111000111000001110110011;
ROM[10046] <= 32'b00000000011100010010000000100011;
ROM[10047] <= 32'b00000000010000010000000100010011;
ROM[10048] <= 32'b00000000001100010010000000100011;
ROM[10049] <= 32'b00000000010000010000000100010011;
ROM[10050] <= 32'b00000000010000010010000000100011;
ROM[10051] <= 32'b00000000010000010000000100010011;
ROM[10052] <= 32'b00000000010100010010000000100011;
ROM[10053] <= 32'b00000000010000010000000100010011;
ROM[10054] <= 32'b00000000011000010010000000100011;
ROM[10055] <= 32'b00000000010000010000000100010011;
ROM[10056] <= 32'b00000001010000000000001110010011;
ROM[10057] <= 32'b00000000010000111000001110010011;
ROM[10058] <= 32'b01000000011100010000001110110011;
ROM[10059] <= 32'b00000000011100000000001000110011;
ROM[10060] <= 32'b00000000001000000000000110110011;
ROM[10061] <= 32'b01010000100000000000000011101111;
ROM[10062] <= 32'b11111111110000010000000100010011;
ROM[10063] <= 32'b00000000000000010010001110000011;
ROM[10064] <= 32'b00000000011100011010000000100011;
ROM[10065] <= 32'b00000000000000011010001110000011;
ROM[10066] <= 32'b00000000011100010010000000100011;
ROM[10067] <= 32'b00000000010000010000000100010011;
ROM[10068] <= 32'b00000000000000000000001110010011;
ROM[10069] <= 32'b11111111110000010000000100010011;
ROM[10070] <= 32'b00000000000000010010010000000011;
ROM[10071] <= 32'b00000000011101000010010010110011;
ROM[10072] <= 32'b00000000100000111010010100110011;
ROM[10073] <= 32'b00000000101001001000001110110011;
ROM[10074] <= 32'b00000000000100111000001110010011;
ROM[10075] <= 32'b00000000000100111111001110010011;
ROM[10076] <= 32'b00000000000000111000101001100011;
ROM[10077] <= 32'b00000000000000001010001110110111;
ROM[10078] <= 32'b11011000100000111000001110010011;
ROM[10079] <= 32'b00000000111000111000001110110011;
ROM[10080] <= 32'b00000000000000111000000011100111;
ROM[10081] <= 32'b00001001100000000000000011101111;
ROM[10082] <= 32'b00000110010001101010001110000011;
ROM[10083] <= 32'b00000000011100010010000000100011;
ROM[10084] <= 32'b00000000010000010000000100010011;
ROM[10085] <= 32'b00000000000000100010001110000011;
ROM[10086] <= 32'b11111111110000010000000100010011;
ROM[10087] <= 32'b00000000000000010010010000000011;
ROM[10088] <= 32'b00000000011101000000001110110011;
ROM[10089] <= 32'b00000000011100010010000000100011;
ROM[10090] <= 32'b00000000010000010000000100010011;
ROM[10091] <= 32'b00000000100000011010001110000011;
ROM[10092] <= 32'b00000000011101100010000000100011;
ROM[10093] <= 32'b11111111110000010000000100010011;
ROM[10094] <= 32'b00000000000000010010001110000011;
ROM[10095] <= 32'b00000000000000111000001100010011;
ROM[10096] <= 32'b00000000000001100010001110000011;
ROM[10097] <= 32'b00000000110100110000010000110011;
ROM[10098] <= 32'b00000000011101000010000000100011;
ROM[10099] <= 32'b00000110100001101010001110000011;
ROM[10100] <= 32'b00000000011100010010000000100011;
ROM[10101] <= 32'b00000000010000010000000100010011;
ROM[10102] <= 32'b00000000000000100010001110000011;
ROM[10103] <= 32'b11111111110000010000000100010011;
ROM[10104] <= 32'b00000000000000010010010000000011;
ROM[10105] <= 32'b00000000011101000000001110110011;
ROM[10106] <= 32'b00000000011100010010000000100011;
ROM[10107] <= 32'b00000000010000010000000100010011;
ROM[10108] <= 32'b00000110000001101010001110000011;
ROM[10109] <= 32'b00000000011101100010000000100011;
ROM[10110] <= 32'b11111111110000010000000100010011;
ROM[10111] <= 32'b00000000000000010010001110000011;
ROM[10112] <= 32'b00000000000000111000001100010011;
ROM[10113] <= 32'b00000000000001100010001110000011;
ROM[10114] <= 32'b00000000110100110000010000110011;
ROM[10115] <= 32'b00000000011101000010000000100011;
ROM[10116] <= 32'b00000000000000100010001110000011;
ROM[10117] <= 32'b00000110011101101010000000100011;
ROM[10118] <= 32'b00100000000000000000000011101111;
ROM[10119] <= 32'b00000000000000011010001110000011;
ROM[10120] <= 32'b00000000011100010010000000100011;
ROM[10121] <= 32'b00000000010000010000000100010011;
ROM[10122] <= 32'b00000110010001101010001110000011;
ROM[10123] <= 32'b00000000011100010010000000100011;
ROM[10124] <= 32'b00000000010000010000000100010011;
ROM[10125] <= 32'b00000000000000011010001110000011;
ROM[10126] <= 32'b11111111110000010000000100010011;
ROM[10127] <= 32'b00000000000000010010010000000011;
ROM[10128] <= 32'b00000000011101000000001110110011;
ROM[10129] <= 32'b00000000000000111000001100010011;
ROM[10130] <= 32'b00000000110100110000010000110011;
ROM[10131] <= 32'b00000000000001000010001110000011;
ROM[10132] <= 32'b11111111110000010000000100010011;
ROM[10133] <= 32'b00000000000000010010010000000011;
ROM[10134] <= 32'b01000000011101000000001110110011;
ROM[10135] <= 32'b00000000011100010010000000100011;
ROM[10136] <= 32'b00000000010000010000000100010011;
ROM[10137] <= 32'b00000000000000100010001110000011;
ROM[10138] <= 32'b11111111110000010000000100010011;
ROM[10139] <= 32'b00000000000000010010010000000011;
ROM[10140] <= 32'b00000000011101000010010010110011;
ROM[10141] <= 32'b00000000100000111010010100110011;
ROM[10142] <= 32'b00000000101001001000001110110011;
ROM[10143] <= 32'b00000000000100111000001110010011;
ROM[10144] <= 32'b00000000000100111111001110010011;
ROM[10145] <= 32'b00000000000000111000101001100011;
ROM[10146] <= 32'b00000000000000001010001110110111;
ROM[10147] <= 32'b11101001110000111000001110010011;
ROM[10148] <= 32'b00000000111000111000001110110011;
ROM[10149] <= 32'b00000000000000111000000011100111;
ROM[10150] <= 32'b00001001000000000000000011101111;
ROM[10151] <= 32'b00000110010001101010001110000011;
ROM[10152] <= 32'b00000000011100010010000000100011;
ROM[10153] <= 32'b00000000010000010000000100010011;
ROM[10154] <= 32'b00000000000000011010001110000011;
ROM[10155] <= 32'b11111111110000010000000100010011;
ROM[10156] <= 32'b00000000000000010010010000000011;
ROM[10157] <= 32'b00000000011101000000001110110011;
ROM[10158] <= 32'b00000000011100010010000000100011;
ROM[10159] <= 32'b00000000010000010000000100010011;
ROM[10160] <= 32'b00000110010001101010001110000011;
ROM[10161] <= 32'b00000000011100010010000000100011;
ROM[10162] <= 32'b00000000010000010000000100010011;
ROM[10163] <= 32'b00000000000000011010001110000011;
ROM[10164] <= 32'b11111111110000010000000100010011;
ROM[10165] <= 32'b00000000000000010010010000000011;
ROM[10166] <= 32'b00000000011101000000001110110011;
ROM[10167] <= 32'b00000000000000111000001100010011;
ROM[10168] <= 32'b00000000110100110000010000110011;
ROM[10169] <= 32'b00000000000001000010001110000011;
ROM[10170] <= 32'b00000000011100010010000000100011;
ROM[10171] <= 32'b00000000010000010000000100010011;
ROM[10172] <= 32'b00000000100000011010001110000011;
ROM[10173] <= 32'b11111111110000010000000100010011;
ROM[10174] <= 32'b00000000000000010010010000000011;
ROM[10175] <= 32'b00000000011101000000001110110011;
ROM[10176] <= 32'b00000000011101100010000000100011;
ROM[10177] <= 32'b11111111110000010000000100010011;
ROM[10178] <= 32'b00000000000000010010001110000011;
ROM[10179] <= 32'b00000000000000111000001100010011;
ROM[10180] <= 32'b00000000000001100010001110000011;
ROM[10181] <= 32'b00000000110100110000010000110011;
ROM[10182] <= 32'b00000000011101000010000000100011;
ROM[10183] <= 32'b00000000000000011010001110000011;
ROM[10184] <= 32'b00000000011100100010000000100011;
ROM[10185] <= 32'b00001111010000000000000011101111;
ROM[10186] <= 32'b00000110010001101010001110000011;
ROM[10187] <= 32'b00000000011100010010000000100011;
ROM[10188] <= 32'b00000000010000010000000100010011;
ROM[10189] <= 32'b00000000000000100010001110000011;
ROM[10190] <= 32'b11111111110000010000000100010011;
ROM[10191] <= 32'b00000000000000010010010000000011;
ROM[10192] <= 32'b00000000011101000000001110110011;
ROM[10193] <= 32'b00000000011100010010000000100011;
ROM[10194] <= 32'b00000000010000010000000100010011;
ROM[10195] <= 32'b00000000100000011010001110000011;
ROM[10196] <= 32'b00000000011101100010000000100011;
ROM[10197] <= 32'b11111111110000010000000100010011;
ROM[10198] <= 32'b00000000000000010010001110000011;
ROM[10199] <= 32'b00000000000000111000001100010011;
ROM[10200] <= 32'b00000000000001100010001110000011;
ROM[10201] <= 32'b00000000110100110000010000110011;
ROM[10202] <= 32'b00000000011101000010000000100011;
ROM[10203] <= 32'b00000110100001101010001110000011;
ROM[10204] <= 32'b00000000011100010010000000100011;
ROM[10205] <= 32'b00000000010000010000000100010011;
ROM[10206] <= 32'b00000000000000100010001110000011;
ROM[10207] <= 32'b11111111110000010000000100010011;
ROM[10208] <= 32'b00000000000000010010010000000011;
ROM[10209] <= 32'b00000000011101000000001110110011;
ROM[10210] <= 32'b00000000011100010010000000100011;
ROM[10211] <= 32'b00000000010000010000000100010011;
ROM[10212] <= 32'b00000110100001101010001110000011;
ROM[10213] <= 32'b00000000011100010010000000100011;
ROM[10214] <= 32'b00000000010000010000000100010011;
ROM[10215] <= 32'b00000000000000011010001110000011;
ROM[10216] <= 32'b11111111110000010000000100010011;
ROM[10217] <= 32'b00000000000000010010010000000011;
ROM[10218] <= 32'b00000000011101000000001110110011;
ROM[10219] <= 32'b00000000000000111000001100010011;
ROM[10220] <= 32'b00000000110100110000010000110011;
ROM[10221] <= 32'b00000000000001000010001110000011;
ROM[10222] <= 32'b00000000011101100010000000100011;
ROM[10223] <= 32'b11111111110000010000000100010011;
ROM[10224] <= 32'b00000000000000010010001110000011;
ROM[10225] <= 32'b00000000000000111000001100010011;
ROM[10226] <= 32'b00000000000001100010001110000011;
ROM[10227] <= 32'b00000000110100110000010000110011;
ROM[10228] <= 32'b00000000011101000010000000100011;
ROM[10229] <= 32'b00000110100001101010001110000011;
ROM[10230] <= 32'b00000000011100010010000000100011;
ROM[10231] <= 32'b00000000010000010000000100010011;
ROM[10232] <= 32'b00000000000000011010001110000011;
ROM[10233] <= 32'b11111111110000010000000100010011;
ROM[10234] <= 32'b00000000000000010010010000000011;
ROM[10235] <= 32'b00000000011101000000001110110011;
ROM[10236] <= 32'b00000000011100010010000000100011;
ROM[10237] <= 32'b00000000010000010000000100010011;
ROM[10238] <= 32'b00000000000000100010001110000011;
ROM[10239] <= 32'b00000000011101100010000000100011;
ROM[10240] <= 32'b11111111110000010000000100010011;
ROM[10241] <= 32'b00000000000000010010001110000011;
ROM[10242] <= 32'b00000000000000111000001100010011;
ROM[10243] <= 32'b00000000000001100010001110000011;
ROM[10244] <= 32'b00000000110100110000010000110011;
ROM[10245] <= 32'b00000000011101000010000000100011;
ROM[10246] <= 32'b00000000000000100010001110000011;
ROM[10247] <= 32'b00000000011100010010000000100011;
ROM[10248] <= 32'b00000000010000010000000100010011;
ROM[10249] <= 32'b00000110010001101010001110000011;
ROM[10250] <= 32'b00000000011100010010000000100011;
ROM[10251] <= 32'b00000000010000010000000100010011;
ROM[10252] <= 32'b00000000000000100010001110000011;
ROM[10253] <= 32'b11111111110000010000000100010011;
ROM[10254] <= 32'b00000000000000010010010000000011;
ROM[10255] <= 32'b00000000011101000000001110110011;
ROM[10256] <= 32'b00000000000000111000001100010011;
ROM[10257] <= 32'b00000000110100110000010000110011;
ROM[10258] <= 32'b00000000000001000010001110000011;
ROM[10259] <= 32'b11111111110000010000000100010011;
ROM[10260] <= 32'b00000000000000010010010000000011;
ROM[10261] <= 32'b01000000011101000000001110110011;
ROM[10262] <= 32'b00000000011100010010000000100011;
ROM[10263] <= 32'b00000000010000010000000100010011;
ROM[10264] <= 32'b00000110100001101010001110000011;
ROM[10265] <= 32'b00000000011100010010000000100011;
ROM[10266] <= 32'b00000000010000010000000100010011;
ROM[10267] <= 32'b00000000000000100010001110000011;
ROM[10268] <= 32'b11111111110000010000000100010011;
ROM[10269] <= 32'b00000000000000010010010000000011;
ROM[10270] <= 32'b00000000011101000000001110110011;
ROM[10271] <= 32'b00000000000000111000001100010011;
ROM[10272] <= 32'b00000000110100110000010000110011;
ROM[10273] <= 32'b00000000000001000010001110000011;
ROM[10274] <= 32'b11111111110000010000000100010011;
ROM[10275] <= 32'b00000000000000010010010000000011;
ROM[10276] <= 32'b00000000011101000010010010110011;
ROM[10277] <= 32'b00000000100000111010010100110011;
ROM[10278] <= 32'b00000000101001001000001110110011;
ROM[10279] <= 32'b00000000000100111000001110010011;
ROM[10280] <= 32'b00000000000100111111001110010011;
ROM[10281] <= 32'b00000000000000111000101001100011;
ROM[10282] <= 32'b00000000000000001010001110110111;
ROM[10283] <= 32'b00001011110000111000001110010011;
ROM[10284] <= 32'b00000000111000111000001110110011;
ROM[10285] <= 32'b00000000000000111000000011100111;
ROM[10286] <= 32'b00010100000000000000000011101111;
ROM[10287] <= 32'b00000110100001101010001110000011;
ROM[10288] <= 32'b00000000011100010010000000100011;
ROM[10289] <= 32'b00000000010000010000000100010011;
ROM[10290] <= 32'b00000000000000100010001110000011;
ROM[10291] <= 32'b11111111110000010000000100010011;
ROM[10292] <= 32'b00000000000000010010010000000011;
ROM[10293] <= 32'b00000000011101000000001110110011;
ROM[10294] <= 32'b00000000000000111000001100010011;
ROM[10295] <= 32'b00000000110100110000010000110011;
ROM[10296] <= 32'b00000000000001000010001110000011;
ROM[10297] <= 32'b00000000011100011010001000100011;
ROM[10298] <= 32'b00000110010001101010001110000011;
ROM[10299] <= 32'b00000000011100010010000000100011;
ROM[10300] <= 32'b00000000010000010000000100010011;
ROM[10301] <= 32'b00000000000000100010001110000011;
ROM[10302] <= 32'b11111111110000010000000100010011;
ROM[10303] <= 32'b00000000000000010010010000000011;
ROM[10304] <= 32'b00000000011101000000001110110011;
ROM[10305] <= 32'b00000000011100010010000000100011;
ROM[10306] <= 32'b00000000010000010000000100010011;
ROM[10307] <= 32'b00000110010001101010001110000011;
ROM[10308] <= 32'b00000000011100010010000000100011;
ROM[10309] <= 32'b00000000010000010000000100010011;
ROM[10310] <= 32'b00000000000000100010001110000011;
ROM[10311] <= 32'b11111111110000010000000100010011;
ROM[10312] <= 32'b00000000000000010010010000000011;
ROM[10313] <= 32'b00000000011101000000001110110011;
ROM[10314] <= 32'b00000000000000111000001100010011;
ROM[10315] <= 32'b00000000110100110000010000110011;
ROM[10316] <= 32'b00000000000001000010001110000011;
ROM[10317] <= 32'b00000000011100010010000000100011;
ROM[10318] <= 32'b00000000010000010000000100010011;
ROM[10319] <= 32'b00000110010001101010001110000011;
ROM[10320] <= 32'b00000000011100010010000000100011;
ROM[10321] <= 32'b00000000010000010000000100010011;
ROM[10322] <= 32'b00000000010000011010001110000011;
ROM[10323] <= 32'b11111111110000010000000100010011;
ROM[10324] <= 32'b00000000000000010010010000000011;
ROM[10325] <= 32'b00000000011101000000001110110011;
ROM[10326] <= 32'b00000000000000111000001100010011;
ROM[10327] <= 32'b00000000110100110000010000110011;
ROM[10328] <= 32'b00000000000001000010001110000011;
ROM[10329] <= 32'b11111111110000010000000100010011;
ROM[10330] <= 32'b00000000000000010010010000000011;
ROM[10331] <= 32'b00000000011101000000001110110011;
ROM[10332] <= 32'b00000000011101100010000000100011;
ROM[10333] <= 32'b11111111110000010000000100010011;
ROM[10334] <= 32'b00000000000000010010001110000011;
ROM[10335] <= 32'b00000000000000111000001100010011;
ROM[10336] <= 32'b00000000000001100010001110000011;
ROM[10337] <= 32'b00000000110100110000010000110011;
ROM[10338] <= 32'b00000000011101000010000000100011;
ROM[10339] <= 32'b00000110100001101010001110000011;
ROM[10340] <= 32'b00000000011100010010000000100011;
ROM[10341] <= 32'b00000000010000010000000100010011;
ROM[10342] <= 32'b00000000000000100010001110000011;
ROM[10343] <= 32'b11111111110000010000000100010011;
ROM[10344] <= 32'b00000000000000010010010000000011;
ROM[10345] <= 32'b00000000011101000000001110110011;
ROM[10346] <= 32'b00000000011100010010000000100011;
ROM[10347] <= 32'b00000000010000010000000100010011;
ROM[10348] <= 32'b00000110100001101010001110000011;
ROM[10349] <= 32'b00000000011100010010000000100011;
ROM[10350] <= 32'b00000000010000010000000100010011;
ROM[10351] <= 32'b00000000010000011010001110000011;
ROM[10352] <= 32'b11111111110000010000000100010011;
ROM[10353] <= 32'b00000000000000010010010000000011;
ROM[10354] <= 32'b00000000011101000000001110110011;
ROM[10355] <= 32'b00000000000000111000001100010011;
ROM[10356] <= 32'b00000000110100110000010000110011;
ROM[10357] <= 32'b00000000000001000010001110000011;
ROM[10358] <= 32'b00000000011101100010000000100011;
ROM[10359] <= 32'b11111111110000010000000100010011;
ROM[10360] <= 32'b00000000000000010010001110000011;
ROM[10361] <= 32'b00000000000000111000001100010011;
ROM[10362] <= 32'b00000000000001100010001110000011;
ROM[10363] <= 32'b00000000110100110000010000110011;
ROM[10364] <= 32'b00000000011101000010000000100011;
ROM[10365] <= 32'b00000000010000000000000011101111;
ROM[10366] <= 32'b00000000000000000000001110010011;
ROM[10367] <= 32'b00000000011100010010000000100011;
ROM[10368] <= 32'b00000000010000010000000100010011;
ROM[10369] <= 32'b00000001010000000000001110010011;
ROM[10370] <= 32'b01000000011100011000001110110011;
ROM[10371] <= 32'b00000000000000111010000010000011;
ROM[10372] <= 32'b11111111110000010000000100010011;
ROM[10373] <= 32'b00000000000000010010001110000011;
ROM[10374] <= 32'b00000000011100100010000000100011;
ROM[10375] <= 32'b00000000010000100000000100010011;
ROM[10376] <= 32'b00000001010000000000001110010011;
ROM[10377] <= 32'b01000000011100011000001110110011;
ROM[10378] <= 32'b00000000010000111010000110000011;
ROM[10379] <= 32'b00000000100000111010001000000011;
ROM[10380] <= 32'b00000000110000111010001010000011;
ROM[10381] <= 32'b00000001000000111010001100000011;
ROM[10382] <= 32'b00000000000000001000000011100111;
ROM[10383] <= 32'b00000000000000010010000000100011;
ROM[10384] <= 32'b00000000010000010000000100010011;
ROM[10385] <= 32'b00000110000001101010001110000011;
ROM[10386] <= 32'b00000000011100010010000000100011;
ROM[10387] <= 32'b00000000010000010000000100010011;
ROM[10388] <= 32'b00000000000000100010001110000011;
ROM[10389] <= 32'b11111111110000010000000100010011;
ROM[10390] <= 32'b00000000000000010010010000000011;
ROM[10391] <= 32'b00000000011101000010001110110011;
ROM[10392] <= 32'b00000000000000111000101001100011;
ROM[10393] <= 32'b00000000000000001010001110110111;
ROM[10394] <= 32'b00100111100000111000001110010011;
ROM[10395] <= 32'b00000000111000111000001110110011;
ROM[10396] <= 32'b00000000000000111000000011100111;
ROM[10397] <= 32'b00000100110000000000000011101111;
ROM[10398] <= 32'b00000000000000000000001110010011;
ROM[10399] <= 32'b00000000011100010010000000100011;
ROM[10400] <= 32'b00000000010000010000000100010011;
ROM[10401] <= 32'b00000001010000000000001110010011;
ROM[10402] <= 32'b01000000011100011000001110110011;
ROM[10403] <= 32'b00000000000000111010000010000011;
ROM[10404] <= 32'b11111111110000010000000100010011;
ROM[10405] <= 32'b00000000000000010010001110000011;
ROM[10406] <= 32'b00000000011100100010000000100011;
ROM[10407] <= 32'b00000000010000100000000100010011;
ROM[10408] <= 32'b00000001010000000000001110010011;
ROM[10409] <= 32'b01000000011100011000001110110011;
ROM[10410] <= 32'b00000000010000111010000110000011;
ROM[10411] <= 32'b00000000100000111010001000000011;
ROM[10412] <= 32'b00000000110000111010001010000011;
ROM[10413] <= 32'b00000001000000111010001100000011;
ROM[10414] <= 32'b00000000000000001000000011100111;
ROM[10415] <= 32'b00000000010000000000000011101111;
ROM[10416] <= 32'b00000110000001101010001110000011;
ROM[10417] <= 32'b00000000011100011010000000100011;
ROM[10418] <= 32'b00000110100001101010001110000011;
ROM[10419] <= 32'b00000000011100010010000000100011;
ROM[10420] <= 32'b00000000010000010000000100010011;
ROM[10421] <= 32'b00000000000000011010001110000011;
ROM[10422] <= 32'b11111111110000010000000100010011;
ROM[10423] <= 32'b00000000000000010010010000000011;
ROM[10424] <= 32'b00000000011101000000001110110011;
ROM[10425] <= 32'b00000000000000111000001100010011;
ROM[10426] <= 32'b00000000110100110000010000110011;
ROM[10427] <= 32'b00000000000001000010001110000011;
ROM[10428] <= 32'b00000000011100010010000000100011;
ROM[10429] <= 32'b00000000010000010000000100010011;
ROM[10430] <= 32'b00000000000000000000001110010011;
ROM[10431] <= 32'b11111111110000010000000100010011;
ROM[10432] <= 32'b00000000000000010010010000000011;
ROM[10433] <= 32'b00000000011101000010010010110011;
ROM[10434] <= 32'b00000000100000111010010100110011;
ROM[10435] <= 32'b00000000101001001000001110110011;
ROM[10436] <= 32'b00000000000100111000001110010011;
ROM[10437] <= 32'b00000000000100111111001110010011;
ROM[10438] <= 32'b01000000011100000000001110110011;
ROM[10439] <= 32'b00000000000100111000001110010011;
ROM[10440] <= 32'b00000000011100010010000000100011;
ROM[10441] <= 32'b00000000010000010000000100010011;
ROM[10442] <= 32'b00000110100001101010001110000011;
ROM[10443] <= 32'b00000000011100010010000000100011;
ROM[10444] <= 32'b00000000010000010000000100010011;
ROM[10445] <= 32'b00000000000000011010001110000011;
ROM[10446] <= 32'b11111111110000010000000100010011;
ROM[10447] <= 32'b00000000000000010010010000000011;
ROM[10448] <= 32'b00000000011101000000001110110011;
ROM[10449] <= 32'b00000000000000111000001100010011;
ROM[10450] <= 32'b00000000110100110000010000110011;
ROM[10451] <= 32'b00000000000001000010001110000011;
ROM[10452] <= 32'b00000000011100010010000000100011;
ROM[10453] <= 32'b00000000010000010000000100010011;
ROM[10454] <= 32'b00000000000000100010001110000011;
ROM[10455] <= 32'b11111111110000010000000100010011;
ROM[10456] <= 32'b00000000000000010010010000000011;
ROM[10457] <= 32'b00000000100000111010001110110011;
ROM[10458] <= 32'b11111111110000010000000100010011;
ROM[10459] <= 32'b00000000000000010010010000000011;
ROM[10460] <= 32'b00000000011101000111001110110011;
ROM[10461] <= 32'b01000000011100000000001110110011;
ROM[10462] <= 32'b00000000000100111000001110010011;
ROM[10463] <= 32'b00000000000000111000101001100011;
ROM[10464] <= 32'b00000000000000001010001110110111;
ROM[10465] <= 32'b00111100000000111000001110010011;
ROM[10466] <= 32'b00000000111000111000001110110011;
ROM[10467] <= 32'b00000000000000111000000011100111;
ROM[10468] <= 32'b00000110100001101010001110000011;
ROM[10469] <= 32'b00000000011100010010000000100011;
ROM[10470] <= 32'b00000000010000010000000100010011;
ROM[10471] <= 32'b00000000000000011010001110000011;
ROM[10472] <= 32'b11111111110000010000000100010011;
ROM[10473] <= 32'b00000000000000010010010000000011;
ROM[10474] <= 32'b00000000011101000000001110110011;
ROM[10475] <= 32'b00000000000000111000001100010011;
ROM[10476] <= 32'b00000000110100110000010000110011;
ROM[10477] <= 32'b00000000000001000010001110000011;
ROM[10478] <= 32'b00000000011100011010000000100011;
ROM[10479] <= 32'b11110000110111111111000011101111;
ROM[10480] <= 32'b00000000000000011010001110000011;
ROM[10481] <= 32'b00000000011100010010000000100011;
ROM[10482] <= 32'b00000000010000010000000100010011;
ROM[10483] <= 32'b00000001010000000000001110010011;
ROM[10484] <= 32'b01000000011100011000001110110011;
ROM[10485] <= 32'b00000000000000111010000010000011;
ROM[10486] <= 32'b11111111110000010000000100010011;
ROM[10487] <= 32'b00000000000000010010001110000011;
ROM[10488] <= 32'b00000000011100100010000000100011;
ROM[10489] <= 32'b00000000010000100000000100010011;
ROM[10490] <= 32'b00000001010000000000001110010011;
ROM[10491] <= 32'b01000000011100011000001110110011;
ROM[10492] <= 32'b00000000010000111010000110000011;
ROM[10493] <= 32'b00000000100000111010001000000011;
ROM[10494] <= 32'b00000000110000111010001010000011;
ROM[10495] <= 32'b00000001000000111010001100000011;
ROM[10496] <= 32'b00000000000000001000000011100111;
ROM[10497] <= 32'b00000000000000010010000000100011;
ROM[10498] <= 32'b00000000010000010000000100010011;
ROM[10499] <= 32'b00000000000000010010000000100011;
ROM[10500] <= 32'b00000000010000010000000100010011;
ROM[10501] <= 32'b00000000000000010010000000100011;
ROM[10502] <= 32'b00000000010000010000000100010011;
ROM[10503] <= 32'b00000000000000100010001110000011;
ROM[10504] <= 32'b00000000011100010010000000100011;
ROM[10505] <= 32'b00000000010000010000000100010011;
ROM[10506] <= 32'b00000000000000001010001110110111;
ROM[10507] <= 32'b01000111010000111000001110010011;
ROM[10508] <= 32'b00000000111000111000001110110011;
ROM[10509] <= 32'b00000000011100010010000000100011;
ROM[10510] <= 32'b00000000010000010000000100010011;
ROM[10511] <= 32'b00000000001100010010000000100011;
ROM[10512] <= 32'b00000000010000010000000100010011;
ROM[10513] <= 32'b00000000010000010010000000100011;
ROM[10514] <= 32'b00000000010000010000000100010011;
ROM[10515] <= 32'b00000000010100010010000000100011;
ROM[10516] <= 32'b00000000010000010000000100010011;
ROM[10517] <= 32'b00000000011000010010000000100011;
ROM[10518] <= 32'b00000000010000010000000100010011;
ROM[10519] <= 32'b00000001010000000000001110010011;
ROM[10520] <= 32'b00000000010000111000001110010011;
ROM[10521] <= 32'b01000000011100010000001110110011;
ROM[10522] <= 32'b00000000011100000000001000110011;
ROM[10523] <= 32'b00000000001000000000000110110011;
ROM[10524] <= 32'b11011000010011111111000011101111;
ROM[10525] <= 32'b11111111110000010000000100010011;
ROM[10526] <= 32'b00000000000000010010001110000011;
ROM[10527] <= 32'b00000000011100011010000000100011;
ROM[10528] <= 32'b00000000000000011010001110000011;
ROM[10529] <= 32'b00000000011100010010000000100011;
ROM[10530] <= 32'b00000000010000010000000100010011;
ROM[10531] <= 32'b00000000010000000000001110010011;
ROM[10532] <= 32'b11111111110000010000000100010011;
ROM[10533] <= 32'b00000000000000010010010000000011;
ROM[10534] <= 32'b00000000011101000000001110110011;
ROM[10535] <= 32'b00000000011100011010010000100011;
ROM[10536] <= 32'b00000000100000011010001110000011;
ROM[10537] <= 32'b00000110011101101010100000100011;
ROM[10538] <= 32'b00000000000000011010001110000011;
ROM[10539] <= 32'b00000000011100010010000000100011;
ROM[10540] <= 32'b00000000010000010000000100010011;
ROM[10541] <= 32'b00000000000000000000001110010011;
ROM[10542] <= 32'b11111111110000010000000100010011;
ROM[10543] <= 32'b00000000000000010010010000000011;
ROM[10544] <= 32'b00000000011101000010010010110011;
ROM[10545] <= 32'b00000000100000111010010100110011;
ROM[10546] <= 32'b00000000101001001000001110110011;
ROM[10547] <= 32'b00000000000100111000001110010011;
ROM[10548] <= 32'b00000000000100111111001110010011;
ROM[10549] <= 32'b01000000011100000000001110110011;
ROM[10550] <= 32'b00000000000100111000001110010011;
ROM[10551] <= 32'b00000000000000111000101001100011;
ROM[10552] <= 32'b00000000000000001010001110110111;
ROM[10553] <= 32'b01001111010000111000001110010011;
ROM[10554] <= 32'b00000000111000111000001110110011;
ROM[10555] <= 32'b00000000000000111000000011100111;
ROM[10556] <= 32'b00110000110000000000000011101111;
ROM[10557] <= 32'b00000110010001101010001110000011;
ROM[10558] <= 32'b00000000011100010010000000100011;
ROM[10559] <= 32'b00000000010000010000000100010011;
ROM[10560] <= 32'b00000000000000011010001110000011;
ROM[10561] <= 32'b11111111110000010000000100010011;
ROM[10562] <= 32'b00000000000000010010010000000011;
ROM[10563] <= 32'b00000000011101000000001110110011;
ROM[10564] <= 32'b00000000000000111000001100010011;
ROM[10565] <= 32'b00000000110100110000010000110011;
ROM[10566] <= 32'b00000000000001000010001110000011;
ROM[10567] <= 32'b00000000011100010010000000100011;
ROM[10568] <= 32'b00000000010000010000000100010011;
ROM[10569] <= 32'b00000000000000100010001110000011;
ROM[10570] <= 32'b00000000011100010010000000100011;
ROM[10571] <= 32'b00000000010000010000000100010011;
ROM[10572] <= 32'b00000000001100000000001110010011;
ROM[10573] <= 32'b11111111110000010000000100010011;
ROM[10574] <= 32'b00000000000000010010010000000011;
ROM[10575] <= 32'b00000000011101000000001110110011;
ROM[10576] <= 32'b11111111110000010000000100010011;
ROM[10577] <= 32'b00000000000000010010010000000011;
ROM[10578] <= 32'b00000000100000111010001110110011;
ROM[10579] <= 32'b00000000000000111000101001100011;
ROM[10580] <= 32'b00000000000000001010001110110111;
ROM[10581] <= 32'b01010110010000111000001110010011;
ROM[10582] <= 32'b00000000111000111000001110110011;
ROM[10583] <= 32'b00000000000000111000000011100111;
ROM[10584] <= 32'b00011111110000000000000011101111;
ROM[10585] <= 32'b00000000000000011010001110000011;
ROM[10586] <= 32'b00000000011100010010000000100011;
ROM[10587] <= 32'b00000000010000010000000100010011;
ROM[10588] <= 32'b00000000000000100010001110000011;
ROM[10589] <= 32'b11111111110000010000000100010011;
ROM[10590] <= 32'b00000000000000010010010000000011;
ROM[10591] <= 32'b00000000011101000000001110110011;
ROM[10592] <= 32'b00000000011100010010000000100011;
ROM[10593] <= 32'b00000000010000010000000100010011;
ROM[10594] <= 32'b00000000000000100010001110000011;
ROM[10595] <= 32'b11111111110000010000000100010011;
ROM[10596] <= 32'b00000000000000010010010000000011;
ROM[10597] <= 32'b00000000011101000000001110110011;
ROM[10598] <= 32'b00000000011100010010000000100011;
ROM[10599] <= 32'b00000000010000010000000100010011;
ROM[10600] <= 32'b00000000000000100010001110000011;
ROM[10601] <= 32'b11111111110000010000000100010011;
ROM[10602] <= 32'b00000000000000010010010000000011;
ROM[10603] <= 32'b00000000011101000000001110110011;
ROM[10604] <= 32'b00000000011100010010000000100011;
ROM[10605] <= 32'b00000000010000010000000100010011;
ROM[10606] <= 32'b00000000000000100010001110000011;
ROM[10607] <= 32'b11111111110000010000000100010011;
ROM[10608] <= 32'b00000000000000010010010000000011;
ROM[10609] <= 32'b00000000011101000000001110110011;
ROM[10610] <= 32'b00000000011100010010000000100011;
ROM[10611] <= 32'b00000000010000010000000100010011;
ROM[10612] <= 32'b00000000010000000000001110010011;
ROM[10613] <= 32'b11111111110000010000000100010011;
ROM[10614] <= 32'b00000000000000010010010000000011;
ROM[10615] <= 32'b00000000011101000000001110110011;
ROM[10616] <= 32'b00000000011100011010001000100011;
ROM[10617] <= 32'b00000110100001101010001110000011;
ROM[10618] <= 32'b00000000011100010010000000100011;
ROM[10619] <= 32'b00000000010000010000000100010011;
ROM[10620] <= 32'b00000000010000011010001110000011;
ROM[10621] <= 32'b11111111110000010000000100010011;
ROM[10622] <= 32'b00000000000000010010010000000011;
ROM[10623] <= 32'b00000000011101000000001110110011;
ROM[10624] <= 32'b00000000011100010010000000100011;
ROM[10625] <= 32'b00000000010000010000000100010011;
ROM[10626] <= 32'b00000110100001101010001110000011;
ROM[10627] <= 32'b00000000011100010010000000100011;
ROM[10628] <= 32'b00000000010000010000000100010011;
ROM[10629] <= 32'b00000000000000011010001110000011;
ROM[10630] <= 32'b11111111110000010000000100010011;
ROM[10631] <= 32'b00000000000000010010010000000011;
ROM[10632] <= 32'b00000000011101000000001110110011;
ROM[10633] <= 32'b00000000000000111000001100010011;
ROM[10634] <= 32'b00000000110100110000010000110011;
ROM[10635] <= 32'b00000000000001000010001110000011;
ROM[10636] <= 32'b00000000011101100010000000100011;
ROM[10637] <= 32'b11111111110000010000000100010011;
ROM[10638] <= 32'b00000000000000010010001110000011;
ROM[10639] <= 32'b00000000000000111000001100010011;
ROM[10640] <= 32'b00000000000001100010001110000011;
ROM[10641] <= 32'b00000000110100110000010000110011;
ROM[10642] <= 32'b00000000011101000010000000100011;
ROM[10643] <= 32'b00000110010001101010001110000011;
ROM[10644] <= 32'b00000000011100010010000000100011;
ROM[10645] <= 32'b00000000010000010000000100010011;
ROM[10646] <= 32'b00000000010000011010001110000011;
ROM[10647] <= 32'b11111111110000010000000100010011;
ROM[10648] <= 32'b00000000000000010010010000000011;
ROM[10649] <= 32'b00000000011101000000001110110011;
ROM[10650] <= 32'b00000000011100010010000000100011;
ROM[10651] <= 32'b00000000010000010000000100010011;
ROM[10652] <= 32'b00000110010001101010001110000011;
ROM[10653] <= 32'b00000000011100010010000000100011;
ROM[10654] <= 32'b00000000010000010000000100010011;
ROM[10655] <= 32'b00000000000000011010001110000011;
ROM[10656] <= 32'b11111111110000010000000100010011;
ROM[10657] <= 32'b00000000000000010010010000000011;
ROM[10658] <= 32'b00000000011101000000001110110011;
ROM[10659] <= 32'b00000000000000111000001100010011;
ROM[10660] <= 32'b00000000110100110000010000110011;
ROM[10661] <= 32'b00000000000001000010001110000011;
ROM[10662] <= 32'b00000000011100010010000000100011;
ROM[10663] <= 32'b00000000010000010000000100010011;
ROM[10664] <= 32'b00000000000000100010001110000011;
ROM[10665] <= 32'b11111111110000010000000100010011;
ROM[10666] <= 32'b00000000000000010010010000000011;
ROM[10667] <= 32'b01000000011101000000001110110011;
ROM[10668] <= 32'b00000000011100010010000000100011;
ROM[10669] <= 32'b00000000010000010000000100010011;
ROM[10670] <= 32'b00000000000100000000001110010011;
ROM[10671] <= 32'b11111111110000010000000100010011;
ROM[10672] <= 32'b00000000000000010010010000000011;
ROM[10673] <= 32'b01000000011101000000001110110011;
ROM[10674] <= 32'b00000000011101100010000000100011;
ROM[10675] <= 32'b11111111110000010000000100010011;
ROM[10676] <= 32'b00000000000000010010001110000011;
ROM[10677] <= 32'b00000000000000111000001100010011;
ROM[10678] <= 32'b00000000000001100010001110000011;
ROM[10679] <= 32'b00000000110100110000010000110011;
ROM[10680] <= 32'b00000000011101000010000000100011;
ROM[10681] <= 32'b00000110110001101010001110000011;
ROM[10682] <= 32'b00000000011100010010000000100011;
ROM[10683] <= 32'b00000000010000010000000100010011;
ROM[10684] <= 32'b00000000100000011010001110000011;
ROM[10685] <= 32'b11111111110000010000000100010011;
ROM[10686] <= 32'b00000000000000010010010000000011;
ROM[10687] <= 32'b00000000011101000000001110110011;
ROM[10688] <= 32'b00000000011100010010000000100011;
ROM[10689] <= 32'b00000000010000010000000100010011;
ROM[10690] <= 32'b00000000000000100010001110000011;
ROM[10691] <= 32'b00000000011100010010000000100011;
ROM[10692] <= 32'b00000000010000010000000100010011;
ROM[10693] <= 32'b00000000000100000000001110010011;
ROM[10694] <= 32'b11111111110000010000000100010011;
ROM[10695] <= 32'b00000000000000010010010000000011;
ROM[10696] <= 32'b00000000011101000000001110110011;
ROM[10697] <= 32'b00000000011101100010000000100011;
ROM[10698] <= 32'b11111111110000010000000100010011;
ROM[10699] <= 32'b00000000000000010010001110000011;
ROM[10700] <= 32'b00000000000000111000001100010011;
ROM[10701] <= 32'b00000000000001100010001110000011;
ROM[10702] <= 32'b00000000110100110000010000110011;
ROM[10703] <= 32'b00000000011101000010000000100011;
ROM[10704] <= 32'b00000000100000011010001110000011;
ROM[10705] <= 32'b00000110011101101010101000100011;
ROM[10706] <= 32'b00000000010000011010001110000011;
ROM[10707] <= 32'b00000110011101101010000000100011;
ROM[10708] <= 32'b00000000000100000000001110010011;
ROM[10709] <= 32'b00000110011101101010110000100011;
ROM[10710] <= 32'b00001010000000000000000011101111;
ROM[10711] <= 32'b00000110100001101010001110000011;
ROM[10712] <= 32'b00000000011100010010000000100011;
ROM[10713] <= 32'b00000000010000010000000100010011;
ROM[10714] <= 32'b00000000000000011010001110000011;
ROM[10715] <= 32'b11111111110000010000000100010011;
ROM[10716] <= 32'b00000000000000010010010000000011;
ROM[10717] <= 32'b00000000011101000000001110110011;
ROM[10718] <= 32'b00000000000000111000001100010011;
ROM[10719] <= 32'b00000000110100110000010000110011;
ROM[10720] <= 32'b00000000000001000010001110000011;
ROM[10721] <= 32'b00000000011100011010001000100011;
ROM[10722] <= 32'b00000110110001101010001110000011;
ROM[10723] <= 32'b00000000011100010010000000100011;
ROM[10724] <= 32'b00000000010000010000000100010011;
ROM[10725] <= 32'b00000000100000011010001110000011;
ROM[10726] <= 32'b11111111110000010000000100010011;
ROM[10727] <= 32'b00000000000000010010010000000011;
ROM[10728] <= 32'b00000000011101000000001110110011;
ROM[10729] <= 32'b00000000011100010010000000100011;
ROM[10730] <= 32'b00000000010000010000000100010011;
ROM[10731] <= 32'b00000110010001101010001110000011;
ROM[10732] <= 32'b00000000011100010010000000100011;
ROM[10733] <= 32'b00000000010000010000000100010011;
ROM[10734] <= 32'b00000000000000011010001110000011;
ROM[10735] <= 32'b11111111110000010000000100010011;
ROM[10736] <= 32'b00000000000000010010010000000011;
ROM[10737] <= 32'b00000000011101000000001110110011;
ROM[10738] <= 32'b00000000000000111000001100010011;
ROM[10739] <= 32'b00000000110100110000010000110011;
ROM[10740] <= 32'b00000000000001000010001110000011;
ROM[10741] <= 32'b00000000011101100010000000100011;
ROM[10742] <= 32'b11111111110000010000000100010011;
ROM[10743] <= 32'b00000000000000010010001110000011;
ROM[10744] <= 32'b00000000000000111000001100010011;
ROM[10745] <= 32'b00000000000001100010001110000011;
ROM[10746] <= 32'b00000000110100110000010000110011;
ROM[10747] <= 32'b00000000011101000010000000100011;
ROM[10748] <= 32'b00000000001000000000001110010011;
ROM[10749] <= 32'b00000110011101101010110000100011;
ROM[10750] <= 32'b00000000010000000000000011101111;
ROM[10751] <= 32'b00000000100000011010001110000011;
ROM[10752] <= 32'b00000000011100010010000000100011;
ROM[10753] <= 32'b00000000010000010000000100010011;
ROM[10754] <= 32'b00000001010000000000001110010011;
ROM[10755] <= 32'b01000000011100011000001110110011;
ROM[10756] <= 32'b00000000000000111010000010000011;
ROM[10757] <= 32'b11111111110000010000000100010011;
ROM[10758] <= 32'b00000000000000010010001110000011;
ROM[10759] <= 32'b00000000011100100010000000100011;
ROM[10760] <= 32'b00000000010000100000000100010011;
ROM[10761] <= 32'b00000001010000000000001110010011;
ROM[10762] <= 32'b01000000011100011000001110110011;
ROM[10763] <= 32'b00000000010000111010000110000011;
ROM[10764] <= 32'b00000000100000111010001000000011;
ROM[10765] <= 32'b00000000110000111010001010000011;
ROM[10766] <= 32'b00000001000000111010001100000011;
ROM[10767] <= 32'b00000000000000001000000011100111;
ROM[10768] <= 32'b00000000000000010010000000100011;
ROM[10769] <= 32'b00000000010000010000000100010011;
ROM[10770] <= 32'b00000000110000000000001110010011;
ROM[10771] <= 32'b00000000011100010010000000100011;
ROM[10772] <= 32'b00000000010000010000000100010011;
ROM[10773] <= 32'b00000000000000001011001110110111;
ROM[10774] <= 32'b10001010000000111000001110010011;
ROM[10775] <= 32'b00000000111000111000001110110011;
ROM[10776] <= 32'b00000000011100010010000000100011;
ROM[10777] <= 32'b00000000010000010000000100010011;
ROM[10778] <= 32'b00000000001100010010000000100011;
ROM[10779] <= 32'b00000000010000010000000100010011;
ROM[10780] <= 32'b00000000010000010010000000100011;
ROM[10781] <= 32'b00000000010000010000000100010011;
ROM[10782] <= 32'b00000000010100010010000000100011;
ROM[10783] <= 32'b00000000010000010000000100010011;
ROM[10784] <= 32'b00000000011000010010000000100011;
ROM[10785] <= 32'b00000000010000010000000100010011;
ROM[10786] <= 32'b00000001010000000000001110010011;
ROM[10787] <= 32'b00000000010000111000001110010011;
ROM[10788] <= 32'b01000000011100010000001110110011;
ROM[10789] <= 32'b00000000011100000000001000110011;
ROM[10790] <= 32'b00000000001000000000000110110011;
ROM[10791] <= 32'b11010110000111111110000011101111;
ROM[10792] <= 32'b11111111110000010000000100010011;
ROM[10793] <= 32'b00000000000000010010001110000011;
ROM[10794] <= 32'b00000000011100011010000000100011;
ROM[10795] <= 32'b00000010001000000000001110010011;
ROM[10796] <= 32'b00000000011100010010000000100011;
ROM[10797] <= 32'b00000000010000010000000100010011;
ROM[10798] <= 32'b00000000000000011010001110000011;
ROM[10799] <= 32'b00000000011100010010000000100011;
ROM[10800] <= 32'b00000000010000010000000100010011;
ROM[10801] <= 32'b00000000000000001011001110110111;
ROM[10802] <= 32'b10010001000000111000001110010011;
ROM[10803] <= 32'b00000000111000111000001110110011;
ROM[10804] <= 32'b00000000011100010010000000100011;
ROM[10805] <= 32'b00000000010000010000000100010011;
ROM[10806] <= 32'b00000000001100010010000000100011;
ROM[10807] <= 32'b00000000010000010000000100010011;
ROM[10808] <= 32'b00000000010000010010000000100011;
ROM[10809] <= 32'b00000000010000010000000100010011;
ROM[10810] <= 32'b00000000010100010010000000100011;
ROM[10811] <= 32'b00000000010000010000000100010011;
ROM[10812] <= 32'b00000000011000010010000000100011;
ROM[10813] <= 32'b00000000010000010000000100010011;
ROM[10814] <= 32'b00000001010000000000001110010011;
ROM[10815] <= 32'b00000000100000111000001110010011;
ROM[10816] <= 32'b01000000011100010000001110110011;
ROM[10817] <= 32'b00000000011100000000001000110011;
ROM[10818] <= 32'b00000000001000000000000110110011;
ROM[10819] <= 32'b11111100100011111110000011101111;
ROM[10820] <= 32'b11111111110000010000000100010011;
ROM[10821] <= 32'b00000000000000010010001110000011;
ROM[10822] <= 32'b00000000011100011010000000100011;
ROM[10823] <= 32'b00000000000000011010001110000011;
ROM[10824] <= 32'b00000000011100010010000000100011;
ROM[10825] <= 32'b00000000010000010000000100010011;
ROM[10826] <= 32'b01011000000000000000001110010011;
ROM[10827] <= 32'b11111111110000010000000100010011;
ROM[10828] <= 32'b00000000000000010010010000000011;
ROM[10829] <= 32'b00000000011101000000001110110011;
ROM[10830] <= 32'b00000000011100011010000000100011;
ROM[10831] <= 32'b00000000000000000000001110010011;
ROM[10832] <= 32'b00000000011100010010000000100011;
ROM[10833] <= 32'b00000000010000010000000100010011;
ROM[10834] <= 32'b00000000000000011010001110000011;
ROM[10835] <= 32'b11111111110000010000000100010011;
ROM[10836] <= 32'b00000000000000010010010000000011;
ROM[10837] <= 32'b01000000011101000000001110110011;
ROM[10838] <= 32'b00000110011101101010111000100011;
ROM[10839] <= 32'b00000000000000000000001110010011;
ROM[10840] <= 32'b00001000011101101010000000100011;
ROM[10841] <= 32'b00000000000000000000001110010011;
ROM[10842] <= 32'b00001000011101101010001000100011;
ROM[10843] <= 32'b00000000000000001011001110110111;
ROM[10844] <= 32'b10011011100000111000001110010011;
ROM[10845] <= 32'b00000000111000111000001110110011;
ROM[10846] <= 32'b00000000011100010010000000100011;
ROM[10847] <= 32'b00000000010000010000000100010011;
ROM[10848] <= 32'b00000000001100010010000000100011;
ROM[10849] <= 32'b00000000010000010000000100010011;
ROM[10850] <= 32'b00000000010000010010000000100011;
ROM[10851] <= 32'b00000000010000010000000100010011;
ROM[10852] <= 32'b00000000010100010010000000100011;
ROM[10853] <= 32'b00000000010000010000000100010011;
ROM[10854] <= 32'b00000000011000010010000000100011;
ROM[10855] <= 32'b00000000010000010000000100010011;
ROM[10856] <= 32'b00000001010000000000001110010011;
ROM[10857] <= 32'b00000000000000111000001110010011;
ROM[10858] <= 32'b01000000011100010000001110110011;
ROM[10859] <= 32'b00000000011100000000001000110011;
ROM[10860] <= 32'b00000000001000000000000110110011;
ROM[10861] <= 32'b00000101010000000000000011101111;
ROM[10862] <= 32'b11111111110000010000000100010011;
ROM[10863] <= 32'b00000000000000010010001110000011;
ROM[10864] <= 32'b00000000011101100010000000100011;
ROM[10865] <= 32'b00000000000000000000001110010011;
ROM[10866] <= 32'b00000000011100010010000000100011;
ROM[10867] <= 32'b00000000010000010000000100010011;
ROM[10868] <= 32'b00000001010000000000001110010011;
ROM[10869] <= 32'b01000000011100011000001110110011;
ROM[10870] <= 32'b00000000000000111010000010000011;
ROM[10871] <= 32'b11111111110000010000000100010011;
ROM[10872] <= 32'b00000000000000010010001110000011;
ROM[10873] <= 32'b00000000011100100010000000100011;
ROM[10874] <= 32'b00000000010000100000000100010011;
ROM[10875] <= 32'b00000001010000000000001110010011;
ROM[10876] <= 32'b01000000011100011000001110110011;
ROM[10877] <= 32'b00000000010000111010000110000011;
ROM[10878] <= 32'b00000000100000111010001000000011;
ROM[10879] <= 32'b00000000110000111010001010000011;
ROM[10880] <= 32'b00000001000000111010001100000011;
ROM[10881] <= 32'b00000000000000001000000011100111;
ROM[10882] <= 32'b00000000000000010010000000100011;
ROM[10883] <= 32'b00000000010000010000000100010011;
ROM[10884] <= 32'b00000111111100000000001110010011;
ROM[10885] <= 32'b00000000011100010010000000100011;
ROM[10886] <= 32'b00000000010000010000000100010011;
ROM[10887] <= 32'b00000000000000001011001110110111;
ROM[10888] <= 32'b10100110100000111000001110010011;
ROM[10889] <= 32'b00000000111000111000001110110011;
ROM[10890] <= 32'b00000000011100010010000000100011;
ROM[10891] <= 32'b00000000010000010000000100010011;
ROM[10892] <= 32'b00000000001100010010000000100011;
ROM[10893] <= 32'b00000000010000010000000100010011;
ROM[10894] <= 32'b00000000010000010010000000100011;
ROM[10895] <= 32'b00000000010000010000000100010011;
ROM[10896] <= 32'b00000000010100010010000000100011;
ROM[10897] <= 32'b00000000010000010000000100010011;
ROM[10898] <= 32'b00000000011000010010000000100011;
ROM[10899] <= 32'b00000000010000010000000100010011;
ROM[10900] <= 32'b00000001010000000000001110010011;
ROM[10901] <= 32'b00000000010000111000001110010011;
ROM[10902] <= 32'b01000000011100010000001110110011;
ROM[10903] <= 32'b00000000011100000000001000110011;
ROM[10904] <= 32'b00000000001000000000000110110011;
ROM[10905] <= 32'b10011101110111110101000011101111;
ROM[10906] <= 32'b11111111110000010000000100010011;
ROM[10907] <= 32'b00000000000000010010001110000011;
ROM[10908] <= 32'b00001000011101101010010000100011;
ROM[10909] <= 32'b00000000000000000000001110010011;
ROM[10910] <= 32'b00000000011100010010000000100011;
ROM[10911] <= 32'b00000000010000010000000100010011;
ROM[10912] <= 32'b00000011111100000000001110010011;
ROM[10913] <= 32'b00000000011100010010000000100011;
ROM[10914] <= 32'b00000000010000010000000100010011;
ROM[10915] <= 32'b00000011111100000000001110010011;
ROM[10916] <= 32'b00000000011100010010000000100011;
ROM[10917] <= 32'b00000000010000010000000100010011;
ROM[10918] <= 32'b00000011111100000000001110010011;
ROM[10919] <= 32'b00000000011100010010000000100011;
ROM[10920] <= 32'b00000000010000010000000100010011;
ROM[10921] <= 32'b00000011111100000000001110010011;
ROM[10922] <= 32'b00000000011100010010000000100011;
ROM[10923] <= 32'b00000000010000010000000100010011;
ROM[10924] <= 32'b00000011111100000000001110010011;
ROM[10925] <= 32'b00000000011100010010000000100011;
ROM[10926] <= 32'b00000000010000010000000100010011;
ROM[10927] <= 32'b00000011111100000000001110010011;
ROM[10928] <= 32'b00000000011100010010000000100011;
ROM[10929] <= 32'b00000000010000010000000100010011;
ROM[10930] <= 32'b00000000000000000000001110010011;
ROM[10931] <= 32'b00000000011100010010000000100011;
ROM[10932] <= 32'b00000000010000010000000100010011;
ROM[10933] <= 32'b00000000000000000000001110010011;
ROM[10934] <= 32'b00000000011100010010000000100011;
ROM[10935] <= 32'b00000000010000010000000100010011;
ROM[10936] <= 32'b00000000000000001011001110110111;
ROM[10937] <= 32'b10110010110000111000001110010011;
ROM[10938] <= 32'b00000000111000111000001110110011;
ROM[10939] <= 32'b00000000011100010010000000100011;
ROM[10940] <= 32'b00000000010000010000000100010011;
ROM[10941] <= 32'b00000000001100010010000000100011;
ROM[10942] <= 32'b00000000010000010000000100010011;
ROM[10943] <= 32'b00000000010000010010000000100011;
ROM[10944] <= 32'b00000000010000010000000100010011;
ROM[10945] <= 32'b00000000010100010010000000100011;
ROM[10946] <= 32'b00000000010000010000000100010011;
ROM[10947] <= 32'b00000000011000010010000000100011;
ROM[10948] <= 32'b00000000010000010000000100010011;
ROM[10949] <= 32'b00000001010000000000001110010011;
ROM[10950] <= 32'b00000010010000111000001110010011;
ROM[10951] <= 32'b01000000011100010000001110110011;
ROM[10952] <= 32'b00000000011100000000001000110011;
ROM[10953] <= 32'b00000000001000000000000110110011;
ROM[10954] <= 32'b00010001000100000100000011101111;
ROM[10955] <= 32'b11111111110000010000000100010011;
ROM[10956] <= 32'b00000000000000010010001110000011;
ROM[10957] <= 32'b00000000011101100010000000100011;
ROM[10958] <= 32'b00000010000000000000001110010011;
ROM[10959] <= 32'b00000000011100010010000000100011;
ROM[10960] <= 32'b00000000010000010000000100010011;
ROM[10961] <= 32'b00000000000000000000001110010011;
ROM[10962] <= 32'b00000000011100010010000000100011;
ROM[10963] <= 32'b00000000010000010000000100010011;
ROM[10964] <= 32'b00000000000000000000001110010011;
ROM[10965] <= 32'b00000000011100010010000000100011;
ROM[10966] <= 32'b00000000010000010000000100010011;
ROM[10967] <= 32'b00000000000000000000001110010011;
ROM[10968] <= 32'b00000000011100010010000000100011;
ROM[10969] <= 32'b00000000010000010000000100010011;
ROM[10970] <= 32'b00000000000000000000001110010011;
ROM[10971] <= 32'b00000000011100010010000000100011;
ROM[10972] <= 32'b00000000010000010000000100010011;
ROM[10973] <= 32'b00000000000000000000001110010011;
ROM[10974] <= 32'b00000000011100010010000000100011;
ROM[10975] <= 32'b00000000010000010000000100010011;
ROM[10976] <= 32'b00000000000000000000001110010011;
ROM[10977] <= 32'b00000000011100010010000000100011;
ROM[10978] <= 32'b00000000010000010000000100010011;
ROM[10979] <= 32'b00000000000000000000001110010011;
ROM[10980] <= 32'b00000000011100010010000000100011;
ROM[10981] <= 32'b00000000010000010000000100010011;
ROM[10982] <= 32'b00000000000000000000001110010011;
ROM[10983] <= 32'b00000000011100010010000000100011;
ROM[10984] <= 32'b00000000010000010000000100010011;
ROM[10985] <= 32'b00000000000000001011001110110111;
ROM[10986] <= 32'b10111111000000111000001110010011;
ROM[10987] <= 32'b00000000111000111000001110110011;
ROM[10988] <= 32'b00000000011100010010000000100011;
ROM[10989] <= 32'b00000000010000010000000100010011;
ROM[10990] <= 32'b00000000001100010010000000100011;
ROM[10991] <= 32'b00000000010000010000000100010011;
ROM[10992] <= 32'b00000000010000010010000000100011;
ROM[10993] <= 32'b00000000010000010000000100010011;
ROM[10994] <= 32'b00000000010100010010000000100011;
ROM[10995] <= 32'b00000000010000010000000100010011;
ROM[10996] <= 32'b00000000011000010010000000100011;
ROM[10997] <= 32'b00000000010000010000000100010011;
ROM[10998] <= 32'b00000001010000000000001110010011;
ROM[10999] <= 32'b00000010010000111000001110010011;
ROM[11000] <= 32'b01000000011100010000001110110011;
ROM[11001] <= 32'b00000000011100000000001000110011;
ROM[11002] <= 32'b00000000001000000000000110110011;
ROM[11003] <= 32'b00000100110100000100000011101111;
ROM[11004] <= 32'b11111111110000010000000100010011;
ROM[11005] <= 32'b00000000000000010010001110000011;
ROM[11006] <= 32'b00000000011101100010000000100011;
ROM[11007] <= 32'b00000010000100000000001110010011;
ROM[11008] <= 32'b00000000011100010010000000100011;
ROM[11009] <= 32'b00000000010000010000000100010011;
ROM[11010] <= 32'b00000001100000000000001110010011;
ROM[11011] <= 32'b00000000011100010010000000100011;
ROM[11012] <= 32'b00000000010000010000000100010011;
ROM[11013] <= 32'b00000011110000000000001110010011;
ROM[11014] <= 32'b00000000011100010010000000100011;
ROM[11015] <= 32'b00000000010000010000000100010011;
ROM[11016] <= 32'b00000011110000000000001110010011;
ROM[11017] <= 32'b00000000011100010010000000100011;
ROM[11018] <= 32'b00000000010000010000000100010011;
ROM[11019] <= 32'b00000001100000000000001110010011;
ROM[11020] <= 32'b00000000011100010010000000100011;
ROM[11021] <= 32'b00000000010000010000000100010011;
ROM[11022] <= 32'b00000001100000000000001110010011;
ROM[11023] <= 32'b00000000011100010010000000100011;
ROM[11024] <= 32'b00000000010000010000000100010011;
ROM[11025] <= 32'b00000000000000000000001110010011;
ROM[11026] <= 32'b00000000011100010010000000100011;
ROM[11027] <= 32'b00000000010000010000000100010011;
ROM[11028] <= 32'b00000001100000000000001110010011;
ROM[11029] <= 32'b00000000011100010010000000100011;
ROM[11030] <= 32'b00000000010000010000000100010011;
ROM[11031] <= 32'b00000000000000000000001110010011;
ROM[11032] <= 32'b00000000011100010010000000100011;
ROM[11033] <= 32'b00000000010000010000000100010011;
ROM[11034] <= 32'b00000000000000001011001110110111;
ROM[11035] <= 32'b11001011010000111000001110010011;
ROM[11036] <= 32'b00000000111000111000001110110011;
ROM[11037] <= 32'b00000000011100010010000000100011;
ROM[11038] <= 32'b00000000010000010000000100010011;
ROM[11039] <= 32'b00000000001100010010000000100011;
ROM[11040] <= 32'b00000000010000010000000100010011;
ROM[11041] <= 32'b00000000010000010010000000100011;
ROM[11042] <= 32'b00000000010000010000000100010011;
ROM[11043] <= 32'b00000000010100010010000000100011;
ROM[11044] <= 32'b00000000010000010000000100010011;
ROM[11045] <= 32'b00000000011000010010000000100011;
ROM[11046] <= 32'b00000000010000010000000100010011;
ROM[11047] <= 32'b00000001010000000000001110010011;
ROM[11048] <= 32'b00000010010000111000001110010011;
ROM[11049] <= 32'b01000000011100010000001110110011;
ROM[11050] <= 32'b00000000011100000000001000110011;
ROM[11051] <= 32'b00000000001000000000000110110011;
ROM[11052] <= 32'b01111000100000000100000011101111;
ROM[11053] <= 32'b11111111110000010000000100010011;
ROM[11054] <= 32'b00000000000000010010001110000011;
ROM[11055] <= 32'b00000000011101100010000000100011;
ROM[11056] <= 32'b00000010001000000000001110010011;
ROM[11057] <= 32'b00000000011100010010000000100011;
ROM[11058] <= 32'b00000000010000010000000100010011;
ROM[11059] <= 32'b00000110110000000000001110010011;
ROM[11060] <= 32'b00000000011100010010000000100011;
ROM[11061] <= 32'b00000000010000010000000100010011;
ROM[11062] <= 32'b00000110110000000000001110010011;
ROM[11063] <= 32'b00000000011100010010000000100011;
ROM[11064] <= 32'b00000000010000010000000100010011;
ROM[11065] <= 32'b00000000000000000000001110010011;
ROM[11066] <= 32'b00000000011100010010000000100011;
ROM[11067] <= 32'b00000000010000010000000100010011;
ROM[11068] <= 32'b00000000000000000000001110010011;
ROM[11069] <= 32'b00000000011100010010000000100011;
ROM[11070] <= 32'b00000000010000010000000100010011;
ROM[11071] <= 32'b00000000000000000000001110010011;
ROM[11072] <= 32'b00000000011100010010000000100011;
ROM[11073] <= 32'b00000000010000010000000100010011;
ROM[11074] <= 32'b00000000000000000000001110010011;
ROM[11075] <= 32'b00000000011100010010000000100011;
ROM[11076] <= 32'b00000000010000010000000100010011;
ROM[11077] <= 32'b00000000000000000000001110010011;
ROM[11078] <= 32'b00000000011100010010000000100011;
ROM[11079] <= 32'b00000000010000010000000100010011;
ROM[11080] <= 32'b00000000000000000000001110010011;
ROM[11081] <= 32'b00000000011100010010000000100011;
ROM[11082] <= 32'b00000000010000010000000100010011;
ROM[11083] <= 32'b00000000000000001011001110110111;
ROM[11084] <= 32'b11010111100000111000001110010011;
ROM[11085] <= 32'b00000000111000111000001110110011;
ROM[11086] <= 32'b00000000011100010010000000100011;
ROM[11087] <= 32'b00000000010000010000000100010011;
ROM[11088] <= 32'b00000000001100010010000000100011;
ROM[11089] <= 32'b00000000010000010000000100010011;
ROM[11090] <= 32'b00000000010000010010000000100011;
ROM[11091] <= 32'b00000000010000010000000100010011;
ROM[11092] <= 32'b00000000010100010010000000100011;
ROM[11093] <= 32'b00000000010000010000000100010011;
ROM[11094] <= 32'b00000000011000010010000000100011;
ROM[11095] <= 32'b00000000010000010000000100010011;
ROM[11096] <= 32'b00000001010000000000001110010011;
ROM[11097] <= 32'b00000010010000111000001110010011;
ROM[11098] <= 32'b01000000011100010000001110110011;
ROM[11099] <= 32'b00000000011100000000001000110011;
ROM[11100] <= 32'b00000000001000000000000110110011;
ROM[11101] <= 32'b01101100010000000100000011101111;
ROM[11102] <= 32'b11111111110000010000000100010011;
ROM[11103] <= 32'b00000000000000010010001110000011;
ROM[11104] <= 32'b00000000011101100010000000100011;
ROM[11105] <= 32'b00000010001100000000001110010011;
ROM[11106] <= 32'b00000000011100010010000000100011;
ROM[11107] <= 32'b00000000010000010000000100010011;
ROM[11108] <= 32'b00000110110000000000001110010011;
ROM[11109] <= 32'b00000000011100010010000000100011;
ROM[11110] <= 32'b00000000010000010000000100010011;
ROM[11111] <= 32'b00000110110000000000001110010011;
ROM[11112] <= 32'b00000000011100010010000000100011;
ROM[11113] <= 32'b00000000010000010000000100010011;
ROM[11114] <= 32'b00001111111000000000001110010011;
ROM[11115] <= 32'b00000000011100010010000000100011;
ROM[11116] <= 32'b00000000010000010000000100010011;
ROM[11117] <= 32'b00000110110000000000001110010011;
ROM[11118] <= 32'b00000000011100010010000000100011;
ROM[11119] <= 32'b00000000010000010000000100010011;
ROM[11120] <= 32'b00001111111000000000001110010011;
ROM[11121] <= 32'b00000000011100010010000000100011;
ROM[11122] <= 32'b00000000010000010000000100010011;
ROM[11123] <= 32'b00000110110000000000001110010011;
ROM[11124] <= 32'b00000000011100010010000000100011;
ROM[11125] <= 32'b00000000010000010000000100010011;
ROM[11126] <= 32'b00000110110000000000001110010011;
ROM[11127] <= 32'b00000000011100010010000000100011;
ROM[11128] <= 32'b00000000010000010000000100010011;
ROM[11129] <= 32'b00000000000000000000001110010011;
ROM[11130] <= 32'b00000000011100010010000000100011;
ROM[11131] <= 32'b00000000010000010000000100010011;
ROM[11132] <= 32'b00000000000000001011001110110111;
ROM[11133] <= 32'b11100011110000111000001110010011;
ROM[11134] <= 32'b00000000111000111000001110110011;
ROM[11135] <= 32'b00000000011100010010000000100011;
ROM[11136] <= 32'b00000000010000010000000100010011;
ROM[11137] <= 32'b00000000001100010010000000100011;
ROM[11138] <= 32'b00000000010000010000000100010011;
ROM[11139] <= 32'b00000000010000010010000000100011;
ROM[11140] <= 32'b00000000010000010000000100010011;
ROM[11141] <= 32'b00000000010100010010000000100011;
ROM[11142] <= 32'b00000000010000010000000100010011;
ROM[11143] <= 32'b00000000011000010010000000100011;
ROM[11144] <= 32'b00000000010000010000000100010011;
ROM[11145] <= 32'b00000001010000000000001110010011;
ROM[11146] <= 32'b00000010010000111000001110010011;
ROM[11147] <= 32'b01000000011100010000001110110011;
ROM[11148] <= 32'b00000000011100000000001000110011;
ROM[11149] <= 32'b00000000001000000000000110110011;
ROM[11150] <= 32'b01100000000000000100000011101111;
ROM[11151] <= 32'b11111111110000010000000100010011;
ROM[11152] <= 32'b00000000000000010010001110000011;
ROM[11153] <= 32'b00000000011101100010000000100011;
ROM[11154] <= 32'b00000010010000000000001110010011;
ROM[11155] <= 32'b00000000011100010010000000100011;
ROM[11156] <= 32'b00000000010000010000000100010011;
ROM[11157] <= 32'b00000011000000000000001110010011;
ROM[11158] <= 32'b00000000011100010010000000100011;
ROM[11159] <= 32'b00000000010000010000000100010011;
ROM[11160] <= 32'b00000111110000000000001110010011;
ROM[11161] <= 32'b00000000011100010010000000100011;
ROM[11162] <= 32'b00000000010000010000000100010011;
ROM[11163] <= 32'b00001100000000000000001110010011;
ROM[11164] <= 32'b00000000011100010010000000100011;
ROM[11165] <= 32'b00000000010000010000000100010011;
ROM[11166] <= 32'b00000111100000000000001110010011;
ROM[11167] <= 32'b00000000011100010010000000100011;
ROM[11168] <= 32'b00000000010000010000000100010011;
ROM[11169] <= 32'b00000000110000000000001110010011;
ROM[11170] <= 32'b00000000011100010010000000100011;
ROM[11171] <= 32'b00000000010000010000000100010011;
ROM[11172] <= 32'b00001111100000000000001110010011;
ROM[11173] <= 32'b00000000011100010010000000100011;
ROM[11174] <= 32'b00000000010000010000000100010011;
ROM[11175] <= 32'b00000011000000000000001110010011;
ROM[11176] <= 32'b00000000011100010010000000100011;
ROM[11177] <= 32'b00000000010000010000000100010011;
ROM[11178] <= 32'b00000000000000000000001110010011;
ROM[11179] <= 32'b00000000011100010010000000100011;
ROM[11180] <= 32'b00000000010000010000000100010011;
ROM[11181] <= 32'b00000000000000001011001110110111;
ROM[11182] <= 32'b11110000000000111000001110010011;
ROM[11183] <= 32'b00000000111000111000001110110011;
ROM[11184] <= 32'b00000000011100010010000000100011;
ROM[11185] <= 32'b00000000010000010000000100010011;
ROM[11186] <= 32'b00000000001100010010000000100011;
ROM[11187] <= 32'b00000000010000010000000100010011;
ROM[11188] <= 32'b00000000010000010010000000100011;
ROM[11189] <= 32'b00000000010000010000000100010011;
ROM[11190] <= 32'b00000000010100010010000000100011;
ROM[11191] <= 32'b00000000010000010000000100010011;
ROM[11192] <= 32'b00000000011000010010000000100011;
ROM[11193] <= 32'b00000000010000010000000100010011;
ROM[11194] <= 32'b00000001010000000000001110010011;
ROM[11195] <= 32'b00000010010000111000001110010011;
ROM[11196] <= 32'b01000000011100010000001110110011;
ROM[11197] <= 32'b00000000011100000000001000110011;
ROM[11198] <= 32'b00000000001000000000000110110011;
ROM[11199] <= 32'b01010011110000000100000011101111;
ROM[11200] <= 32'b11111111110000010000000100010011;
ROM[11201] <= 32'b00000000000000010010001110000011;
ROM[11202] <= 32'b00000000011101100010000000100011;
ROM[11203] <= 32'b00000010010100000000001110010011;
ROM[11204] <= 32'b00000000011100010010000000100011;
ROM[11205] <= 32'b00000000010000010000000100010011;
ROM[11206] <= 32'b00000000000000000000001110010011;
ROM[11207] <= 32'b00000000011100010010000000100011;
ROM[11208] <= 32'b00000000010000010000000100010011;
ROM[11209] <= 32'b00001100011000000000001110010011;
ROM[11210] <= 32'b00000000011100010010000000100011;
ROM[11211] <= 32'b00000000010000010000000100010011;
ROM[11212] <= 32'b00001100110000000000001110010011;
ROM[11213] <= 32'b00000000011100010010000000100011;
ROM[11214] <= 32'b00000000010000010000000100010011;
ROM[11215] <= 32'b00000001100000000000001110010011;
ROM[11216] <= 32'b00000000011100010010000000100011;
ROM[11217] <= 32'b00000000010000010000000100010011;
ROM[11218] <= 32'b00000011000000000000001110010011;
ROM[11219] <= 32'b00000000011100010010000000100011;
ROM[11220] <= 32'b00000000010000010000000100010011;
ROM[11221] <= 32'b00000110011000000000001110010011;
ROM[11222] <= 32'b00000000011100010010000000100011;
ROM[11223] <= 32'b00000000010000010000000100010011;
ROM[11224] <= 32'b00001100011000000000001110010011;
ROM[11225] <= 32'b00000000011100010010000000100011;
ROM[11226] <= 32'b00000000010000010000000100010011;
ROM[11227] <= 32'b00000000000000000000001110010011;
ROM[11228] <= 32'b00000000011100010010000000100011;
ROM[11229] <= 32'b00000000010000010000000100010011;
ROM[11230] <= 32'b00000000000000001011001110110111;
ROM[11231] <= 32'b11111100010000111000001110010011;
ROM[11232] <= 32'b00000000111000111000001110110011;
ROM[11233] <= 32'b00000000011100010010000000100011;
ROM[11234] <= 32'b00000000010000010000000100010011;
ROM[11235] <= 32'b00000000001100010010000000100011;
ROM[11236] <= 32'b00000000010000010000000100010011;
ROM[11237] <= 32'b00000000010000010010000000100011;
ROM[11238] <= 32'b00000000010000010000000100010011;
ROM[11239] <= 32'b00000000010100010010000000100011;
ROM[11240] <= 32'b00000000010000010000000100010011;
ROM[11241] <= 32'b00000000011000010010000000100011;
ROM[11242] <= 32'b00000000010000010000000100010011;
ROM[11243] <= 32'b00000001010000000000001110010011;
ROM[11244] <= 32'b00000010010000111000001110010011;
ROM[11245] <= 32'b01000000011100010000001110110011;
ROM[11246] <= 32'b00000000011100000000001000110011;
ROM[11247] <= 32'b00000000001000000000000110110011;
ROM[11248] <= 32'b01000111100000000100000011101111;
ROM[11249] <= 32'b11111111110000010000000100010011;
ROM[11250] <= 32'b00000000000000010010001110000011;
ROM[11251] <= 32'b00000000011101100010000000100011;
ROM[11252] <= 32'b00000010011000000000001110010011;
ROM[11253] <= 32'b00000000011100010010000000100011;
ROM[11254] <= 32'b00000000010000010000000100010011;
ROM[11255] <= 32'b00000011100000000000001110010011;
ROM[11256] <= 32'b00000000011100010010000000100011;
ROM[11257] <= 32'b00000000010000010000000100010011;
ROM[11258] <= 32'b00000110110000000000001110010011;
ROM[11259] <= 32'b00000000011100010010000000100011;
ROM[11260] <= 32'b00000000010000010000000100010011;
ROM[11261] <= 32'b00000011100000000000001110010011;
ROM[11262] <= 32'b00000000011100010010000000100011;
ROM[11263] <= 32'b00000000010000010000000100010011;
ROM[11264] <= 32'b00000111011000000000001110010011;
ROM[11265] <= 32'b00000000011100010010000000100011;
ROM[11266] <= 32'b00000000010000010000000100010011;
ROM[11267] <= 32'b00001101110000000000001110010011;
ROM[11268] <= 32'b00000000011100010010000000100011;
ROM[11269] <= 32'b00000000010000010000000100010011;
ROM[11270] <= 32'b00001100110000000000001110010011;
ROM[11271] <= 32'b00000000011100010010000000100011;
ROM[11272] <= 32'b00000000010000010000000100010011;
ROM[11273] <= 32'b00000111011000000000001110010011;
ROM[11274] <= 32'b00000000011100010010000000100011;
ROM[11275] <= 32'b00000000010000010000000100010011;
ROM[11276] <= 32'b00000000000000000000001110010011;
ROM[11277] <= 32'b00000000011100010010000000100011;
ROM[11278] <= 32'b00000000010000010000000100010011;
ROM[11279] <= 32'b00000000000000001011001110110111;
ROM[11280] <= 32'b00001000100000111000001110010011;
ROM[11281] <= 32'b00000000111000111000001110110011;
ROM[11282] <= 32'b00000000011100010010000000100011;
ROM[11283] <= 32'b00000000010000010000000100010011;
ROM[11284] <= 32'b00000000001100010010000000100011;
ROM[11285] <= 32'b00000000010000010000000100010011;
ROM[11286] <= 32'b00000000010000010010000000100011;
ROM[11287] <= 32'b00000000010000010000000100010011;
ROM[11288] <= 32'b00000000010100010010000000100011;
ROM[11289] <= 32'b00000000010000010000000100010011;
ROM[11290] <= 32'b00000000011000010010000000100011;
ROM[11291] <= 32'b00000000010000010000000100010011;
ROM[11292] <= 32'b00000001010000000000001110010011;
ROM[11293] <= 32'b00000010010000111000001110010011;
ROM[11294] <= 32'b01000000011100010000001110110011;
ROM[11295] <= 32'b00000000011100000000001000110011;
ROM[11296] <= 32'b00000000001000000000000110110011;
ROM[11297] <= 32'b00111011010000000100000011101111;
ROM[11298] <= 32'b11111111110000010000000100010011;
ROM[11299] <= 32'b00000000000000010010001110000011;
ROM[11300] <= 32'b00000000011101100010000000100011;
ROM[11301] <= 32'b00000010011100000000001110010011;
ROM[11302] <= 32'b00000000011100010010000000100011;
ROM[11303] <= 32'b00000000010000010000000100010011;
ROM[11304] <= 32'b00000110000000000000001110010011;
ROM[11305] <= 32'b00000000011100010010000000100011;
ROM[11306] <= 32'b00000000010000010000000100010011;
ROM[11307] <= 32'b00000110000000000000001110010011;
ROM[11308] <= 32'b00000000011100010010000000100011;
ROM[11309] <= 32'b00000000010000010000000100010011;
ROM[11310] <= 32'b00001100000000000000001110010011;
ROM[11311] <= 32'b00000000011100010010000000100011;
ROM[11312] <= 32'b00000000010000010000000100010011;
ROM[11313] <= 32'b00000000000000000000001110010011;
ROM[11314] <= 32'b00000000011100010010000000100011;
ROM[11315] <= 32'b00000000010000010000000100010011;
ROM[11316] <= 32'b00000000000000000000001110010011;
ROM[11317] <= 32'b00000000011100010010000000100011;
ROM[11318] <= 32'b00000000010000010000000100010011;
ROM[11319] <= 32'b00000000000000000000001110010011;
ROM[11320] <= 32'b00000000011100010010000000100011;
ROM[11321] <= 32'b00000000010000010000000100010011;
ROM[11322] <= 32'b00000000000000000000001110010011;
ROM[11323] <= 32'b00000000011100010010000000100011;
ROM[11324] <= 32'b00000000010000010000000100010011;
ROM[11325] <= 32'b00000000000000000000001110010011;
ROM[11326] <= 32'b00000000011100010010000000100011;
ROM[11327] <= 32'b00000000010000010000000100010011;
ROM[11328] <= 32'b00000000000000001011001110110111;
ROM[11329] <= 32'b00010100110000111000001110010011;
ROM[11330] <= 32'b00000000111000111000001110110011;
ROM[11331] <= 32'b00000000011100010010000000100011;
ROM[11332] <= 32'b00000000010000010000000100010011;
ROM[11333] <= 32'b00000000001100010010000000100011;
ROM[11334] <= 32'b00000000010000010000000100010011;
ROM[11335] <= 32'b00000000010000010010000000100011;
ROM[11336] <= 32'b00000000010000010000000100010011;
ROM[11337] <= 32'b00000000010100010010000000100011;
ROM[11338] <= 32'b00000000010000010000000100010011;
ROM[11339] <= 32'b00000000011000010010000000100011;
ROM[11340] <= 32'b00000000010000010000000100010011;
ROM[11341] <= 32'b00000001010000000000001110010011;
ROM[11342] <= 32'b00000010010000111000001110010011;
ROM[11343] <= 32'b01000000011100010000001110110011;
ROM[11344] <= 32'b00000000011100000000001000110011;
ROM[11345] <= 32'b00000000001000000000000110110011;
ROM[11346] <= 32'b00101111000000000100000011101111;
ROM[11347] <= 32'b11111111110000010000000100010011;
ROM[11348] <= 32'b00000000000000010010001110000011;
ROM[11349] <= 32'b00000000011101100010000000100011;
ROM[11350] <= 32'b00000010100000000000001110010011;
ROM[11351] <= 32'b00000000011100010010000000100011;
ROM[11352] <= 32'b00000000010000010000000100010011;
ROM[11353] <= 32'b00000001100000000000001110010011;
ROM[11354] <= 32'b00000000011100010010000000100011;
ROM[11355] <= 32'b00000000010000010000000100010011;
ROM[11356] <= 32'b00000011000000000000001110010011;
ROM[11357] <= 32'b00000000011100010010000000100011;
ROM[11358] <= 32'b00000000010000010000000100010011;
ROM[11359] <= 32'b00000110000000000000001110010011;
ROM[11360] <= 32'b00000000011100010010000000100011;
ROM[11361] <= 32'b00000000010000010000000100010011;
ROM[11362] <= 32'b00000110000000000000001110010011;
ROM[11363] <= 32'b00000000011100010010000000100011;
ROM[11364] <= 32'b00000000010000010000000100010011;
ROM[11365] <= 32'b00000110000000000000001110010011;
ROM[11366] <= 32'b00000000011100010010000000100011;
ROM[11367] <= 32'b00000000010000010000000100010011;
ROM[11368] <= 32'b00000011000000000000001110010011;
ROM[11369] <= 32'b00000000011100010010000000100011;
ROM[11370] <= 32'b00000000010000010000000100010011;
ROM[11371] <= 32'b00000001100000000000001110010011;
ROM[11372] <= 32'b00000000011100010010000000100011;
ROM[11373] <= 32'b00000000010000010000000100010011;
ROM[11374] <= 32'b00000000000000000000001110010011;
ROM[11375] <= 32'b00000000011100010010000000100011;
ROM[11376] <= 32'b00000000010000010000000100010011;
ROM[11377] <= 32'b00000000000000001011001110110111;
ROM[11378] <= 32'b00100001000000111000001110010011;
ROM[11379] <= 32'b00000000111000111000001110110011;
ROM[11380] <= 32'b00000000011100010010000000100011;
ROM[11381] <= 32'b00000000010000010000000100010011;
ROM[11382] <= 32'b00000000001100010010000000100011;
ROM[11383] <= 32'b00000000010000010000000100010011;
ROM[11384] <= 32'b00000000010000010010000000100011;
ROM[11385] <= 32'b00000000010000010000000100010011;
ROM[11386] <= 32'b00000000010100010010000000100011;
ROM[11387] <= 32'b00000000010000010000000100010011;
ROM[11388] <= 32'b00000000011000010010000000100011;
ROM[11389] <= 32'b00000000010000010000000100010011;
ROM[11390] <= 32'b00000001010000000000001110010011;
ROM[11391] <= 32'b00000010010000111000001110010011;
ROM[11392] <= 32'b01000000011100010000001110110011;
ROM[11393] <= 32'b00000000011100000000001000110011;
ROM[11394] <= 32'b00000000001000000000000110110011;
ROM[11395] <= 32'b00100010110000000100000011101111;
ROM[11396] <= 32'b11111111110000010000000100010011;
ROM[11397] <= 32'b00000000000000010010001110000011;
ROM[11398] <= 32'b00000000011101100010000000100011;
ROM[11399] <= 32'b00000010100100000000001110010011;
ROM[11400] <= 32'b00000000011100010010000000100011;
ROM[11401] <= 32'b00000000010000010000000100010011;
ROM[11402] <= 32'b00000110000000000000001110010011;
ROM[11403] <= 32'b00000000011100010010000000100011;
ROM[11404] <= 32'b00000000010000010000000100010011;
ROM[11405] <= 32'b00000011000000000000001110010011;
ROM[11406] <= 32'b00000000011100010010000000100011;
ROM[11407] <= 32'b00000000010000010000000100010011;
ROM[11408] <= 32'b00000001100000000000001110010011;
ROM[11409] <= 32'b00000000011100010010000000100011;
ROM[11410] <= 32'b00000000010000010000000100010011;
ROM[11411] <= 32'b00000001100000000000001110010011;
ROM[11412] <= 32'b00000000011100010010000000100011;
ROM[11413] <= 32'b00000000010000010000000100010011;
ROM[11414] <= 32'b00000001100000000000001110010011;
ROM[11415] <= 32'b00000000011100010010000000100011;
ROM[11416] <= 32'b00000000010000010000000100010011;
ROM[11417] <= 32'b00000011000000000000001110010011;
ROM[11418] <= 32'b00000000011100010010000000100011;
ROM[11419] <= 32'b00000000010000010000000100010011;
ROM[11420] <= 32'b00000110000000000000001110010011;
ROM[11421] <= 32'b00000000011100010010000000100011;
ROM[11422] <= 32'b00000000010000010000000100010011;
ROM[11423] <= 32'b00000000000000000000001110010011;
ROM[11424] <= 32'b00000000011100010010000000100011;
ROM[11425] <= 32'b00000000010000010000000100010011;
ROM[11426] <= 32'b00000000000000001011001110110111;
ROM[11427] <= 32'b00101101010000111000001110010011;
ROM[11428] <= 32'b00000000111000111000001110110011;
ROM[11429] <= 32'b00000000011100010010000000100011;
ROM[11430] <= 32'b00000000010000010000000100010011;
ROM[11431] <= 32'b00000000001100010010000000100011;
ROM[11432] <= 32'b00000000010000010000000100010011;
ROM[11433] <= 32'b00000000010000010010000000100011;
ROM[11434] <= 32'b00000000010000010000000100010011;
ROM[11435] <= 32'b00000000010100010010000000100011;
ROM[11436] <= 32'b00000000010000010000000100010011;
ROM[11437] <= 32'b00000000011000010010000000100011;
ROM[11438] <= 32'b00000000010000010000000100010011;
ROM[11439] <= 32'b00000001010000000000001110010011;
ROM[11440] <= 32'b00000010010000111000001110010011;
ROM[11441] <= 32'b01000000011100010000001110110011;
ROM[11442] <= 32'b00000000011100000000001000110011;
ROM[11443] <= 32'b00000000001000000000000110110011;
ROM[11444] <= 32'b00010110100000000100000011101111;
ROM[11445] <= 32'b11111111110000010000000100010011;
ROM[11446] <= 32'b00000000000000010010001110000011;
ROM[11447] <= 32'b00000000011101100010000000100011;
ROM[11448] <= 32'b00000010101000000000001110010011;
ROM[11449] <= 32'b00000000011100010010000000100011;
ROM[11450] <= 32'b00000000010000010000000100010011;
ROM[11451] <= 32'b00000000000000000000001110010011;
ROM[11452] <= 32'b00000000011100010010000000100011;
ROM[11453] <= 32'b00000000010000010000000100010011;
ROM[11454] <= 32'b00000110011000000000001110010011;
ROM[11455] <= 32'b00000000011100010010000000100011;
ROM[11456] <= 32'b00000000010000010000000100010011;
ROM[11457] <= 32'b00000011110000000000001110010011;
ROM[11458] <= 32'b00000000011100010010000000100011;
ROM[11459] <= 32'b00000000010000010000000100010011;
ROM[11460] <= 32'b00001111111100000000001110010011;
ROM[11461] <= 32'b00000000011100010010000000100011;
ROM[11462] <= 32'b00000000010000010000000100010011;
ROM[11463] <= 32'b00000011110000000000001110010011;
ROM[11464] <= 32'b00000000011100010010000000100011;
ROM[11465] <= 32'b00000000010000010000000100010011;
ROM[11466] <= 32'b00000110011000000000001110010011;
ROM[11467] <= 32'b00000000011100010010000000100011;
ROM[11468] <= 32'b00000000010000010000000100010011;
ROM[11469] <= 32'b00000000000000000000001110010011;
ROM[11470] <= 32'b00000000011100010010000000100011;
ROM[11471] <= 32'b00000000010000010000000100010011;
ROM[11472] <= 32'b00000000000000000000001110010011;
ROM[11473] <= 32'b00000000011100010010000000100011;
ROM[11474] <= 32'b00000000010000010000000100010011;
ROM[11475] <= 32'b00000000000000001011001110110111;
ROM[11476] <= 32'b00111001100000111000001110010011;
ROM[11477] <= 32'b00000000111000111000001110110011;
ROM[11478] <= 32'b00000000011100010010000000100011;
ROM[11479] <= 32'b00000000010000010000000100010011;
ROM[11480] <= 32'b00000000001100010010000000100011;
ROM[11481] <= 32'b00000000010000010000000100010011;
ROM[11482] <= 32'b00000000010000010010000000100011;
ROM[11483] <= 32'b00000000010000010000000100010011;
ROM[11484] <= 32'b00000000010100010010000000100011;
ROM[11485] <= 32'b00000000010000010000000100010011;
ROM[11486] <= 32'b00000000011000010010000000100011;
ROM[11487] <= 32'b00000000010000010000000100010011;
ROM[11488] <= 32'b00000001010000000000001110010011;
ROM[11489] <= 32'b00000010010000111000001110010011;
ROM[11490] <= 32'b01000000011100010000001110110011;
ROM[11491] <= 32'b00000000011100000000001000110011;
ROM[11492] <= 32'b00000000001000000000000110110011;
ROM[11493] <= 32'b00001010010000000100000011101111;
ROM[11494] <= 32'b11111111110000010000000100010011;
ROM[11495] <= 32'b00000000000000010010001110000011;
ROM[11496] <= 32'b00000000011101100010000000100011;
ROM[11497] <= 32'b00000010101100000000001110010011;
ROM[11498] <= 32'b00000000011100010010000000100011;
ROM[11499] <= 32'b00000000010000010000000100010011;
ROM[11500] <= 32'b00000000000000000000001110010011;
ROM[11501] <= 32'b00000000011100010010000000100011;
ROM[11502] <= 32'b00000000010000010000000100010011;
ROM[11503] <= 32'b00000011000000000000001110010011;
ROM[11504] <= 32'b00000000011100010010000000100011;
ROM[11505] <= 32'b00000000010000010000000100010011;
ROM[11506] <= 32'b00000011000000000000001110010011;
ROM[11507] <= 32'b00000000011100010010000000100011;
ROM[11508] <= 32'b00000000010000010000000100010011;
ROM[11509] <= 32'b00001111110000000000001110010011;
ROM[11510] <= 32'b00000000011100010010000000100011;
ROM[11511] <= 32'b00000000010000010000000100010011;
ROM[11512] <= 32'b00000011000000000000001110010011;
ROM[11513] <= 32'b00000000011100010010000000100011;
ROM[11514] <= 32'b00000000010000010000000100010011;
ROM[11515] <= 32'b00000011000000000000001110010011;
ROM[11516] <= 32'b00000000011100010010000000100011;
ROM[11517] <= 32'b00000000010000010000000100010011;
ROM[11518] <= 32'b00000000000000000000001110010011;
ROM[11519] <= 32'b00000000011100010010000000100011;
ROM[11520] <= 32'b00000000010000010000000100010011;
ROM[11521] <= 32'b00000000000000000000001110010011;
ROM[11522] <= 32'b00000000011100010010000000100011;
ROM[11523] <= 32'b00000000010000010000000100010011;
ROM[11524] <= 32'b00000000000000001011001110110111;
ROM[11525] <= 32'b01000101110000111000001110010011;
ROM[11526] <= 32'b00000000111000111000001110110011;
ROM[11527] <= 32'b00000000011100010010000000100011;
ROM[11528] <= 32'b00000000010000010000000100010011;
ROM[11529] <= 32'b00000000001100010010000000100011;
ROM[11530] <= 32'b00000000010000010000000100010011;
ROM[11531] <= 32'b00000000010000010010000000100011;
ROM[11532] <= 32'b00000000010000010000000100010011;
ROM[11533] <= 32'b00000000010100010010000000100011;
ROM[11534] <= 32'b00000000010000010000000100010011;
ROM[11535] <= 32'b00000000011000010010000000100011;
ROM[11536] <= 32'b00000000010000010000000100010011;
ROM[11537] <= 32'b00000001010000000000001110010011;
ROM[11538] <= 32'b00000010010000111000001110010011;
ROM[11539] <= 32'b01000000011100010000001110110011;
ROM[11540] <= 32'b00000000011100000000001000110011;
ROM[11541] <= 32'b00000000001000000000000110110011;
ROM[11542] <= 32'b01111110000100000011000011101111;
ROM[11543] <= 32'b11111111110000010000000100010011;
ROM[11544] <= 32'b00000000000000010010001110000011;
ROM[11545] <= 32'b00000000011101100010000000100011;
ROM[11546] <= 32'b00000010110000000000001110010011;
ROM[11547] <= 32'b00000000011100010010000000100011;
ROM[11548] <= 32'b00000000010000010000000100010011;
ROM[11549] <= 32'b00000000000000000000001110010011;
ROM[11550] <= 32'b00000000011100010010000000100011;
ROM[11551] <= 32'b00000000010000010000000100010011;
ROM[11552] <= 32'b00000000000000000000001110010011;
ROM[11553] <= 32'b00000000011100010010000000100011;
ROM[11554] <= 32'b00000000010000010000000100010011;
ROM[11555] <= 32'b00000000000000000000001110010011;
ROM[11556] <= 32'b00000000011100010010000000100011;
ROM[11557] <= 32'b00000000010000010000000100010011;
ROM[11558] <= 32'b00000000000000000000001110010011;
ROM[11559] <= 32'b00000000011100010010000000100011;
ROM[11560] <= 32'b00000000010000010000000100010011;
ROM[11561] <= 32'b00000000000000000000001110010011;
ROM[11562] <= 32'b00000000011100010010000000100011;
ROM[11563] <= 32'b00000000010000010000000100010011;
ROM[11564] <= 32'b00000011000000000000001110010011;
ROM[11565] <= 32'b00000000011100010010000000100011;
ROM[11566] <= 32'b00000000010000010000000100010011;
ROM[11567] <= 32'b00000011000000000000001110010011;
ROM[11568] <= 32'b00000000011100010010000000100011;
ROM[11569] <= 32'b00000000010000010000000100010011;
ROM[11570] <= 32'b00000110000000000000001110010011;
ROM[11571] <= 32'b00000000011100010010000000100011;
ROM[11572] <= 32'b00000000010000010000000100010011;
ROM[11573] <= 32'b00000000000000001011001110110111;
ROM[11574] <= 32'b01010010000000111000001110010011;
ROM[11575] <= 32'b00000000111000111000001110110011;
ROM[11576] <= 32'b00000000011100010010000000100011;
ROM[11577] <= 32'b00000000010000010000000100010011;
ROM[11578] <= 32'b00000000001100010010000000100011;
ROM[11579] <= 32'b00000000010000010000000100010011;
ROM[11580] <= 32'b00000000010000010010000000100011;
ROM[11581] <= 32'b00000000010000010000000100010011;
ROM[11582] <= 32'b00000000010100010010000000100011;
ROM[11583] <= 32'b00000000010000010000000100010011;
ROM[11584] <= 32'b00000000011000010010000000100011;
ROM[11585] <= 32'b00000000010000010000000100010011;
ROM[11586] <= 32'b00000001010000000000001110010011;
ROM[11587] <= 32'b00000010010000111000001110010011;
ROM[11588] <= 32'b01000000011100010000001110110011;
ROM[11589] <= 32'b00000000011100000000001000110011;
ROM[11590] <= 32'b00000000001000000000000110110011;
ROM[11591] <= 32'b01110001110100000011000011101111;
ROM[11592] <= 32'b11111111110000010000000100010011;
ROM[11593] <= 32'b00000000000000010010001110000011;
ROM[11594] <= 32'b00000000011101100010000000100011;
ROM[11595] <= 32'b00000010110100000000001110010011;
ROM[11596] <= 32'b00000000011100010010000000100011;
ROM[11597] <= 32'b00000000010000010000000100010011;
ROM[11598] <= 32'b00000000000000000000001110010011;
ROM[11599] <= 32'b00000000011100010010000000100011;
ROM[11600] <= 32'b00000000010000010000000100010011;
ROM[11601] <= 32'b00000000000000000000001110010011;
ROM[11602] <= 32'b00000000011100010010000000100011;
ROM[11603] <= 32'b00000000010000010000000100010011;
ROM[11604] <= 32'b00000000000000000000001110010011;
ROM[11605] <= 32'b00000000011100010010000000100011;
ROM[11606] <= 32'b00000000010000010000000100010011;
ROM[11607] <= 32'b00001111110000000000001110010011;
ROM[11608] <= 32'b00000000011100010010000000100011;
ROM[11609] <= 32'b00000000010000010000000100010011;
ROM[11610] <= 32'b00000000000000000000001110010011;
ROM[11611] <= 32'b00000000011100010010000000100011;
ROM[11612] <= 32'b00000000010000010000000100010011;
ROM[11613] <= 32'b00000000000000000000001110010011;
ROM[11614] <= 32'b00000000011100010010000000100011;
ROM[11615] <= 32'b00000000010000010000000100010011;
ROM[11616] <= 32'b00000000000000000000001110010011;
ROM[11617] <= 32'b00000000011100010010000000100011;
ROM[11618] <= 32'b00000000010000010000000100010011;
ROM[11619] <= 32'b00000000000000000000001110010011;
ROM[11620] <= 32'b00000000011100010010000000100011;
ROM[11621] <= 32'b00000000010000010000000100010011;
ROM[11622] <= 32'b00000000000000001011001110110111;
ROM[11623] <= 32'b01011110010000111000001110010011;
ROM[11624] <= 32'b00000000111000111000001110110011;
ROM[11625] <= 32'b00000000011100010010000000100011;
ROM[11626] <= 32'b00000000010000010000000100010011;
ROM[11627] <= 32'b00000000001100010010000000100011;
ROM[11628] <= 32'b00000000010000010000000100010011;
ROM[11629] <= 32'b00000000010000010010000000100011;
ROM[11630] <= 32'b00000000010000010000000100010011;
ROM[11631] <= 32'b00000000010100010010000000100011;
ROM[11632] <= 32'b00000000010000010000000100010011;
ROM[11633] <= 32'b00000000011000010010000000100011;
ROM[11634] <= 32'b00000000010000010000000100010011;
ROM[11635] <= 32'b00000001010000000000001110010011;
ROM[11636] <= 32'b00000010010000111000001110010011;
ROM[11637] <= 32'b01000000011100010000001110110011;
ROM[11638] <= 32'b00000000011100000000001000110011;
ROM[11639] <= 32'b00000000001000000000000110110011;
ROM[11640] <= 32'b01100101100100000011000011101111;
ROM[11641] <= 32'b11111111110000010000000100010011;
ROM[11642] <= 32'b00000000000000010010001110000011;
ROM[11643] <= 32'b00000000011101100010000000100011;
ROM[11644] <= 32'b00000010111000000000001110010011;
ROM[11645] <= 32'b00000000011100010010000000100011;
ROM[11646] <= 32'b00000000010000010000000100010011;
ROM[11647] <= 32'b00000000000000000000001110010011;
ROM[11648] <= 32'b00000000011100010010000000100011;
ROM[11649] <= 32'b00000000010000010000000100010011;
ROM[11650] <= 32'b00000000000000000000001110010011;
ROM[11651] <= 32'b00000000011100010010000000100011;
ROM[11652] <= 32'b00000000010000010000000100010011;
ROM[11653] <= 32'b00000000000000000000001110010011;
ROM[11654] <= 32'b00000000011100010010000000100011;
ROM[11655] <= 32'b00000000010000010000000100010011;
ROM[11656] <= 32'b00000000000000000000001110010011;
ROM[11657] <= 32'b00000000011100010010000000100011;
ROM[11658] <= 32'b00000000010000010000000100010011;
ROM[11659] <= 32'b00000000000000000000001110010011;
ROM[11660] <= 32'b00000000011100010010000000100011;
ROM[11661] <= 32'b00000000010000010000000100010011;
ROM[11662] <= 32'b00000011000000000000001110010011;
ROM[11663] <= 32'b00000000011100010010000000100011;
ROM[11664] <= 32'b00000000010000010000000100010011;
ROM[11665] <= 32'b00000011000000000000001110010011;
ROM[11666] <= 32'b00000000011100010010000000100011;
ROM[11667] <= 32'b00000000010000010000000100010011;
ROM[11668] <= 32'b00000000000000000000001110010011;
ROM[11669] <= 32'b00000000011100010010000000100011;
ROM[11670] <= 32'b00000000010000010000000100010011;
ROM[11671] <= 32'b00000000000000001011001110110111;
ROM[11672] <= 32'b01101010100000111000001110010011;
ROM[11673] <= 32'b00000000111000111000001110110011;
ROM[11674] <= 32'b00000000011100010010000000100011;
ROM[11675] <= 32'b00000000010000010000000100010011;
ROM[11676] <= 32'b00000000001100010010000000100011;
ROM[11677] <= 32'b00000000010000010000000100010011;
ROM[11678] <= 32'b00000000010000010010000000100011;
ROM[11679] <= 32'b00000000010000010000000100010011;
ROM[11680] <= 32'b00000000010100010010000000100011;
ROM[11681] <= 32'b00000000010000010000000100010011;
ROM[11682] <= 32'b00000000011000010010000000100011;
ROM[11683] <= 32'b00000000010000010000000100010011;
ROM[11684] <= 32'b00000001010000000000001110010011;
ROM[11685] <= 32'b00000010010000111000001110010011;
ROM[11686] <= 32'b01000000011100010000001110110011;
ROM[11687] <= 32'b00000000011100000000001000110011;
ROM[11688] <= 32'b00000000001000000000000110110011;
ROM[11689] <= 32'b01011001010100000011000011101111;
ROM[11690] <= 32'b11111111110000010000000100010011;
ROM[11691] <= 32'b00000000000000010010001110000011;
ROM[11692] <= 32'b00000000011101100010000000100011;
ROM[11693] <= 32'b00000010111100000000001110010011;
ROM[11694] <= 32'b00000000011100010010000000100011;
ROM[11695] <= 32'b00000000010000010000000100010011;
ROM[11696] <= 32'b00000000011000000000001110010011;
ROM[11697] <= 32'b00000000011100010010000000100011;
ROM[11698] <= 32'b00000000010000010000000100010011;
ROM[11699] <= 32'b00000000110000000000001110010011;
ROM[11700] <= 32'b00000000011100010010000000100011;
ROM[11701] <= 32'b00000000010000010000000100010011;
ROM[11702] <= 32'b00000001100000000000001110010011;
ROM[11703] <= 32'b00000000011100010010000000100011;
ROM[11704] <= 32'b00000000010000010000000100010011;
ROM[11705] <= 32'b00000011000000000000001110010011;
ROM[11706] <= 32'b00000000011100010010000000100011;
ROM[11707] <= 32'b00000000010000010000000100010011;
ROM[11708] <= 32'b00000110000000000000001110010011;
ROM[11709] <= 32'b00000000011100010010000000100011;
ROM[11710] <= 32'b00000000010000010000000100010011;
ROM[11711] <= 32'b00001100000000000000001110010011;
ROM[11712] <= 32'b00000000011100010010000000100011;
ROM[11713] <= 32'b00000000010000010000000100010011;
ROM[11714] <= 32'b00001000000000000000001110010011;
ROM[11715] <= 32'b00000000011100010010000000100011;
ROM[11716] <= 32'b00000000010000010000000100010011;
ROM[11717] <= 32'b00000000000000000000001110010011;
ROM[11718] <= 32'b00000000011100010010000000100011;
ROM[11719] <= 32'b00000000010000010000000100010011;
ROM[11720] <= 32'b00000000000000001011001110110111;
ROM[11721] <= 32'b01110110110000111000001110010011;
ROM[11722] <= 32'b00000000111000111000001110110011;
ROM[11723] <= 32'b00000000011100010010000000100011;
ROM[11724] <= 32'b00000000010000010000000100010011;
ROM[11725] <= 32'b00000000001100010010000000100011;
ROM[11726] <= 32'b00000000010000010000000100010011;
ROM[11727] <= 32'b00000000010000010010000000100011;
ROM[11728] <= 32'b00000000010000010000000100010011;
ROM[11729] <= 32'b00000000010100010010000000100011;
ROM[11730] <= 32'b00000000010000010000000100010011;
ROM[11731] <= 32'b00000000011000010010000000100011;
ROM[11732] <= 32'b00000000010000010000000100010011;
ROM[11733] <= 32'b00000001010000000000001110010011;
ROM[11734] <= 32'b00000010010000111000001110010011;
ROM[11735] <= 32'b01000000011100010000001110110011;
ROM[11736] <= 32'b00000000011100000000001000110011;
ROM[11737] <= 32'b00000000001000000000000110110011;
ROM[11738] <= 32'b01001101000100000011000011101111;
ROM[11739] <= 32'b11111111110000010000000100010011;
ROM[11740] <= 32'b00000000000000010010001110000011;
ROM[11741] <= 32'b00000000011101100010000000100011;
ROM[11742] <= 32'b00000011000000000000001110010011;
ROM[11743] <= 32'b00000000011100010010000000100011;
ROM[11744] <= 32'b00000000010000010000000100010011;
ROM[11745] <= 32'b00000111110000000000001110010011;
ROM[11746] <= 32'b00000000011100010010000000100011;
ROM[11747] <= 32'b00000000010000010000000100010011;
ROM[11748] <= 32'b00001100011000000000001110010011;
ROM[11749] <= 32'b00000000011100010010000000100011;
ROM[11750] <= 32'b00000000010000010000000100010011;
ROM[11751] <= 32'b00001100111000000000001110010011;
ROM[11752] <= 32'b00000000011100010010000000100011;
ROM[11753] <= 32'b00000000010000010000000100010011;
ROM[11754] <= 32'b00001101111000000000001110010011;
ROM[11755] <= 32'b00000000011100010010000000100011;
ROM[11756] <= 32'b00000000010000010000000100010011;
ROM[11757] <= 32'b00001111011000000000001110010011;
ROM[11758] <= 32'b00000000011100010010000000100011;
ROM[11759] <= 32'b00000000010000010000000100010011;
ROM[11760] <= 32'b00001110011000000000001110010011;
ROM[11761] <= 32'b00000000011100010010000000100011;
ROM[11762] <= 32'b00000000010000010000000100010011;
ROM[11763] <= 32'b00000111110000000000001110010011;
ROM[11764] <= 32'b00000000011100010010000000100011;
ROM[11765] <= 32'b00000000010000010000000100010011;
ROM[11766] <= 32'b00000000000000000000001110010011;
ROM[11767] <= 32'b00000000011100010010000000100011;
ROM[11768] <= 32'b00000000010000010000000100010011;
ROM[11769] <= 32'b00000000000000001100001110110111;
ROM[11770] <= 32'b10000011000000111000001110010011;
ROM[11771] <= 32'b00000000111000111000001110110011;
ROM[11772] <= 32'b00000000011100010010000000100011;
ROM[11773] <= 32'b00000000010000010000000100010011;
ROM[11774] <= 32'b00000000001100010010000000100011;
ROM[11775] <= 32'b00000000010000010000000100010011;
ROM[11776] <= 32'b00000000010000010010000000100011;
ROM[11777] <= 32'b00000000010000010000000100010011;
ROM[11778] <= 32'b00000000010100010010000000100011;
ROM[11779] <= 32'b00000000010000010000000100010011;
ROM[11780] <= 32'b00000000011000010010000000100011;
ROM[11781] <= 32'b00000000010000010000000100010011;
ROM[11782] <= 32'b00000001010000000000001110010011;
ROM[11783] <= 32'b00000010010000111000001110010011;
ROM[11784] <= 32'b01000000011100010000001110110011;
ROM[11785] <= 32'b00000000011100000000001000110011;
ROM[11786] <= 32'b00000000001000000000000110110011;
ROM[11787] <= 32'b01000000110100000011000011101111;
ROM[11788] <= 32'b11111111110000010000000100010011;
ROM[11789] <= 32'b00000000000000010010001110000011;
ROM[11790] <= 32'b00000000011101100010000000100011;
ROM[11791] <= 32'b00000011000100000000001110010011;
ROM[11792] <= 32'b00000000011100010010000000100011;
ROM[11793] <= 32'b00000000010000010000000100010011;
ROM[11794] <= 32'b00000011000000000000001110010011;
ROM[11795] <= 32'b00000000011100010010000000100011;
ROM[11796] <= 32'b00000000010000010000000100010011;
ROM[11797] <= 32'b00000111000000000000001110010011;
ROM[11798] <= 32'b00000000011100010010000000100011;
ROM[11799] <= 32'b00000000010000010000000100010011;
ROM[11800] <= 32'b00000011000000000000001110010011;
ROM[11801] <= 32'b00000000011100010010000000100011;
ROM[11802] <= 32'b00000000010000010000000100010011;
ROM[11803] <= 32'b00000011000000000000001110010011;
ROM[11804] <= 32'b00000000011100010010000000100011;
ROM[11805] <= 32'b00000000010000010000000100010011;
ROM[11806] <= 32'b00000011000000000000001110010011;
ROM[11807] <= 32'b00000000011100010010000000100011;
ROM[11808] <= 32'b00000000010000010000000100010011;
ROM[11809] <= 32'b00000011000000000000001110010011;
ROM[11810] <= 32'b00000000011100010010000000100011;
ROM[11811] <= 32'b00000000010000010000000100010011;
ROM[11812] <= 32'b00001111110000000000001110010011;
ROM[11813] <= 32'b00000000011100010010000000100011;
ROM[11814] <= 32'b00000000010000010000000100010011;
ROM[11815] <= 32'b00000000000000000000001110010011;
ROM[11816] <= 32'b00000000011100010010000000100011;
ROM[11817] <= 32'b00000000010000010000000100010011;
ROM[11818] <= 32'b00000000000000001100001110110111;
ROM[11819] <= 32'b10001111010000111000001110010011;
ROM[11820] <= 32'b00000000111000111000001110110011;
ROM[11821] <= 32'b00000000011100010010000000100011;
ROM[11822] <= 32'b00000000010000010000000100010011;
ROM[11823] <= 32'b00000000001100010010000000100011;
ROM[11824] <= 32'b00000000010000010000000100010011;
ROM[11825] <= 32'b00000000010000010010000000100011;
ROM[11826] <= 32'b00000000010000010000000100010011;
ROM[11827] <= 32'b00000000010100010010000000100011;
ROM[11828] <= 32'b00000000010000010000000100010011;
ROM[11829] <= 32'b00000000011000010010000000100011;
ROM[11830] <= 32'b00000000010000010000000100010011;
ROM[11831] <= 32'b00000001010000000000001110010011;
ROM[11832] <= 32'b00000010010000111000001110010011;
ROM[11833] <= 32'b01000000011100010000001110110011;
ROM[11834] <= 32'b00000000011100000000001000110011;
ROM[11835] <= 32'b00000000001000000000000110110011;
ROM[11836] <= 32'b00110100100100000011000011101111;
ROM[11837] <= 32'b11111111110000010000000100010011;
ROM[11838] <= 32'b00000000000000010010001110000011;
ROM[11839] <= 32'b00000000011101100010000000100011;
ROM[11840] <= 32'b00000011001000000000001110010011;
ROM[11841] <= 32'b00000000011100010010000000100011;
ROM[11842] <= 32'b00000000010000010000000100010011;
ROM[11843] <= 32'b00000111100000000000001110010011;
ROM[11844] <= 32'b00000000011100010010000000100011;
ROM[11845] <= 32'b00000000010000010000000100010011;
ROM[11846] <= 32'b00001100110000000000001110010011;
ROM[11847] <= 32'b00000000011100010010000000100011;
ROM[11848] <= 32'b00000000010000010000000100010011;
ROM[11849] <= 32'b00000000110000000000001110010011;
ROM[11850] <= 32'b00000000011100010010000000100011;
ROM[11851] <= 32'b00000000010000010000000100010011;
ROM[11852] <= 32'b00000011100000000000001110010011;
ROM[11853] <= 32'b00000000011100010010000000100011;
ROM[11854] <= 32'b00000000010000010000000100010011;
ROM[11855] <= 32'b00000110000000000000001110010011;
ROM[11856] <= 32'b00000000011100010010000000100011;
ROM[11857] <= 32'b00000000010000010000000100010011;
ROM[11858] <= 32'b00001100110000000000001110010011;
ROM[11859] <= 32'b00000000011100010010000000100011;
ROM[11860] <= 32'b00000000010000010000000100010011;
ROM[11861] <= 32'b00001111110000000000001110010011;
ROM[11862] <= 32'b00000000011100010010000000100011;
ROM[11863] <= 32'b00000000010000010000000100010011;
ROM[11864] <= 32'b00000000000000000000001110010011;
ROM[11865] <= 32'b00000000011100010010000000100011;
ROM[11866] <= 32'b00000000010000010000000100010011;
ROM[11867] <= 32'b00000000000000001100001110110111;
ROM[11868] <= 32'b10011011100000111000001110010011;
ROM[11869] <= 32'b00000000111000111000001110110011;
ROM[11870] <= 32'b00000000011100010010000000100011;
ROM[11871] <= 32'b00000000010000010000000100010011;
ROM[11872] <= 32'b00000000001100010010000000100011;
ROM[11873] <= 32'b00000000010000010000000100010011;
ROM[11874] <= 32'b00000000010000010010000000100011;
ROM[11875] <= 32'b00000000010000010000000100010011;
ROM[11876] <= 32'b00000000010100010010000000100011;
ROM[11877] <= 32'b00000000010000010000000100010011;
ROM[11878] <= 32'b00000000011000010010000000100011;
ROM[11879] <= 32'b00000000010000010000000100010011;
ROM[11880] <= 32'b00000001010000000000001110010011;
ROM[11881] <= 32'b00000010010000111000001110010011;
ROM[11882] <= 32'b01000000011100010000001110110011;
ROM[11883] <= 32'b00000000011100000000001000110011;
ROM[11884] <= 32'b00000000001000000000000110110011;
ROM[11885] <= 32'b00101000010100000011000011101111;
ROM[11886] <= 32'b11111111110000010000000100010011;
ROM[11887] <= 32'b00000000000000010010001110000011;
ROM[11888] <= 32'b00000000011101100010000000100011;
ROM[11889] <= 32'b00000011001100000000001110010011;
ROM[11890] <= 32'b00000000011100010010000000100011;
ROM[11891] <= 32'b00000000010000010000000100010011;
ROM[11892] <= 32'b00000111100000000000001110010011;
ROM[11893] <= 32'b00000000011100010010000000100011;
ROM[11894] <= 32'b00000000010000010000000100010011;
ROM[11895] <= 32'b00001100110000000000001110010011;
ROM[11896] <= 32'b00000000011100010010000000100011;
ROM[11897] <= 32'b00000000010000010000000100010011;
ROM[11898] <= 32'b00000000110000000000001110010011;
ROM[11899] <= 32'b00000000011100010010000000100011;
ROM[11900] <= 32'b00000000010000010000000100010011;
ROM[11901] <= 32'b00000011100000000000001110010011;
ROM[11902] <= 32'b00000000011100010010000000100011;
ROM[11903] <= 32'b00000000010000010000000100010011;
ROM[11904] <= 32'b00000000110000000000001110010011;
ROM[11905] <= 32'b00000000011100010010000000100011;
ROM[11906] <= 32'b00000000010000010000000100010011;
ROM[11907] <= 32'b00001100110000000000001110010011;
ROM[11908] <= 32'b00000000011100010010000000100011;
ROM[11909] <= 32'b00000000010000010000000100010011;
ROM[11910] <= 32'b00000111100000000000001110010011;
ROM[11911] <= 32'b00000000011100010010000000100011;
ROM[11912] <= 32'b00000000010000010000000100010011;
ROM[11913] <= 32'b00000000000000000000001110010011;
ROM[11914] <= 32'b00000000011100010010000000100011;
ROM[11915] <= 32'b00000000010000010000000100010011;
ROM[11916] <= 32'b00000000000000001100001110110111;
ROM[11917] <= 32'b10100111110000111000001110010011;
ROM[11918] <= 32'b00000000111000111000001110110011;
ROM[11919] <= 32'b00000000011100010010000000100011;
ROM[11920] <= 32'b00000000010000010000000100010011;
ROM[11921] <= 32'b00000000001100010010000000100011;
ROM[11922] <= 32'b00000000010000010000000100010011;
ROM[11923] <= 32'b00000000010000010010000000100011;
ROM[11924] <= 32'b00000000010000010000000100010011;
ROM[11925] <= 32'b00000000010100010010000000100011;
ROM[11926] <= 32'b00000000010000010000000100010011;
ROM[11927] <= 32'b00000000011000010010000000100011;
ROM[11928] <= 32'b00000000010000010000000100010011;
ROM[11929] <= 32'b00000001010000000000001110010011;
ROM[11930] <= 32'b00000010010000111000001110010011;
ROM[11931] <= 32'b01000000011100010000001110110011;
ROM[11932] <= 32'b00000000011100000000001000110011;
ROM[11933] <= 32'b00000000001000000000000110110011;
ROM[11934] <= 32'b00011100000100000011000011101111;
ROM[11935] <= 32'b11111111110000010000000100010011;
ROM[11936] <= 32'b00000000000000010010001110000011;
ROM[11937] <= 32'b00000000011101100010000000100011;
ROM[11938] <= 32'b00000011010000000000001110010011;
ROM[11939] <= 32'b00000000011100010010000000100011;
ROM[11940] <= 32'b00000000010000010000000100010011;
ROM[11941] <= 32'b00000001110000000000001110010011;
ROM[11942] <= 32'b00000000011100010010000000100011;
ROM[11943] <= 32'b00000000010000010000000100010011;
ROM[11944] <= 32'b00000011110000000000001110010011;
ROM[11945] <= 32'b00000000011100010010000000100011;
ROM[11946] <= 32'b00000000010000010000000100010011;
ROM[11947] <= 32'b00000110110000000000001110010011;
ROM[11948] <= 32'b00000000011100010010000000100011;
ROM[11949] <= 32'b00000000010000010000000100010011;
ROM[11950] <= 32'b00001100110000000000001110010011;
ROM[11951] <= 32'b00000000011100010010000000100011;
ROM[11952] <= 32'b00000000010000010000000100010011;
ROM[11953] <= 32'b00001111111000000000001110010011;
ROM[11954] <= 32'b00000000011100010010000000100011;
ROM[11955] <= 32'b00000000010000010000000100010011;
ROM[11956] <= 32'b00000000110000000000001110010011;
ROM[11957] <= 32'b00000000011100010010000000100011;
ROM[11958] <= 32'b00000000010000010000000100010011;
ROM[11959] <= 32'b00000001111000000000001110010011;
ROM[11960] <= 32'b00000000011100010010000000100011;
ROM[11961] <= 32'b00000000010000010000000100010011;
ROM[11962] <= 32'b00000000000000000000001110010011;
ROM[11963] <= 32'b00000000011100010010000000100011;
ROM[11964] <= 32'b00000000010000010000000100010011;
ROM[11965] <= 32'b00000000000000001100001110110111;
ROM[11966] <= 32'b10110100000000111000001110010011;
ROM[11967] <= 32'b00000000111000111000001110110011;
ROM[11968] <= 32'b00000000011100010010000000100011;
ROM[11969] <= 32'b00000000010000010000000100010011;
ROM[11970] <= 32'b00000000001100010010000000100011;
ROM[11971] <= 32'b00000000010000010000000100010011;
ROM[11972] <= 32'b00000000010000010010000000100011;
ROM[11973] <= 32'b00000000010000010000000100010011;
ROM[11974] <= 32'b00000000010100010010000000100011;
ROM[11975] <= 32'b00000000010000010000000100010011;
ROM[11976] <= 32'b00000000011000010010000000100011;
ROM[11977] <= 32'b00000000010000010000000100010011;
ROM[11978] <= 32'b00000001010000000000001110010011;
ROM[11979] <= 32'b00000010010000111000001110010011;
ROM[11980] <= 32'b01000000011100010000001110110011;
ROM[11981] <= 32'b00000000011100000000001000110011;
ROM[11982] <= 32'b00000000001000000000000110110011;
ROM[11983] <= 32'b00001111110100000011000011101111;
ROM[11984] <= 32'b11111111110000010000000100010011;
ROM[11985] <= 32'b00000000000000010010001110000011;
ROM[11986] <= 32'b00000000011101100010000000100011;
ROM[11987] <= 32'b00000011010100000000001110010011;
ROM[11988] <= 32'b00000000011100010010000000100011;
ROM[11989] <= 32'b00000000010000010000000100010011;
ROM[11990] <= 32'b00001111110000000000001110010011;
ROM[11991] <= 32'b00000000011100010010000000100011;
ROM[11992] <= 32'b00000000010000010000000100010011;
ROM[11993] <= 32'b00001100000000000000001110010011;
ROM[11994] <= 32'b00000000011100010010000000100011;
ROM[11995] <= 32'b00000000010000010000000100010011;
ROM[11996] <= 32'b00001111100000000000001110010011;
ROM[11997] <= 32'b00000000011100010010000000100011;
ROM[11998] <= 32'b00000000010000010000000100010011;
ROM[11999] <= 32'b00000000110000000000001110010011;
ROM[12000] <= 32'b00000000011100010010000000100011;
ROM[12001] <= 32'b00000000010000010000000100010011;
ROM[12002] <= 32'b00000000110000000000001110010011;
ROM[12003] <= 32'b00000000011100010010000000100011;
ROM[12004] <= 32'b00000000010000010000000100010011;
ROM[12005] <= 32'b00001100110000000000001110010011;
ROM[12006] <= 32'b00000000011100010010000000100011;
ROM[12007] <= 32'b00000000010000010000000100010011;
ROM[12008] <= 32'b00000111100000000000001110010011;
ROM[12009] <= 32'b00000000011100010010000000100011;
ROM[12010] <= 32'b00000000010000010000000100010011;
ROM[12011] <= 32'b00000000000000000000001110010011;
ROM[12012] <= 32'b00000000011100010010000000100011;
ROM[12013] <= 32'b00000000010000010000000100010011;
ROM[12014] <= 32'b00000000000000001100001110110111;
ROM[12015] <= 32'b11000000010000111000001110010011;
ROM[12016] <= 32'b00000000111000111000001110110011;
ROM[12017] <= 32'b00000000011100010010000000100011;
ROM[12018] <= 32'b00000000010000010000000100010011;
ROM[12019] <= 32'b00000000001100010010000000100011;
ROM[12020] <= 32'b00000000010000010000000100010011;
ROM[12021] <= 32'b00000000010000010010000000100011;
ROM[12022] <= 32'b00000000010000010000000100010011;
ROM[12023] <= 32'b00000000010100010010000000100011;
ROM[12024] <= 32'b00000000010000010000000100010011;
ROM[12025] <= 32'b00000000011000010010000000100011;
ROM[12026] <= 32'b00000000010000010000000100010011;
ROM[12027] <= 32'b00000001010000000000001110010011;
ROM[12028] <= 32'b00000010010000111000001110010011;
ROM[12029] <= 32'b01000000011100010000001110110011;
ROM[12030] <= 32'b00000000011100000000001000110011;
ROM[12031] <= 32'b00000000001000000000000110110011;
ROM[12032] <= 32'b00000011100100000011000011101111;
ROM[12033] <= 32'b11111111110000010000000100010011;
ROM[12034] <= 32'b00000000000000010010001110000011;
ROM[12035] <= 32'b00000000011101100010000000100011;
ROM[12036] <= 32'b00000011011000000000001110010011;
ROM[12037] <= 32'b00000000011100010010000000100011;
ROM[12038] <= 32'b00000000010000010000000100010011;
ROM[12039] <= 32'b00000011100000000000001110010011;
ROM[12040] <= 32'b00000000011100010010000000100011;
ROM[12041] <= 32'b00000000010000010000000100010011;
ROM[12042] <= 32'b00000110000000000000001110010011;
ROM[12043] <= 32'b00000000011100010010000000100011;
ROM[12044] <= 32'b00000000010000010000000100010011;
ROM[12045] <= 32'b00001100000000000000001110010011;
ROM[12046] <= 32'b00000000011100010010000000100011;
ROM[12047] <= 32'b00000000010000010000000100010011;
ROM[12048] <= 32'b00001111100000000000001110010011;
ROM[12049] <= 32'b00000000011100010010000000100011;
ROM[12050] <= 32'b00000000010000010000000100010011;
ROM[12051] <= 32'b00001100110000000000001110010011;
ROM[12052] <= 32'b00000000011100010010000000100011;
ROM[12053] <= 32'b00000000010000010000000100010011;
ROM[12054] <= 32'b00001100110000000000001110010011;
ROM[12055] <= 32'b00000000011100010010000000100011;
ROM[12056] <= 32'b00000000010000010000000100010011;
ROM[12057] <= 32'b00000111100000000000001110010011;
ROM[12058] <= 32'b00000000011100010010000000100011;
ROM[12059] <= 32'b00000000010000010000000100010011;
ROM[12060] <= 32'b00000000000000000000001110010011;
ROM[12061] <= 32'b00000000011100010010000000100011;
ROM[12062] <= 32'b00000000010000010000000100010011;
ROM[12063] <= 32'b00000000000000001100001110110111;
ROM[12064] <= 32'b11001100100000111000001110010011;
ROM[12065] <= 32'b00000000111000111000001110110011;
ROM[12066] <= 32'b00000000011100010010000000100011;
ROM[12067] <= 32'b00000000010000010000000100010011;
ROM[12068] <= 32'b00000000001100010010000000100011;
ROM[12069] <= 32'b00000000010000010000000100010011;
ROM[12070] <= 32'b00000000010000010010000000100011;
ROM[12071] <= 32'b00000000010000010000000100010011;
ROM[12072] <= 32'b00000000010100010010000000100011;
ROM[12073] <= 32'b00000000010000010000000100010011;
ROM[12074] <= 32'b00000000011000010010000000100011;
ROM[12075] <= 32'b00000000010000010000000100010011;
ROM[12076] <= 32'b00000001010000000000001110010011;
ROM[12077] <= 32'b00000010010000111000001110010011;
ROM[12078] <= 32'b01000000011100010000001110110011;
ROM[12079] <= 32'b00000000011100000000001000110011;
ROM[12080] <= 32'b00000000001000000000000110110011;
ROM[12081] <= 32'b01110111010000000011000011101111;
ROM[12082] <= 32'b11111111110000010000000100010011;
ROM[12083] <= 32'b00000000000000010010001110000011;
ROM[12084] <= 32'b00000000011101100010000000100011;
ROM[12085] <= 32'b00000011011100000000001110010011;
ROM[12086] <= 32'b00000000011100010010000000100011;
ROM[12087] <= 32'b00000000010000010000000100010011;
ROM[12088] <= 32'b00001111110000000000001110010011;
ROM[12089] <= 32'b00000000011100010010000000100011;
ROM[12090] <= 32'b00000000010000010000000100010011;
ROM[12091] <= 32'b00001100110000000000001110010011;
ROM[12092] <= 32'b00000000011100010010000000100011;
ROM[12093] <= 32'b00000000010000010000000100010011;
ROM[12094] <= 32'b00000000110000000000001110010011;
ROM[12095] <= 32'b00000000011100010010000000100011;
ROM[12096] <= 32'b00000000010000010000000100010011;
ROM[12097] <= 32'b00000001100000000000001110010011;
ROM[12098] <= 32'b00000000011100010010000000100011;
ROM[12099] <= 32'b00000000010000010000000100010011;
ROM[12100] <= 32'b00000011000000000000001110010011;
ROM[12101] <= 32'b00000000011100010010000000100011;
ROM[12102] <= 32'b00000000010000010000000100010011;
ROM[12103] <= 32'b00000011000000000000001110010011;
ROM[12104] <= 32'b00000000011100010010000000100011;
ROM[12105] <= 32'b00000000010000010000000100010011;
ROM[12106] <= 32'b00000011000000000000001110010011;
ROM[12107] <= 32'b00000000011100010010000000100011;
ROM[12108] <= 32'b00000000010000010000000100010011;
ROM[12109] <= 32'b00000000000000000000001110010011;
ROM[12110] <= 32'b00000000011100010010000000100011;
ROM[12111] <= 32'b00000000010000010000000100010011;
ROM[12112] <= 32'b00000000000000001100001110110111;
ROM[12113] <= 32'b11011000110000111000001110010011;
ROM[12114] <= 32'b00000000111000111000001110110011;
ROM[12115] <= 32'b00000000011100010010000000100011;
ROM[12116] <= 32'b00000000010000010000000100010011;
ROM[12117] <= 32'b00000000001100010010000000100011;
ROM[12118] <= 32'b00000000010000010000000100010011;
ROM[12119] <= 32'b00000000010000010010000000100011;
ROM[12120] <= 32'b00000000010000010000000100010011;
ROM[12121] <= 32'b00000000010100010010000000100011;
ROM[12122] <= 32'b00000000010000010000000100010011;
ROM[12123] <= 32'b00000000011000010010000000100011;
ROM[12124] <= 32'b00000000010000010000000100010011;
ROM[12125] <= 32'b00000001010000000000001110010011;
ROM[12126] <= 32'b00000010010000111000001110010011;
ROM[12127] <= 32'b01000000011100010000001110110011;
ROM[12128] <= 32'b00000000011100000000001000110011;
ROM[12129] <= 32'b00000000001000000000000110110011;
ROM[12130] <= 32'b01101011000000000011000011101111;
ROM[12131] <= 32'b11111111110000010000000100010011;
ROM[12132] <= 32'b00000000000000010010001110000011;
ROM[12133] <= 32'b00000000011101100010000000100011;
ROM[12134] <= 32'b00000011100000000000001110010011;
ROM[12135] <= 32'b00000000011100010010000000100011;
ROM[12136] <= 32'b00000000010000010000000100010011;
ROM[12137] <= 32'b00000111100000000000001110010011;
ROM[12138] <= 32'b00000000011100010010000000100011;
ROM[12139] <= 32'b00000000010000010000000100010011;
ROM[12140] <= 32'b00001100110000000000001110010011;
ROM[12141] <= 32'b00000000011100010010000000100011;
ROM[12142] <= 32'b00000000010000010000000100010011;
ROM[12143] <= 32'b00001100110000000000001110010011;
ROM[12144] <= 32'b00000000011100010010000000100011;
ROM[12145] <= 32'b00000000010000010000000100010011;
ROM[12146] <= 32'b00000111100000000000001110010011;
ROM[12147] <= 32'b00000000011100010010000000100011;
ROM[12148] <= 32'b00000000010000010000000100010011;
ROM[12149] <= 32'b00001100110000000000001110010011;
ROM[12150] <= 32'b00000000011100010010000000100011;
ROM[12151] <= 32'b00000000010000010000000100010011;
ROM[12152] <= 32'b00001100110000000000001110010011;
ROM[12153] <= 32'b00000000011100010010000000100011;
ROM[12154] <= 32'b00000000010000010000000100010011;
ROM[12155] <= 32'b00000111100000000000001110010011;
ROM[12156] <= 32'b00000000011100010010000000100011;
ROM[12157] <= 32'b00000000010000010000000100010011;
ROM[12158] <= 32'b00000000000000000000001110010011;
ROM[12159] <= 32'b00000000011100010010000000100011;
ROM[12160] <= 32'b00000000010000010000000100010011;
ROM[12161] <= 32'b00000000000000001100001110110111;
ROM[12162] <= 32'b11100101000000111000001110010011;
ROM[12163] <= 32'b00000000111000111000001110110011;
ROM[12164] <= 32'b00000000011100010010000000100011;
ROM[12165] <= 32'b00000000010000010000000100010011;
ROM[12166] <= 32'b00000000001100010010000000100011;
ROM[12167] <= 32'b00000000010000010000000100010011;
ROM[12168] <= 32'b00000000010000010010000000100011;
ROM[12169] <= 32'b00000000010000010000000100010011;
ROM[12170] <= 32'b00000000010100010010000000100011;
ROM[12171] <= 32'b00000000010000010000000100010011;
ROM[12172] <= 32'b00000000011000010010000000100011;
ROM[12173] <= 32'b00000000010000010000000100010011;
ROM[12174] <= 32'b00000001010000000000001110010011;
ROM[12175] <= 32'b00000010010000111000001110010011;
ROM[12176] <= 32'b01000000011100010000001110110011;
ROM[12177] <= 32'b00000000011100000000001000110011;
ROM[12178] <= 32'b00000000001000000000000110110011;
ROM[12179] <= 32'b01011110110000000011000011101111;
ROM[12180] <= 32'b11111111110000010000000100010011;
ROM[12181] <= 32'b00000000000000010010001110000011;
ROM[12182] <= 32'b00000000011101100010000000100011;
ROM[12183] <= 32'b00000011100100000000001110010011;
ROM[12184] <= 32'b00000000011100010010000000100011;
ROM[12185] <= 32'b00000000010000010000000100010011;
ROM[12186] <= 32'b00000111100000000000001110010011;
ROM[12187] <= 32'b00000000011100010010000000100011;
ROM[12188] <= 32'b00000000010000010000000100010011;
ROM[12189] <= 32'b00001100110000000000001110010011;
ROM[12190] <= 32'b00000000011100010010000000100011;
ROM[12191] <= 32'b00000000010000010000000100010011;
ROM[12192] <= 32'b00001100110000000000001110010011;
ROM[12193] <= 32'b00000000011100010010000000100011;
ROM[12194] <= 32'b00000000010000010000000100010011;
ROM[12195] <= 32'b00000111110000000000001110010011;
ROM[12196] <= 32'b00000000011100010010000000100011;
ROM[12197] <= 32'b00000000010000010000000100010011;
ROM[12198] <= 32'b00000000110000000000001110010011;
ROM[12199] <= 32'b00000000011100010010000000100011;
ROM[12200] <= 32'b00000000010000010000000100010011;
ROM[12201] <= 32'b00000001100000000000001110010011;
ROM[12202] <= 32'b00000000011100010010000000100011;
ROM[12203] <= 32'b00000000010000010000000100010011;
ROM[12204] <= 32'b00000111000000000000001110010011;
ROM[12205] <= 32'b00000000011100010010000000100011;
ROM[12206] <= 32'b00000000010000010000000100010011;
ROM[12207] <= 32'b00000000000000000000001110010011;
ROM[12208] <= 32'b00000000011100010010000000100011;
ROM[12209] <= 32'b00000000010000010000000100010011;
ROM[12210] <= 32'b00000000000000001100001110110111;
ROM[12211] <= 32'b11110001010000111000001110010011;
ROM[12212] <= 32'b00000000111000111000001110110011;
ROM[12213] <= 32'b00000000011100010010000000100011;
ROM[12214] <= 32'b00000000010000010000000100010011;
ROM[12215] <= 32'b00000000001100010010000000100011;
ROM[12216] <= 32'b00000000010000010000000100010011;
ROM[12217] <= 32'b00000000010000010010000000100011;
ROM[12218] <= 32'b00000000010000010000000100010011;
ROM[12219] <= 32'b00000000010100010010000000100011;
ROM[12220] <= 32'b00000000010000010000000100010011;
ROM[12221] <= 32'b00000000011000010010000000100011;
ROM[12222] <= 32'b00000000010000010000000100010011;
ROM[12223] <= 32'b00000001010000000000001110010011;
ROM[12224] <= 32'b00000010010000111000001110010011;
ROM[12225] <= 32'b01000000011100010000001110110011;
ROM[12226] <= 32'b00000000011100000000001000110011;
ROM[12227] <= 32'b00000000001000000000000110110011;
ROM[12228] <= 32'b01010010100000000011000011101111;
ROM[12229] <= 32'b11111111110000010000000100010011;
ROM[12230] <= 32'b00000000000000010010001110000011;
ROM[12231] <= 32'b00000000011101100010000000100011;
ROM[12232] <= 32'b00000011101000000000001110010011;
ROM[12233] <= 32'b00000000011100010010000000100011;
ROM[12234] <= 32'b00000000010000010000000100010011;
ROM[12235] <= 32'b00000000000000000000001110010011;
ROM[12236] <= 32'b00000000011100010010000000100011;
ROM[12237] <= 32'b00000000010000010000000100010011;
ROM[12238] <= 32'b00000011000000000000001110010011;
ROM[12239] <= 32'b00000000011100010010000000100011;
ROM[12240] <= 32'b00000000010000010000000100010011;
ROM[12241] <= 32'b00000011000000000000001110010011;
ROM[12242] <= 32'b00000000011100010010000000100011;
ROM[12243] <= 32'b00000000010000010000000100010011;
ROM[12244] <= 32'b00000000000000000000001110010011;
ROM[12245] <= 32'b00000000011100010010000000100011;
ROM[12246] <= 32'b00000000010000010000000100010011;
ROM[12247] <= 32'b00000000000000000000001110010011;
ROM[12248] <= 32'b00000000011100010010000000100011;
ROM[12249] <= 32'b00000000010000010000000100010011;
ROM[12250] <= 32'b00000011000000000000001110010011;
ROM[12251] <= 32'b00000000011100010010000000100011;
ROM[12252] <= 32'b00000000010000010000000100010011;
ROM[12253] <= 32'b00000011000000000000001110010011;
ROM[12254] <= 32'b00000000011100010010000000100011;
ROM[12255] <= 32'b00000000010000010000000100010011;
ROM[12256] <= 32'b00000000000000000000001110010011;
ROM[12257] <= 32'b00000000011100010010000000100011;
ROM[12258] <= 32'b00000000010000010000000100010011;
ROM[12259] <= 32'b00000000000000001100001110110111;
ROM[12260] <= 32'b11111101100000111000001110010011;
ROM[12261] <= 32'b00000000111000111000001110110011;
ROM[12262] <= 32'b00000000011100010010000000100011;
ROM[12263] <= 32'b00000000010000010000000100010011;
ROM[12264] <= 32'b00000000001100010010000000100011;
ROM[12265] <= 32'b00000000010000010000000100010011;
ROM[12266] <= 32'b00000000010000010010000000100011;
ROM[12267] <= 32'b00000000010000010000000100010011;
ROM[12268] <= 32'b00000000010100010010000000100011;
ROM[12269] <= 32'b00000000010000010000000100010011;
ROM[12270] <= 32'b00000000011000010010000000100011;
ROM[12271] <= 32'b00000000010000010000000100010011;
ROM[12272] <= 32'b00000001010000000000001110010011;
ROM[12273] <= 32'b00000010010000111000001110010011;
ROM[12274] <= 32'b01000000011100010000001110110011;
ROM[12275] <= 32'b00000000011100000000001000110011;
ROM[12276] <= 32'b00000000001000000000000110110011;
ROM[12277] <= 32'b01000110010000000011000011101111;
ROM[12278] <= 32'b11111111110000010000000100010011;
ROM[12279] <= 32'b00000000000000010010001110000011;
ROM[12280] <= 32'b00000000011101100010000000100011;
ROM[12281] <= 32'b00000011101100000000001110010011;
ROM[12282] <= 32'b00000000011100010010000000100011;
ROM[12283] <= 32'b00000000010000010000000100010011;
ROM[12284] <= 32'b00000000000000000000001110010011;
ROM[12285] <= 32'b00000000011100010010000000100011;
ROM[12286] <= 32'b00000000010000010000000100010011;
ROM[12287] <= 32'b00000011000000000000001110010011;
ROM[12288] <= 32'b00000000011100010010000000100011;
ROM[12289] <= 32'b00000000010000010000000100010011;
ROM[12290] <= 32'b00000011000000000000001110010011;
ROM[12291] <= 32'b00000000011100010010000000100011;
ROM[12292] <= 32'b00000000010000010000000100010011;
ROM[12293] <= 32'b00000000000000000000001110010011;
ROM[12294] <= 32'b00000000011100010010000000100011;
ROM[12295] <= 32'b00000000010000010000000100010011;
ROM[12296] <= 32'b00000000000000000000001110010011;
ROM[12297] <= 32'b00000000011100010010000000100011;
ROM[12298] <= 32'b00000000010000010000000100010011;
ROM[12299] <= 32'b00000011000000000000001110010011;
ROM[12300] <= 32'b00000000011100010010000000100011;
ROM[12301] <= 32'b00000000010000010000000100010011;
ROM[12302] <= 32'b00000011000000000000001110010011;
ROM[12303] <= 32'b00000000011100010010000000100011;
ROM[12304] <= 32'b00000000010000010000000100010011;
ROM[12305] <= 32'b00000110000000000000001110010011;
ROM[12306] <= 32'b00000000011100010010000000100011;
ROM[12307] <= 32'b00000000010000010000000100010011;
ROM[12308] <= 32'b00000000000000001100001110110111;
ROM[12309] <= 32'b00001001110000111000001110010011;
ROM[12310] <= 32'b00000000111000111000001110110011;
ROM[12311] <= 32'b00000000011100010010000000100011;
ROM[12312] <= 32'b00000000010000010000000100010011;
ROM[12313] <= 32'b00000000001100010010000000100011;
ROM[12314] <= 32'b00000000010000010000000100010011;
ROM[12315] <= 32'b00000000010000010010000000100011;
ROM[12316] <= 32'b00000000010000010000000100010011;
ROM[12317] <= 32'b00000000010100010010000000100011;
ROM[12318] <= 32'b00000000010000010000000100010011;
ROM[12319] <= 32'b00000000011000010010000000100011;
ROM[12320] <= 32'b00000000010000010000000100010011;
ROM[12321] <= 32'b00000001010000000000001110010011;
ROM[12322] <= 32'b00000010010000111000001110010011;
ROM[12323] <= 32'b01000000011100010000001110110011;
ROM[12324] <= 32'b00000000011100000000001000110011;
ROM[12325] <= 32'b00000000001000000000000110110011;
ROM[12326] <= 32'b00111010000000000011000011101111;
ROM[12327] <= 32'b11111111110000010000000100010011;
ROM[12328] <= 32'b00000000000000010010001110000011;
ROM[12329] <= 32'b00000000011101100010000000100011;
ROM[12330] <= 32'b00000011110000000000001110010011;
ROM[12331] <= 32'b00000000011100010010000000100011;
ROM[12332] <= 32'b00000000010000010000000100010011;
ROM[12333] <= 32'b00000001100000000000001110010011;
ROM[12334] <= 32'b00000000011100010010000000100011;
ROM[12335] <= 32'b00000000010000010000000100010011;
ROM[12336] <= 32'b00000011000000000000001110010011;
ROM[12337] <= 32'b00000000011100010010000000100011;
ROM[12338] <= 32'b00000000010000010000000100010011;
ROM[12339] <= 32'b00000110000000000000001110010011;
ROM[12340] <= 32'b00000000011100010010000000100011;
ROM[12341] <= 32'b00000000010000010000000100010011;
ROM[12342] <= 32'b00001100000000000000001110010011;
ROM[12343] <= 32'b00000000011100010010000000100011;
ROM[12344] <= 32'b00000000010000010000000100010011;
ROM[12345] <= 32'b00000110000000000000001110010011;
ROM[12346] <= 32'b00000000011100010010000000100011;
ROM[12347] <= 32'b00000000010000010000000100010011;
ROM[12348] <= 32'b00000011000000000000001110010011;
ROM[12349] <= 32'b00000000011100010010000000100011;
ROM[12350] <= 32'b00000000010000010000000100010011;
ROM[12351] <= 32'b00000001100000000000001110010011;
ROM[12352] <= 32'b00000000011100010010000000100011;
ROM[12353] <= 32'b00000000010000010000000100010011;
ROM[12354] <= 32'b00000000000000000000001110010011;
ROM[12355] <= 32'b00000000011100010010000000100011;
ROM[12356] <= 32'b00000000010000010000000100010011;
ROM[12357] <= 32'b00000000000000001100001110110111;
ROM[12358] <= 32'b00010110000000111000001110010011;
ROM[12359] <= 32'b00000000111000111000001110110011;
ROM[12360] <= 32'b00000000011100010010000000100011;
ROM[12361] <= 32'b00000000010000010000000100010011;
ROM[12362] <= 32'b00000000001100010010000000100011;
ROM[12363] <= 32'b00000000010000010000000100010011;
ROM[12364] <= 32'b00000000010000010010000000100011;
ROM[12365] <= 32'b00000000010000010000000100010011;
ROM[12366] <= 32'b00000000010100010010000000100011;
ROM[12367] <= 32'b00000000010000010000000100010011;
ROM[12368] <= 32'b00000000011000010010000000100011;
ROM[12369] <= 32'b00000000010000010000000100010011;
ROM[12370] <= 32'b00000001010000000000001110010011;
ROM[12371] <= 32'b00000010010000111000001110010011;
ROM[12372] <= 32'b01000000011100010000001110110011;
ROM[12373] <= 32'b00000000011100000000001000110011;
ROM[12374] <= 32'b00000000001000000000000110110011;
ROM[12375] <= 32'b00101101110000000011000011101111;
ROM[12376] <= 32'b11111111110000010000000100010011;
ROM[12377] <= 32'b00000000000000010010001110000011;
ROM[12378] <= 32'b00000000011101100010000000100011;
ROM[12379] <= 32'b00000011110100000000001110010011;
ROM[12380] <= 32'b00000000011100010010000000100011;
ROM[12381] <= 32'b00000000010000010000000100010011;
ROM[12382] <= 32'b00000000000000000000001110010011;
ROM[12383] <= 32'b00000000011100010010000000100011;
ROM[12384] <= 32'b00000000010000010000000100010011;
ROM[12385] <= 32'b00000000000000000000001110010011;
ROM[12386] <= 32'b00000000011100010010000000100011;
ROM[12387] <= 32'b00000000010000010000000100010011;
ROM[12388] <= 32'b00001111110000000000001110010011;
ROM[12389] <= 32'b00000000011100010010000000100011;
ROM[12390] <= 32'b00000000010000010000000100010011;
ROM[12391] <= 32'b00000000000000000000001110010011;
ROM[12392] <= 32'b00000000011100010010000000100011;
ROM[12393] <= 32'b00000000010000010000000100010011;
ROM[12394] <= 32'b00000000000000000000001110010011;
ROM[12395] <= 32'b00000000011100010010000000100011;
ROM[12396] <= 32'b00000000010000010000000100010011;
ROM[12397] <= 32'b00001111110000000000001110010011;
ROM[12398] <= 32'b00000000011100010010000000100011;
ROM[12399] <= 32'b00000000010000010000000100010011;
ROM[12400] <= 32'b00000000000000000000001110010011;
ROM[12401] <= 32'b00000000011100010010000000100011;
ROM[12402] <= 32'b00000000010000010000000100010011;
ROM[12403] <= 32'b00000000000000000000001110010011;
ROM[12404] <= 32'b00000000011100010010000000100011;
ROM[12405] <= 32'b00000000010000010000000100010011;
ROM[12406] <= 32'b00000000000000001100001110110111;
ROM[12407] <= 32'b00100010010000111000001110010011;
ROM[12408] <= 32'b00000000111000111000001110110011;
ROM[12409] <= 32'b00000000011100010010000000100011;
ROM[12410] <= 32'b00000000010000010000000100010011;
ROM[12411] <= 32'b00000000001100010010000000100011;
ROM[12412] <= 32'b00000000010000010000000100010011;
ROM[12413] <= 32'b00000000010000010010000000100011;
ROM[12414] <= 32'b00000000010000010000000100010011;
ROM[12415] <= 32'b00000000010100010010000000100011;
ROM[12416] <= 32'b00000000010000010000000100010011;
ROM[12417] <= 32'b00000000011000010010000000100011;
ROM[12418] <= 32'b00000000010000010000000100010011;
ROM[12419] <= 32'b00000001010000000000001110010011;
ROM[12420] <= 32'b00000010010000111000001110010011;
ROM[12421] <= 32'b01000000011100010000001110110011;
ROM[12422] <= 32'b00000000011100000000001000110011;
ROM[12423] <= 32'b00000000001000000000000110110011;
ROM[12424] <= 32'b00100001100000000011000011101111;
ROM[12425] <= 32'b11111111110000010000000100010011;
ROM[12426] <= 32'b00000000000000010010001110000011;
ROM[12427] <= 32'b00000000011101100010000000100011;
ROM[12428] <= 32'b00000011111000000000001110010011;
ROM[12429] <= 32'b00000000011100010010000000100011;
ROM[12430] <= 32'b00000000010000010000000100010011;
ROM[12431] <= 32'b00000110000000000000001110010011;
ROM[12432] <= 32'b00000000011100010010000000100011;
ROM[12433] <= 32'b00000000010000010000000100010011;
ROM[12434] <= 32'b00000011000000000000001110010011;
ROM[12435] <= 32'b00000000011100010010000000100011;
ROM[12436] <= 32'b00000000010000010000000100010011;
ROM[12437] <= 32'b00000001100000000000001110010011;
ROM[12438] <= 32'b00000000011100010010000000100011;
ROM[12439] <= 32'b00000000010000010000000100010011;
ROM[12440] <= 32'b00000000110000000000001110010011;
ROM[12441] <= 32'b00000000011100010010000000100011;
ROM[12442] <= 32'b00000000010000010000000100010011;
ROM[12443] <= 32'b00000001100000000000001110010011;
ROM[12444] <= 32'b00000000011100010010000000100011;
ROM[12445] <= 32'b00000000010000010000000100010011;
ROM[12446] <= 32'b00000011000000000000001110010011;
ROM[12447] <= 32'b00000000011100010010000000100011;
ROM[12448] <= 32'b00000000010000010000000100010011;
ROM[12449] <= 32'b00000110000000000000001110010011;
ROM[12450] <= 32'b00000000011100010010000000100011;
ROM[12451] <= 32'b00000000010000010000000100010011;
ROM[12452] <= 32'b00000000000000000000001110010011;
ROM[12453] <= 32'b00000000011100010010000000100011;
ROM[12454] <= 32'b00000000010000010000000100010011;
ROM[12455] <= 32'b00000000000000001100001110110111;
ROM[12456] <= 32'b00101110100000111000001110010011;
ROM[12457] <= 32'b00000000111000111000001110110011;
ROM[12458] <= 32'b00000000011100010010000000100011;
ROM[12459] <= 32'b00000000010000010000000100010011;
ROM[12460] <= 32'b00000000001100010010000000100011;
ROM[12461] <= 32'b00000000010000010000000100010011;
ROM[12462] <= 32'b00000000010000010010000000100011;
ROM[12463] <= 32'b00000000010000010000000100010011;
ROM[12464] <= 32'b00000000010100010010000000100011;
ROM[12465] <= 32'b00000000010000010000000100010011;
ROM[12466] <= 32'b00000000011000010010000000100011;
ROM[12467] <= 32'b00000000010000010000000100010011;
ROM[12468] <= 32'b00000001010000000000001110010011;
ROM[12469] <= 32'b00000010010000111000001110010011;
ROM[12470] <= 32'b01000000011100010000001110110011;
ROM[12471] <= 32'b00000000011100000000001000110011;
ROM[12472] <= 32'b00000000001000000000000110110011;
ROM[12473] <= 32'b00010101010000000011000011101111;
ROM[12474] <= 32'b11111111110000010000000100010011;
ROM[12475] <= 32'b00000000000000010010001110000011;
ROM[12476] <= 32'b00000000011101100010000000100011;
ROM[12477] <= 32'b00000011111100000000001110010011;
ROM[12478] <= 32'b00000000011100010010000000100011;
ROM[12479] <= 32'b00000000010000010000000100010011;
ROM[12480] <= 32'b00000111100000000000001110010011;
ROM[12481] <= 32'b00000000011100010010000000100011;
ROM[12482] <= 32'b00000000010000010000000100010011;
ROM[12483] <= 32'b00001100110000000000001110010011;
ROM[12484] <= 32'b00000000011100010010000000100011;
ROM[12485] <= 32'b00000000010000010000000100010011;
ROM[12486] <= 32'b00000000110000000000001110010011;
ROM[12487] <= 32'b00000000011100010010000000100011;
ROM[12488] <= 32'b00000000010000010000000100010011;
ROM[12489] <= 32'b00000001100000000000001110010011;
ROM[12490] <= 32'b00000000011100010010000000100011;
ROM[12491] <= 32'b00000000010000010000000100010011;
ROM[12492] <= 32'b00000011000000000000001110010011;
ROM[12493] <= 32'b00000000011100010010000000100011;
ROM[12494] <= 32'b00000000010000010000000100010011;
ROM[12495] <= 32'b00000000000000000000001110010011;
ROM[12496] <= 32'b00000000011100010010000000100011;
ROM[12497] <= 32'b00000000010000010000000100010011;
ROM[12498] <= 32'b00000011000000000000001110010011;
ROM[12499] <= 32'b00000000011100010010000000100011;
ROM[12500] <= 32'b00000000010000010000000100010011;
ROM[12501] <= 32'b00000000000000000000001110010011;
ROM[12502] <= 32'b00000000011100010010000000100011;
ROM[12503] <= 32'b00000000010000010000000100010011;
ROM[12504] <= 32'b00000000000000001100001110110111;
ROM[12505] <= 32'b00111010110000111000001110010011;
ROM[12506] <= 32'b00000000111000111000001110110011;
ROM[12507] <= 32'b00000000011100010010000000100011;
ROM[12508] <= 32'b00000000010000010000000100010011;
ROM[12509] <= 32'b00000000001100010010000000100011;
ROM[12510] <= 32'b00000000010000010000000100010011;
ROM[12511] <= 32'b00000000010000010010000000100011;
ROM[12512] <= 32'b00000000010000010000000100010011;
ROM[12513] <= 32'b00000000010100010010000000100011;
ROM[12514] <= 32'b00000000010000010000000100010011;
ROM[12515] <= 32'b00000000011000010010000000100011;
ROM[12516] <= 32'b00000000010000010000000100010011;
ROM[12517] <= 32'b00000001010000000000001110010011;
ROM[12518] <= 32'b00000010010000111000001110010011;
ROM[12519] <= 32'b01000000011100010000001110110011;
ROM[12520] <= 32'b00000000011100000000001000110011;
ROM[12521] <= 32'b00000000001000000000000110110011;
ROM[12522] <= 32'b00001001000000000011000011101111;
ROM[12523] <= 32'b11111111110000010000000100010011;
ROM[12524] <= 32'b00000000000000010010001110000011;
ROM[12525] <= 32'b00000000011101100010000000100011;
ROM[12526] <= 32'b00000100000000000000001110010011;
ROM[12527] <= 32'b00000000011100010010000000100011;
ROM[12528] <= 32'b00000000010000010000000100010011;
ROM[12529] <= 32'b00000111110000000000001110010011;
ROM[12530] <= 32'b00000000011100010010000000100011;
ROM[12531] <= 32'b00000000010000010000000100010011;
ROM[12532] <= 32'b00001100011000000000001110010011;
ROM[12533] <= 32'b00000000011100010010000000100011;
ROM[12534] <= 32'b00000000010000010000000100010011;
ROM[12535] <= 32'b00001101111000000000001110010011;
ROM[12536] <= 32'b00000000011100010010000000100011;
ROM[12537] <= 32'b00000000010000010000000100010011;
ROM[12538] <= 32'b00001101111000000000001110010011;
ROM[12539] <= 32'b00000000011100010010000000100011;
ROM[12540] <= 32'b00000000010000010000000100010011;
ROM[12541] <= 32'b00001101111000000000001110010011;
ROM[12542] <= 32'b00000000011100010010000000100011;
ROM[12543] <= 32'b00000000010000010000000100010011;
ROM[12544] <= 32'b00001100000000000000001110010011;
ROM[12545] <= 32'b00000000011100010010000000100011;
ROM[12546] <= 32'b00000000010000010000000100010011;
ROM[12547] <= 32'b00000111100000000000001110010011;
ROM[12548] <= 32'b00000000011100010010000000100011;
ROM[12549] <= 32'b00000000010000010000000100010011;
ROM[12550] <= 32'b00000000000000000000001110010011;
ROM[12551] <= 32'b00000000011100010010000000100011;
ROM[12552] <= 32'b00000000010000010000000100010011;
ROM[12553] <= 32'b00000000000000001100001110110111;
ROM[12554] <= 32'b01000111000000111000001110010011;
ROM[12555] <= 32'b00000000111000111000001110110011;
ROM[12556] <= 32'b00000000011100010010000000100011;
ROM[12557] <= 32'b00000000010000010000000100010011;
ROM[12558] <= 32'b00000000001100010010000000100011;
ROM[12559] <= 32'b00000000010000010000000100010011;
ROM[12560] <= 32'b00000000010000010010000000100011;
ROM[12561] <= 32'b00000000010000010000000100010011;
ROM[12562] <= 32'b00000000010100010010000000100011;
ROM[12563] <= 32'b00000000010000010000000100010011;
ROM[12564] <= 32'b00000000011000010010000000100011;
ROM[12565] <= 32'b00000000010000010000000100010011;
ROM[12566] <= 32'b00000001010000000000001110010011;
ROM[12567] <= 32'b00000010010000111000001110010011;
ROM[12568] <= 32'b01000000011100010000001110110011;
ROM[12569] <= 32'b00000000011100000000001000110011;
ROM[12570] <= 32'b00000000001000000000000110110011;
ROM[12571] <= 32'b01111100110100000010000011101111;
ROM[12572] <= 32'b11111111110000010000000100010011;
ROM[12573] <= 32'b00000000000000010010001110000011;
ROM[12574] <= 32'b00000000011101100010000000100011;
ROM[12575] <= 32'b00000100000100000000001110010011;
ROM[12576] <= 32'b00000000011100010010000000100011;
ROM[12577] <= 32'b00000000010000010000000100010011;
ROM[12578] <= 32'b00000011000000000000001110010011;
ROM[12579] <= 32'b00000000011100010010000000100011;
ROM[12580] <= 32'b00000000010000010000000100010011;
ROM[12581] <= 32'b00000111100000000000001110010011;
ROM[12582] <= 32'b00000000011100010010000000100011;
ROM[12583] <= 32'b00000000010000010000000100010011;
ROM[12584] <= 32'b00001100110000000000001110010011;
ROM[12585] <= 32'b00000000011100010010000000100011;
ROM[12586] <= 32'b00000000010000010000000100010011;
ROM[12587] <= 32'b00001100110000000000001110010011;
ROM[12588] <= 32'b00000000011100010010000000100011;
ROM[12589] <= 32'b00000000010000010000000100010011;
ROM[12590] <= 32'b00001111110000000000001110010011;
ROM[12591] <= 32'b00000000011100010010000000100011;
ROM[12592] <= 32'b00000000010000010000000100010011;
ROM[12593] <= 32'b00001100110000000000001110010011;
ROM[12594] <= 32'b00000000011100010010000000100011;
ROM[12595] <= 32'b00000000010000010000000100010011;
ROM[12596] <= 32'b00001100110000000000001110010011;
ROM[12597] <= 32'b00000000011100010010000000100011;
ROM[12598] <= 32'b00000000010000010000000100010011;
ROM[12599] <= 32'b00000000000000000000001110010011;
ROM[12600] <= 32'b00000000011100010010000000100011;
ROM[12601] <= 32'b00000000010000010000000100010011;
ROM[12602] <= 32'b00000000000000001100001110110111;
ROM[12603] <= 32'b01010011010000111000001110010011;
ROM[12604] <= 32'b00000000111000111000001110110011;
ROM[12605] <= 32'b00000000011100010010000000100011;
ROM[12606] <= 32'b00000000010000010000000100010011;
ROM[12607] <= 32'b00000000001100010010000000100011;
ROM[12608] <= 32'b00000000010000010000000100010011;
ROM[12609] <= 32'b00000000010000010010000000100011;
ROM[12610] <= 32'b00000000010000010000000100010011;
ROM[12611] <= 32'b00000000010100010010000000100011;
ROM[12612] <= 32'b00000000010000010000000100010011;
ROM[12613] <= 32'b00000000011000010010000000100011;
ROM[12614] <= 32'b00000000010000010000000100010011;
ROM[12615] <= 32'b00000001010000000000001110010011;
ROM[12616] <= 32'b00000010010000111000001110010011;
ROM[12617] <= 32'b01000000011100010000001110110011;
ROM[12618] <= 32'b00000000011100000000001000110011;
ROM[12619] <= 32'b00000000001000000000000110110011;
ROM[12620] <= 32'b01110000100100000010000011101111;
ROM[12621] <= 32'b11111111110000010000000100010011;
ROM[12622] <= 32'b00000000000000010010001110000011;
ROM[12623] <= 32'b00000000011101100010000000100011;
ROM[12624] <= 32'b00000100001000000000001110010011;
ROM[12625] <= 32'b00000000011100010010000000100011;
ROM[12626] <= 32'b00000000010000010000000100010011;
ROM[12627] <= 32'b00001111110000000000001110010011;
ROM[12628] <= 32'b00000000011100010010000000100011;
ROM[12629] <= 32'b00000000010000010000000100010011;
ROM[12630] <= 32'b00000110011000000000001110010011;
ROM[12631] <= 32'b00000000011100010010000000100011;
ROM[12632] <= 32'b00000000010000010000000100010011;
ROM[12633] <= 32'b00000110011000000000001110010011;
ROM[12634] <= 32'b00000000011100010010000000100011;
ROM[12635] <= 32'b00000000010000010000000100010011;
ROM[12636] <= 32'b00000111110000000000001110010011;
ROM[12637] <= 32'b00000000011100010010000000100011;
ROM[12638] <= 32'b00000000010000010000000100010011;
ROM[12639] <= 32'b00000110011000000000001110010011;
ROM[12640] <= 32'b00000000011100010010000000100011;
ROM[12641] <= 32'b00000000010000010000000100010011;
ROM[12642] <= 32'b00000110011000000000001110010011;
ROM[12643] <= 32'b00000000011100010010000000100011;
ROM[12644] <= 32'b00000000010000010000000100010011;
ROM[12645] <= 32'b00001111110000000000001110010011;
ROM[12646] <= 32'b00000000011100010010000000100011;
ROM[12647] <= 32'b00000000010000010000000100010011;
ROM[12648] <= 32'b00000000000000000000001110010011;
ROM[12649] <= 32'b00000000011100010010000000100011;
ROM[12650] <= 32'b00000000010000010000000100010011;
ROM[12651] <= 32'b00000000000000001100001110110111;
ROM[12652] <= 32'b01011111100000111000001110010011;
ROM[12653] <= 32'b00000000111000111000001110110011;
ROM[12654] <= 32'b00000000011100010010000000100011;
ROM[12655] <= 32'b00000000010000010000000100010011;
ROM[12656] <= 32'b00000000001100010010000000100011;
ROM[12657] <= 32'b00000000010000010000000100010011;
ROM[12658] <= 32'b00000000010000010010000000100011;
ROM[12659] <= 32'b00000000010000010000000100010011;
ROM[12660] <= 32'b00000000010100010010000000100011;
ROM[12661] <= 32'b00000000010000010000000100010011;
ROM[12662] <= 32'b00000000011000010010000000100011;
ROM[12663] <= 32'b00000000010000010000000100010011;
ROM[12664] <= 32'b00000001010000000000001110010011;
ROM[12665] <= 32'b00000010010000111000001110010011;
ROM[12666] <= 32'b01000000011100010000001110110011;
ROM[12667] <= 32'b00000000011100000000001000110011;
ROM[12668] <= 32'b00000000001000000000000110110011;
ROM[12669] <= 32'b01100100010100000010000011101111;
ROM[12670] <= 32'b11111111110000010000000100010011;
ROM[12671] <= 32'b00000000000000010010001110000011;
ROM[12672] <= 32'b00000000011101100010000000100011;
ROM[12673] <= 32'b00000100001100000000001110010011;
ROM[12674] <= 32'b00000000011100010010000000100011;
ROM[12675] <= 32'b00000000010000010000000100010011;
ROM[12676] <= 32'b00000011110000000000001110010011;
ROM[12677] <= 32'b00000000011100010010000000100011;
ROM[12678] <= 32'b00000000010000010000000100010011;
ROM[12679] <= 32'b00000110011000000000001110010011;
ROM[12680] <= 32'b00000000011100010010000000100011;
ROM[12681] <= 32'b00000000010000010000000100010011;
ROM[12682] <= 32'b00001100000000000000001110010011;
ROM[12683] <= 32'b00000000011100010010000000100011;
ROM[12684] <= 32'b00000000010000010000000100010011;
ROM[12685] <= 32'b00001100000000000000001110010011;
ROM[12686] <= 32'b00000000011100010010000000100011;
ROM[12687] <= 32'b00000000010000010000000100010011;
ROM[12688] <= 32'b00001100000000000000001110010011;
ROM[12689] <= 32'b00000000011100010010000000100011;
ROM[12690] <= 32'b00000000010000010000000100010011;
ROM[12691] <= 32'b00000110011000000000001110010011;
ROM[12692] <= 32'b00000000011100010010000000100011;
ROM[12693] <= 32'b00000000010000010000000100010011;
ROM[12694] <= 32'b00000011110000000000001110010011;
ROM[12695] <= 32'b00000000011100010010000000100011;
ROM[12696] <= 32'b00000000010000010000000100010011;
ROM[12697] <= 32'b00000000000000000000001110010011;
ROM[12698] <= 32'b00000000011100010010000000100011;
ROM[12699] <= 32'b00000000010000010000000100010011;
ROM[12700] <= 32'b00000000000000001100001110110111;
ROM[12701] <= 32'b01101011110000111000001110010011;
ROM[12702] <= 32'b00000000111000111000001110110011;
ROM[12703] <= 32'b00000000011100010010000000100011;
ROM[12704] <= 32'b00000000010000010000000100010011;
ROM[12705] <= 32'b00000000001100010010000000100011;
ROM[12706] <= 32'b00000000010000010000000100010011;
ROM[12707] <= 32'b00000000010000010010000000100011;
ROM[12708] <= 32'b00000000010000010000000100010011;
ROM[12709] <= 32'b00000000010100010010000000100011;
ROM[12710] <= 32'b00000000010000010000000100010011;
ROM[12711] <= 32'b00000000011000010010000000100011;
ROM[12712] <= 32'b00000000010000010000000100010011;
ROM[12713] <= 32'b00000001010000000000001110010011;
ROM[12714] <= 32'b00000010010000111000001110010011;
ROM[12715] <= 32'b01000000011100010000001110110011;
ROM[12716] <= 32'b00000000011100000000001000110011;
ROM[12717] <= 32'b00000000001000000000000110110011;
ROM[12718] <= 32'b01011000000100000010000011101111;
ROM[12719] <= 32'b11111111110000010000000100010011;
ROM[12720] <= 32'b00000000000000010010001110000011;
ROM[12721] <= 32'b00000000011101100010000000100011;
ROM[12722] <= 32'b00000100010000000000001110010011;
ROM[12723] <= 32'b00000000011100010010000000100011;
ROM[12724] <= 32'b00000000010000010000000100010011;
ROM[12725] <= 32'b00001111100000000000001110010011;
ROM[12726] <= 32'b00000000011100010010000000100011;
ROM[12727] <= 32'b00000000010000010000000100010011;
ROM[12728] <= 32'b00000110110000000000001110010011;
ROM[12729] <= 32'b00000000011100010010000000100011;
ROM[12730] <= 32'b00000000010000010000000100010011;
ROM[12731] <= 32'b00000110011000000000001110010011;
ROM[12732] <= 32'b00000000011100010010000000100011;
ROM[12733] <= 32'b00000000010000010000000100010011;
ROM[12734] <= 32'b00000110011000000000001110010011;
ROM[12735] <= 32'b00000000011100010010000000100011;
ROM[12736] <= 32'b00000000010000010000000100010011;
ROM[12737] <= 32'b00000110011000000000001110010011;
ROM[12738] <= 32'b00000000011100010010000000100011;
ROM[12739] <= 32'b00000000010000010000000100010011;
ROM[12740] <= 32'b00000110110000000000001110010011;
ROM[12741] <= 32'b00000000011100010010000000100011;
ROM[12742] <= 32'b00000000010000010000000100010011;
ROM[12743] <= 32'b00001111100000000000001110010011;
ROM[12744] <= 32'b00000000011100010010000000100011;
ROM[12745] <= 32'b00000000010000010000000100010011;
ROM[12746] <= 32'b00000000000000000000001110010011;
ROM[12747] <= 32'b00000000011100010010000000100011;
ROM[12748] <= 32'b00000000010000010000000100010011;
ROM[12749] <= 32'b00000000000000001100001110110111;
ROM[12750] <= 32'b01111000000000111000001110010011;
ROM[12751] <= 32'b00000000111000111000001110110011;
ROM[12752] <= 32'b00000000011100010010000000100011;
ROM[12753] <= 32'b00000000010000010000000100010011;
ROM[12754] <= 32'b00000000001100010010000000100011;
ROM[12755] <= 32'b00000000010000010000000100010011;
ROM[12756] <= 32'b00000000010000010010000000100011;
ROM[12757] <= 32'b00000000010000010000000100010011;
ROM[12758] <= 32'b00000000010100010010000000100011;
ROM[12759] <= 32'b00000000010000010000000100010011;
ROM[12760] <= 32'b00000000011000010010000000100011;
ROM[12761] <= 32'b00000000010000010000000100010011;
ROM[12762] <= 32'b00000001010000000000001110010011;
ROM[12763] <= 32'b00000010010000111000001110010011;
ROM[12764] <= 32'b01000000011100010000001110110011;
ROM[12765] <= 32'b00000000011100000000001000110011;
ROM[12766] <= 32'b00000000001000000000000110110011;
ROM[12767] <= 32'b01001011110100000010000011101111;
ROM[12768] <= 32'b11111111110000010000000100010011;
ROM[12769] <= 32'b00000000000000010010001110000011;
ROM[12770] <= 32'b00000000011101100010000000100011;
ROM[12771] <= 32'b00000100010100000000001110010011;
ROM[12772] <= 32'b00000000011100010010000000100011;
ROM[12773] <= 32'b00000000010000010000000100010011;
ROM[12774] <= 32'b00001111111000000000001110010011;
ROM[12775] <= 32'b00000000011100010010000000100011;
ROM[12776] <= 32'b00000000010000010000000100010011;
ROM[12777] <= 32'b00000110001000000000001110010011;
ROM[12778] <= 32'b00000000011100010010000000100011;
ROM[12779] <= 32'b00000000010000010000000100010011;
ROM[12780] <= 32'b00000110100000000000001110010011;
ROM[12781] <= 32'b00000000011100010010000000100011;
ROM[12782] <= 32'b00000000010000010000000100010011;
ROM[12783] <= 32'b00000111100000000000001110010011;
ROM[12784] <= 32'b00000000011100010010000000100011;
ROM[12785] <= 32'b00000000010000010000000100010011;
ROM[12786] <= 32'b00000110100000000000001110010011;
ROM[12787] <= 32'b00000000011100010010000000100011;
ROM[12788] <= 32'b00000000010000010000000100010011;
ROM[12789] <= 32'b00000110001000000000001110010011;
ROM[12790] <= 32'b00000000011100010010000000100011;
ROM[12791] <= 32'b00000000010000010000000100010011;
ROM[12792] <= 32'b00001111111000000000001110010011;
ROM[12793] <= 32'b00000000011100010010000000100011;
ROM[12794] <= 32'b00000000010000010000000100010011;
ROM[12795] <= 32'b00000000000000000000001110010011;
ROM[12796] <= 32'b00000000011100010010000000100011;
ROM[12797] <= 32'b00000000010000010000000100010011;
ROM[12798] <= 32'b00000000000000001101001110110111;
ROM[12799] <= 32'b10000100010000111000001110010011;
ROM[12800] <= 32'b00000000111000111000001110110011;
ROM[12801] <= 32'b00000000011100010010000000100011;
ROM[12802] <= 32'b00000000010000010000000100010011;
ROM[12803] <= 32'b00000000001100010010000000100011;
ROM[12804] <= 32'b00000000010000010000000100010011;
ROM[12805] <= 32'b00000000010000010010000000100011;
ROM[12806] <= 32'b00000000010000010000000100010011;
ROM[12807] <= 32'b00000000010100010010000000100011;
ROM[12808] <= 32'b00000000010000010000000100010011;
ROM[12809] <= 32'b00000000011000010010000000100011;
ROM[12810] <= 32'b00000000010000010000000100010011;
ROM[12811] <= 32'b00000001010000000000001110010011;
ROM[12812] <= 32'b00000010010000111000001110010011;
ROM[12813] <= 32'b01000000011100010000001110110011;
ROM[12814] <= 32'b00000000011100000000001000110011;
ROM[12815] <= 32'b00000000001000000000000110110011;
ROM[12816] <= 32'b00111111100100000010000011101111;
ROM[12817] <= 32'b11111111110000010000000100010011;
ROM[12818] <= 32'b00000000000000010010001110000011;
ROM[12819] <= 32'b00000000011101100010000000100011;
ROM[12820] <= 32'b00000100011000000000001110010011;
ROM[12821] <= 32'b00000000011100010010000000100011;
ROM[12822] <= 32'b00000000010000010000000100010011;
ROM[12823] <= 32'b00001111111000000000001110010011;
ROM[12824] <= 32'b00000000011100010010000000100011;
ROM[12825] <= 32'b00000000010000010000000100010011;
ROM[12826] <= 32'b00000110001000000000001110010011;
ROM[12827] <= 32'b00000000011100010010000000100011;
ROM[12828] <= 32'b00000000010000010000000100010011;
ROM[12829] <= 32'b00000110100000000000001110010011;
ROM[12830] <= 32'b00000000011100010010000000100011;
ROM[12831] <= 32'b00000000010000010000000100010011;
ROM[12832] <= 32'b00000111100000000000001110010011;
ROM[12833] <= 32'b00000000011100010010000000100011;
ROM[12834] <= 32'b00000000010000010000000100010011;
ROM[12835] <= 32'b00000110100000000000001110010011;
ROM[12836] <= 32'b00000000011100010010000000100011;
ROM[12837] <= 32'b00000000010000010000000100010011;
ROM[12838] <= 32'b00000110000000000000001110010011;
ROM[12839] <= 32'b00000000011100010010000000100011;
ROM[12840] <= 32'b00000000010000010000000100010011;
ROM[12841] <= 32'b00001111000000000000001110010011;
ROM[12842] <= 32'b00000000011100010010000000100011;
ROM[12843] <= 32'b00000000010000010000000100010011;
ROM[12844] <= 32'b00000000000000000000001110010011;
ROM[12845] <= 32'b00000000011100010010000000100011;
ROM[12846] <= 32'b00000000010000010000000100010011;
ROM[12847] <= 32'b00000000000000001101001110110111;
ROM[12848] <= 32'b10010000100000111000001110010011;
ROM[12849] <= 32'b00000000111000111000001110110011;
ROM[12850] <= 32'b00000000011100010010000000100011;
ROM[12851] <= 32'b00000000010000010000000100010011;
ROM[12852] <= 32'b00000000001100010010000000100011;
ROM[12853] <= 32'b00000000010000010000000100010011;
ROM[12854] <= 32'b00000000010000010010000000100011;
ROM[12855] <= 32'b00000000010000010000000100010011;
ROM[12856] <= 32'b00000000010100010010000000100011;
ROM[12857] <= 32'b00000000010000010000000100010011;
ROM[12858] <= 32'b00000000011000010010000000100011;
ROM[12859] <= 32'b00000000010000010000000100010011;
ROM[12860] <= 32'b00000001010000000000001110010011;
ROM[12861] <= 32'b00000010010000111000001110010011;
ROM[12862] <= 32'b01000000011100010000001110110011;
ROM[12863] <= 32'b00000000011100000000001000110011;
ROM[12864] <= 32'b00000000001000000000000110110011;
ROM[12865] <= 32'b00110011010100000010000011101111;
ROM[12866] <= 32'b11111111110000010000000100010011;
ROM[12867] <= 32'b00000000000000010010001110000011;
ROM[12868] <= 32'b00000000011101100010000000100011;
ROM[12869] <= 32'b00000100011100000000001110010011;
ROM[12870] <= 32'b00000000011100010010000000100011;
ROM[12871] <= 32'b00000000010000010000000100010011;
ROM[12872] <= 32'b00000011110000000000001110010011;
ROM[12873] <= 32'b00000000011100010010000000100011;
ROM[12874] <= 32'b00000000010000010000000100010011;
ROM[12875] <= 32'b00000110011000000000001110010011;
ROM[12876] <= 32'b00000000011100010010000000100011;
ROM[12877] <= 32'b00000000010000010000000100010011;
ROM[12878] <= 32'b00001100000000000000001110010011;
ROM[12879] <= 32'b00000000011100010010000000100011;
ROM[12880] <= 32'b00000000010000010000000100010011;
ROM[12881] <= 32'b00001100000000000000001110010011;
ROM[12882] <= 32'b00000000011100010010000000100011;
ROM[12883] <= 32'b00000000010000010000000100010011;
ROM[12884] <= 32'b00001100111000000000001110010011;
ROM[12885] <= 32'b00000000011100010010000000100011;
ROM[12886] <= 32'b00000000010000010000000100010011;
ROM[12887] <= 32'b00000110011000000000001110010011;
ROM[12888] <= 32'b00000000011100010010000000100011;
ROM[12889] <= 32'b00000000010000010000000100010011;
ROM[12890] <= 32'b00000011111000000000001110010011;
ROM[12891] <= 32'b00000000011100010010000000100011;
ROM[12892] <= 32'b00000000010000010000000100010011;
ROM[12893] <= 32'b00000000000000000000001110010011;
ROM[12894] <= 32'b00000000011100010010000000100011;
ROM[12895] <= 32'b00000000010000010000000100010011;
ROM[12896] <= 32'b00000000000000001101001110110111;
ROM[12897] <= 32'b10011100110000111000001110010011;
ROM[12898] <= 32'b00000000111000111000001110110011;
ROM[12899] <= 32'b00000000011100010010000000100011;
ROM[12900] <= 32'b00000000010000010000000100010011;
ROM[12901] <= 32'b00000000001100010010000000100011;
ROM[12902] <= 32'b00000000010000010000000100010011;
ROM[12903] <= 32'b00000000010000010010000000100011;
ROM[12904] <= 32'b00000000010000010000000100010011;
ROM[12905] <= 32'b00000000010100010010000000100011;
ROM[12906] <= 32'b00000000010000010000000100010011;
ROM[12907] <= 32'b00000000011000010010000000100011;
ROM[12908] <= 32'b00000000010000010000000100010011;
ROM[12909] <= 32'b00000001010000000000001110010011;
ROM[12910] <= 32'b00000010010000111000001110010011;
ROM[12911] <= 32'b01000000011100010000001110110011;
ROM[12912] <= 32'b00000000011100000000001000110011;
ROM[12913] <= 32'b00000000001000000000000110110011;
ROM[12914] <= 32'b00100111000100000010000011101111;
ROM[12915] <= 32'b11111111110000010000000100010011;
ROM[12916] <= 32'b00000000000000010010001110000011;
ROM[12917] <= 32'b00000000011101100010000000100011;
ROM[12918] <= 32'b00000100100000000000001110010011;
ROM[12919] <= 32'b00000000011100010010000000100011;
ROM[12920] <= 32'b00000000010000010000000100010011;
ROM[12921] <= 32'b00001100110000000000001110010011;
ROM[12922] <= 32'b00000000011100010010000000100011;
ROM[12923] <= 32'b00000000010000010000000100010011;
ROM[12924] <= 32'b00001100110000000000001110010011;
ROM[12925] <= 32'b00000000011100010010000000100011;
ROM[12926] <= 32'b00000000010000010000000100010011;
ROM[12927] <= 32'b00001100110000000000001110010011;
ROM[12928] <= 32'b00000000011100010010000000100011;
ROM[12929] <= 32'b00000000010000010000000100010011;
ROM[12930] <= 32'b00001111110000000000001110010011;
ROM[12931] <= 32'b00000000011100010010000000100011;
ROM[12932] <= 32'b00000000010000010000000100010011;
ROM[12933] <= 32'b00001100110000000000001110010011;
ROM[12934] <= 32'b00000000011100010010000000100011;
ROM[12935] <= 32'b00000000010000010000000100010011;
ROM[12936] <= 32'b00001100110000000000001110010011;
ROM[12937] <= 32'b00000000011100010010000000100011;
ROM[12938] <= 32'b00000000010000010000000100010011;
ROM[12939] <= 32'b00001100110000000000001110010011;
ROM[12940] <= 32'b00000000011100010010000000100011;
ROM[12941] <= 32'b00000000010000010000000100010011;
ROM[12942] <= 32'b00000000000000000000001110010011;
ROM[12943] <= 32'b00000000011100010010000000100011;
ROM[12944] <= 32'b00000000010000010000000100010011;
ROM[12945] <= 32'b00000000000000001101001110110111;
ROM[12946] <= 32'b10101001000000111000001110010011;
ROM[12947] <= 32'b00000000111000111000001110110011;
ROM[12948] <= 32'b00000000011100010010000000100011;
ROM[12949] <= 32'b00000000010000010000000100010011;
ROM[12950] <= 32'b00000000001100010010000000100011;
ROM[12951] <= 32'b00000000010000010000000100010011;
ROM[12952] <= 32'b00000000010000010010000000100011;
ROM[12953] <= 32'b00000000010000010000000100010011;
ROM[12954] <= 32'b00000000010100010010000000100011;
ROM[12955] <= 32'b00000000010000010000000100010011;
ROM[12956] <= 32'b00000000011000010010000000100011;
ROM[12957] <= 32'b00000000010000010000000100010011;
ROM[12958] <= 32'b00000001010000000000001110010011;
ROM[12959] <= 32'b00000010010000111000001110010011;
ROM[12960] <= 32'b01000000011100010000001110110011;
ROM[12961] <= 32'b00000000011100000000001000110011;
ROM[12962] <= 32'b00000000001000000000000110110011;
ROM[12963] <= 32'b00011010110100000010000011101111;
ROM[12964] <= 32'b11111111110000010000000100010011;
ROM[12965] <= 32'b00000000000000010010001110000011;
ROM[12966] <= 32'b00000000011101100010000000100011;
ROM[12967] <= 32'b00000100100100000000001110010011;
ROM[12968] <= 32'b00000000011100010010000000100011;
ROM[12969] <= 32'b00000000010000010000000100010011;
ROM[12970] <= 32'b00000111100000000000001110010011;
ROM[12971] <= 32'b00000000011100010010000000100011;
ROM[12972] <= 32'b00000000010000010000000100010011;
ROM[12973] <= 32'b00000011000000000000001110010011;
ROM[12974] <= 32'b00000000011100010010000000100011;
ROM[12975] <= 32'b00000000010000010000000100010011;
ROM[12976] <= 32'b00000011000000000000001110010011;
ROM[12977] <= 32'b00000000011100010010000000100011;
ROM[12978] <= 32'b00000000010000010000000100010011;
ROM[12979] <= 32'b00000011000000000000001110010011;
ROM[12980] <= 32'b00000000011100010010000000100011;
ROM[12981] <= 32'b00000000010000010000000100010011;
ROM[12982] <= 32'b00000011000000000000001110010011;
ROM[12983] <= 32'b00000000011100010010000000100011;
ROM[12984] <= 32'b00000000010000010000000100010011;
ROM[12985] <= 32'b00000011000000000000001110010011;
ROM[12986] <= 32'b00000000011100010010000000100011;
ROM[12987] <= 32'b00000000010000010000000100010011;
ROM[12988] <= 32'b00000111100000000000001110010011;
ROM[12989] <= 32'b00000000011100010010000000100011;
ROM[12990] <= 32'b00000000010000010000000100010011;
ROM[12991] <= 32'b00000000000000000000001110010011;
ROM[12992] <= 32'b00000000011100010010000000100011;
ROM[12993] <= 32'b00000000010000010000000100010011;
ROM[12994] <= 32'b00000000000000001101001110110111;
ROM[12995] <= 32'b10110101010000111000001110010011;
ROM[12996] <= 32'b00000000111000111000001110110011;
ROM[12997] <= 32'b00000000011100010010000000100011;
ROM[12998] <= 32'b00000000010000010000000100010011;
ROM[12999] <= 32'b00000000001100010010000000100011;
ROM[13000] <= 32'b00000000010000010000000100010011;
ROM[13001] <= 32'b00000000010000010010000000100011;
ROM[13002] <= 32'b00000000010000010000000100010011;
ROM[13003] <= 32'b00000000010100010010000000100011;
ROM[13004] <= 32'b00000000010000010000000100010011;
ROM[13005] <= 32'b00000000011000010010000000100011;
ROM[13006] <= 32'b00000000010000010000000100010011;
ROM[13007] <= 32'b00000001010000000000001110010011;
ROM[13008] <= 32'b00000010010000111000001110010011;
ROM[13009] <= 32'b01000000011100010000001110110011;
ROM[13010] <= 32'b00000000011100000000001000110011;
ROM[13011] <= 32'b00000000001000000000000110110011;
ROM[13012] <= 32'b00001110100100000010000011101111;
ROM[13013] <= 32'b11111111110000010000000100010011;
ROM[13014] <= 32'b00000000000000010010001110000011;
ROM[13015] <= 32'b00000000011101100010000000100011;
ROM[13016] <= 32'b00000100101000000000001110010011;
ROM[13017] <= 32'b00000000011100010010000000100011;
ROM[13018] <= 32'b00000000010000010000000100010011;
ROM[13019] <= 32'b00000001111000000000001110010011;
ROM[13020] <= 32'b00000000011100010010000000100011;
ROM[13021] <= 32'b00000000010000010000000100010011;
ROM[13022] <= 32'b00000000110000000000001110010011;
ROM[13023] <= 32'b00000000011100010010000000100011;
ROM[13024] <= 32'b00000000010000010000000100010011;
ROM[13025] <= 32'b00000000110000000000001110010011;
ROM[13026] <= 32'b00000000011100010010000000100011;
ROM[13027] <= 32'b00000000010000010000000100010011;
ROM[13028] <= 32'b00000000110000000000001110010011;
ROM[13029] <= 32'b00000000011100010010000000100011;
ROM[13030] <= 32'b00000000010000010000000100010011;
ROM[13031] <= 32'b00001100110000000000001110010011;
ROM[13032] <= 32'b00000000011100010010000000100011;
ROM[13033] <= 32'b00000000010000010000000100010011;
ROM[13034] <= 32'b00001100110000000000001110010011;
ROM[13035] <= 32'b00000000011100010010000000100011;
ROM[13036] <= 32'b00000000010000010000000100010011;
ROM[13037] <= 32'b00000111100000000000001110010011;
ROM[13038] <= 32'b00000000011100010010000000100011;
ROM[13039] <= 32'b00000000010000010000000100010011;
ROM[13040] <= 32'b00000000000000000000001110010011;
ROM[13041] <= 32'b00000000011100010010000000100011;
ROM[13042] <= 32'b00000000010000010000000100010011;
ROM[13043] <= 32'b00000000000000001101001110110111;
ROM[13044] <= 32'b11000001100000111000001110010011;
ROM[13045] <= 32'b00000000111000111000001110110011;
ROM[13046] <= 32'b00000000011100010010000000100011;
ROM[13047] <= 32'b00000000010000010000000100010011;
ROM[13048] <= 32'b00000000001100010010000000100011;
ROM[13049] <= 32'b00000000010000010000000100010011;
ROM[13050] <= 32'b00000000010000010010000000100011;
ROM[13051] <= 32'b00000000010000010000000100010011;
ROM[13052] <= 32'b00000000010100010010000000100011;
ROM[13053] <= 32'b00000000010000010000000100010011;
ROM[13054] <= 32'b00000000011000010010000000100011;
ROM[13055] <= 32'b00000000010000010000000100010011;
ROM[13056] <= 32'b00000001010000000000001110010011;
ROM[13057] <= 32'b00000010010000111000001110010011;
ROM[13058] <= 32'b01000000011100010000001110110011;
ROM[13059] <= 32'b00000000011100000000001000110011;
ROM[13060] <= 32'b00000000001000000000000110110011;
ROM[13061] <= 32'b00000010010100000010000011101111;
ROM[13062] <= 32'b11111111110000010000000100010011;
ROM[13063] <= 32'b00000000000000010010001110000011;
ROM[13064] <= 32'b00000000011101100010000000100011;
ROM[13065] <= 32'b00000100101100000000001110010011;
ROM[13066] <= 32'b00000000011100010010000000100011;
ROM[13067] <= 32'b00000000010000010000000100010011;
ROM[13068] <= 32'b00001110011000000000001110010011;
ROM[13069] <= 32'b00000000011100010010000000100011;
ROM[13070] <= 32'b00000000010000010000000100010011;
ROM[13071] <= 32'b00000110011000000000001110010011;
ROM[13072] <= 32'b00000000011100010010000000100011;
ROM[13073] <= 32'b00000000010000010000000100010011;
ROM[13074] <= 32'b00000110110000000000001110010011;
ROM[13075] <= 32'b00000000011100010010000000100011;
ROM[13076] <= 32'b00000000010000010000000100010011;
ROM[13077] <= 32'b00000111100000000000001110010011;
ROM[13078] <= 32'b00000000011100010010000000100011;
ROM[13079] <= 32'b00000000010000010000000100010011;
ROM[13080] <= 32'b00000110110000000000001110010011;
ROM[13081] <= 32'b00000000011100010010000000100011;
ROM[13082] <= 32'b00000000010000010000000100010011;
ROM[13083] <= 32'b00000110011000000000001110010011;
ROM[13084] <= 32'b00000000011100010010000000100011;
ROM[13085] <= 32'b00000000010000010000000100010011;
ROM[13086] <= 32'b00001110011000000000001110010011;
ROM[13087] <= 32'b00000000011100010010000000100011;
ROM[13088] <= 32'b00000000010000010000000100010011;
ROM[13089] <= 32'b00000000000000000000001110010011;
ROM[13090] <= 32'b00000000011100010010000000100011;
ROM[13091] <= 32'b00000000010000010000000100010011;
ROM[13092] <= 32'b00000000000000001101001110110111;
ROM[13093] <= 32'b11001101110000111000001110010011;
ROM[13094] <= 32'b00000000111000111000001110110011;
ROM[13095] <= 32'b00000000011100010010000000100011;
ROM[13096] <= 32'b00000000010000010000000100010011;
ROM[13097] <= 32'b00000000001100010010000000100011;
ROM[13098] <= 32'b00000000010000010000000100010011;
ROM[13099] <= 32'b00000000010000010010000000100011;
ROM[13100] <= 32'b00000000010000010000000100010011;
ROM[13101] <= 32'b00000000010100010010000000100011;
ROM[13102] <= 32'b00000000010000010000000100010011;
ROM[13103] <= 32'b00000000011000010010000000100011;
ROM[13104] <= 32'b00000000010000010000000100010011;
ROM[13105] <= 32'b00000001010000000000001110010011;
ROM[13106] <= 32'b00000010010000111000001110010011;
ROM[13107] <= 32'b01000000011100010000001110110011;
ROM[13108] <= 32'b00000000011100000000001000110011;
ROM[13109] <= 32'b00000000001000000000000110110011;
ROM[13110] <= 32'b01110110000000000010000011101111;
ROM[13111] <= 32'b11111111110000010000000100010011;
ROM[13112] <= 32'b00000000000000010010001110000011;
ROM[13113] <= 32'b00000000011101100010000000100011;
ROM[13114] <= 32'b00000100110000000000001110010011;
ROM[13115] <= 32'b00000000011100010010000000100011;
ROM[13116] <= 32'b00000000010000010000000100010011;
ROM[13117] <= 32'b00001111000000000000001110010011;
ROM[13118] <= 32'b00000000011100010010000000100011;
ROM[13119] <= 32'b00000000010000010000000100010011;
ROM[13120] <= 32'b00000110000000000000001110010011;
ROM[13121] <= 32'b00000000011100010010000000100011;
ROM[13122] <= 32'b00000000010000010000000100010011;
ROM[13123] <= 32'b00000110000000000000001110010011;
ROM[13124] <= 32'b00000000011100010010000000100011;
ROM[13125] <= 32'b00000000010000010000000100010011;
ROM[13126] <= 32'b00000110000000000000001110010011;
ROM[13127] <= 32'b00000000011100010010000000100011;
ROM[13128] <= 32'b00000000010000010000000100010011;
ROM[13129] <= 32'b00000110001000000000001110010011;
ROM[13130] <= 32'b00000000011100010010000000100011;
ROM[13131] <= 32'b00000000010000010000000100010011;
ROM[13132] <= 32'b00000110011000000000001110010011;
ROM[13133] <= 32'b00000000011100010010000000100011;
ROM[13134] <= 32'b00000000010000010000000100010011;
ROM[13135] <= 32'b00001111111000000000001110010011;
ROM[13136] <= 32'b00000000011100010010000000100011;
ROM[13137] <= 32'b00000000010000010000000100010011;
ROM[13138] <= 32'b00000000000000000000001110010011;
ROM[13139] <= 32'b00000000011100010010000000100011;
ROM[13140] <= 32'b00000000010000010000000100010011;
ROM[13141] <= 32'b00000000000000001101001110110111;
ROM[13142] <= 32'b11011010000000111000001110010011;
ROM[13143] <= 32'b00000000111000111000001110110011;
ROM[13144] <= 32'b00000000011100010010000000100011;
ROM[13145] <= 32'b00000000010000010000000100010011;
ROM[13146] <= 32'b00000000001100010010000000100011;
ROM[13147] <= 32'b00000000010000010000000100010011;
ROM[13148] <= 32'b00000000010000010010000000100011;
ROM[13149] <= 32'b00000000010000010000000100010011;
ROM[13150] <= 32'b00000000010100010010000000100011;
ROM[13151] <= 32'b00000000010000010000000100010011;
ROM[13152] <= 32'b00000000011000010010000000100011;
ROM[13153] <= 32'b00000000010000010000000100010011;
ROM[13154] <= 32'b00000001010000000000001110010011;
ROM[13155] <= 32'b00000010010000111000001110010011;
ROM[13156] <= 32'b01000000011100010000001110110011;
ROM[13157] <= 32'b00000000011100000000001000110011;
ROM[13158] <= 32'b00000000001000000000000110110011;
ROM[13159] <= 32'b01101001110000000010000011101111;
ROM[13160] <= 32'b11111111110000010000000100010011;
ROM[13161] <= 32'b00000000000000010010001110000011;
ROM[13162] <= 32'b00000000011101100010000000100011;
ROM[13163] <= 32'b00000100110100000000001110010011;
ROM[13164] <= 32'b00000000011100010010000000100011;
ROM[13165] <= 32'b00000000010000010000000100010011;
ROM[13166] <= 32'b00001100011000000000001110010011;
ROM[13167] <= 32'b00000000011100010010000000100011;
ROM[13168] <= 32'b00000000010000010000000100010011;
ROM[13169] <= 32'b00001110111000000000001110010011;
ROM[13170] <= 32'b00000000011100010010000000100011;
ROM[13171] <= 32'b00000000010000010000000100010011;
ROM[13172] <= 32'b00001111111000000000001110010011;
ROM[13173] <= 32'b00000000011100010010000000100011;
ROM[13174] <= 32'b00000000010000010000000100010011;
ROM[13175] <= 32'b00001111111000000000001110010011;
ROM[13176] <= 32'b00000000011100010010000000100011;
ROM[13177] <= 32'b00000000010000010000000100010011;
ROM[13178] <= 32'b00001101011000000000001110010011;
ROM[13179] <= 32'b00000000011100010010000000100011;
ROM[13180] <= 32'b00000000010000010000000100010011;
ROM[13181] <= 32'b00001100011000000000001110010011;
ROM[13182] <= 32'b00000000011100010010000000100011;
ROM[13183] <= 32'b00000000010000010000000100010011;
ROM[13184] <= 32'b00001100011000000000001110010011;
ROM[13185] <= 32'b00000000011100010010000000100011;
ROM[13186] <= 32'b00000000010000010000000100010011;
ROM[13187] <= 32'b00000000000000000000001110010011;
ROM[13188] <= 32'b00000000011100010010000000100011;
ROM[13189] <= 32'b00000000010000010000000100010011;
ROM[13190] <= 32'b00000000000000001101001110110111;
ROM[13191] <= 32'b11100110010000111000001110010011;
ROM[13192] <= 32'b00000000111000111000001110110011;
ROM[13193] <= 32'b00000000011100010010000000100011;
ROM[13194] <= 32'b00000000010000010000000100010011;
ROM[13195] <= 32'b00000000001100010010000000100011;
ROM[13196] <= 32'b00000000010000010000000100010011;
ROM[13197] <= 32'b00000000010000010010000000100011;
ROM[13198] <= 32'b00000000010000010000000100010011;
ROM[13199] <= 32'b00000000010100010010000000100011;
ROM[13200] <= 32'b00000000010000010000000100010011;
ROM[13201] <= 32'b00000000011000010010000000100011;
ROM[13202] <= 32'b00000000010000010000000100010011;
ROM[13203] <= 32'b00000001010000000000001110010011;
ROM[13204] <= 32'b00000010010000111000001110010011;
ROM[13205] <= 32'b01000000011100010000001110110011;
ROM[13206] <= 32'b00000000011100000000001000110011;
ROM[13207] <= 32'b00000000001000000000000110110011;
ROM[13208] <= 32'b01011101100000000010000011101111;
ROM[13209] <= 32'b11111111110000010000000100010011;
ROM[13210] <= 32'b00000000000000010010001110000011;
ROM[13211] <= 32'b00000000011101100010000000100011;
ROM[13212] <= 32'b00000100111000000000001110010011;
ROM[13213] <= 32'b00000000011100010010000000100011;
ROM[13214] <= 32'b00000000010000010000000100010011;
ROM[13215] <= 32'b00001100011000000000001110010011;
ROM[13216] <= 32'b00000000011100010010000000100011;
ROM[13217] <= 32'b00000000010000010000000100010011;
ROM[13218] <= 32'b00001110011000000000001110010011;
ROM[13219] <= 32'b00000000011100010010000000100011;
ROM[13220] <= 32'b00000000010000010000000100010011;
ROM[13221] <= 32'b00001111011000000000001110010011;
ROM[13222] <= 32'b00000000011100010010000000100011;
ROM[13223] <= 32'b00000000010000010000000100010011;
ROM[13224] <= 32'b00001101111000000000001110010011;
ROM[13225] <= 32'b00000000011100010010000000100011;
ROM[13226] <= 32'b00000000010000010000000100010011;
ROM[13227] <= 32'b00001100111000000000001110010011;
ROM[13228] <= 32'b00000000011100010010000000100011;
ROM[13229] <= 32'b00000000010000010000000100010011;
ROM[13230] <= 32'b00001100011000000000001110010011;
ROM[13231] <= 32'b00000000011100010010000000100011;
ROM[13232] <= 32'b00000000010000010000000100010011;
ROM[13233] <= 32'b00001100011000000000001110010011;
ROM[13234] <= 32'b00000000011100010010000000100011;
ROM[13235] <= 32'b00000000010000010000000100010011;
ROM[13236] <= 32'b00000000000000000000001110010011;
ROM[13237] <= 32'b00000000011100010010000000100011;
ROM[13238] <= 32'b00000000010000010000000100010011;
ROM[13239] <= 32'b00000000000000001101001110110111;
ROM[13240] <= 32'b11110010100000111000001110010011;
ROM[13241] <= 32'b00000000111000111000001110110011;
ROM[13242] <= 32'b00000000011100010010000000100011;
ROM[13243] <= 32'b00000000010000010000000100010011;
ROM[13244] <= 32'b00000000001100010010000000100011;
ROM[13245] <= 32'b00000000010000010000000100010011;
ROM[13246] <= 32'b00000000010000010010000000100011;
ROM[13247] <= 32'b00000000010000010000000100010011;
ROM[13248] <= 32'b00000000010100010010000000100011;
ROM[13249] <= 32'b00000000010000010000000100010011;
ROM[13250] <= 32'b00000000011000010010000000100011;
ROM[13251] <= 32'b00000000010000010000000100010011;
ROM[13252] <= 32'b00000001010000000000001110010011;
ROM[13253] <= 32'b00000010010000111000001110010011;
ROM[13254] <= 32'b01000000011100010000001110110011;
ROM[13255] <= 32'b00000000011100000000001000110011;
ROM[13256] <= 32'b00000000001000000000000110110011;
ROM[13257] <= 32'b01010001010000000010000011101111;
ROM[13258] <= 32'b11111111110000010000000100010011;
ROM[13259] <= 32'b00000000000000010010001110000011;
ROM[13260] <= 32'b00000000011101100010000000100011;
ROM[13261] <= 32'b00000100111100000000001110010011;
ROM[13262] <= 32'b00000000011100010010000000100011;
ROM[13263] <= 32'b00000000010000010000000100010011;
ROM[13264] <= 32'b00000011100000000000001110010011;
ROM[13265] <= 32'b00000000011100010010000000100011;
ROM[13266] <= 32'b00000000010000010000000100010011;
ROM[13267] <= 32'b00000110110000000000001110010011;
ROM[13268] <= 32'b00000000011100010010000000100011;
ROM[13269] <= 32'b00000000010000010000000100010011;
ROM[13270] <= 32'b00001100011000000000001110010011;
ROM[13271] <= 32'b00000000011100010010000000100011;
ROM[13272] <= 32'b00000000010000010000000100010011;
ROM[13273] <= 32'b00001100011000000000001110010011;
ROM[13274] <= 32'b00000000011100010010000000100011;
ROM[13275] <= 32'b00000000010000010000000100010011;
ROM[13276] <= 32'b00001100011000000000001110010011;
ROM[13277] <= 32'b00000000011100010010000000100011;
ROM[13278] <= 32'b00000000010000010000000100010011;
ROM[13279] <= 32'b00000110110000000000001110010011;
ROM[13280] <= 32'b00000000011100010010000000100011;
ROM[13281] <= 32'b00000000010000010000000100010011;
ROM[13282] <= 32'b00000011100000000000001110010011;
ROM[13283] <= 32'b00000000011100010010000000100011;
ROM[13284] <= 32'b00000000010000010000000100010011;
ROM[13285] <= 32'b00000000000000000000001110010011;
ROM[13286] <= 32'b00000000011100010010000000100011;
ROM[13287] <= 32'b00000000010000010000000100010011;
ROM[13288] <= 32'b00000000000000001101001110110111;
ROM[13289] <= 32'b11111110110000111000001110010011;
ROM[13290] <= 32'b00000000111000111000001110110011;
ROM[13291] <= 32'b00000000011100010010000000100011;
ROM[13292] <= 32'b00000000010000010000000100010011;
ROM[13293] <= 32'b00000000001100010010000000100011;
ROM[13294] <= 32'b00000000010000010000000100010011;
ROM[13295] <= 32'b00000000010000010010000000100011;
ROM[13296] <= 32'b00000000010000010000000100010011;
ROM[13297] <= 32'b00000000010100010010000000100011;
ROM[13298] <= 32'b00000000010000010000000100010011;
ROM[13299] <= 32'b00000000011000010010000000100011;
ROM[13300] <= 32'b00000000010000010000000100010011;
ROM[13301] <= 32'b00000001010000000000001110010011;
ROM[13302] <= 32'b00000010010000111000001110010011;
ROM[13303] <= 32'b01000000011100010000001110110011;
ROM[13304] <= 32'b00000000011100000000001000110011;
ROM[13305] <= 32'b00000000001000000000000110110011;
ROM[13306] <= 32'b01000101000000000010000011101111;
ROM[13307] <= 32'b11111111110000010000000100010011;
ROM[13308] <= 32'b00000000000000010010001110000011;
ROM[13309] <= 32'b00000000011101100010000000100011;
ROM[13310] <= 32'b00000101000000000000001110010011;
ROM[13311] <= 32'b00000000011100010010000000100011;
ROM[13312] <= 32'b00000000010000010000000100010011;
ROM[13313] <= 32'b00001111110000000000001110010011;
ROM[13314] <= 32'b00000000011100010010000000100011;
ROM[13315] <= 32'b00000000010000010000000100010011;
ROM[13316] <= 32'b00000110011000000000001110010011;
ROM[13317] <= 32'b00000000011100010010000000100011;
ROM[13318] <= 32'b00000000010000010000000100010011;
ROM[13319] <= 32'b00000110011000000000001110010011;
ROM[13320] <= 32'b00000000011100010010000000100011;
ROM[13321] <= 32'b00000000010000010000000100010011;
ROM[13322] <= 32'b00000111110000000000001110010011;
ROM[13323] <= 32'b00000000011100010010000000100011;
ROM[13324] <= 32'b00000000010000010000000100010011;
ROM[13325] <= 32'b00000110000000000000001110010011;
ROM[13326] <= 32'b00000000011100010010000000100011;
ROM[13327] <= 32'b00000000010000010000000100010011;
ROM[13328] <= 32'b00000110000000000000001110010011;
ROM[13329] <= 32'b00000000011100010010000000100011;
ROM[13330] <= 32'b00000000010000010000000100010011;
ROM[13331] <= 32'b00001111000000000000001110010011;
ROM[13332] <= 32'b00000000011100010010000000100011;
ROM[13333] <= 32'b00000000010000010000000100010011;
ROM[13334] <= 32'b00000000000000000000001110010011;
ROM[13335] <= 32'b00000000011100010010000000100011;
ROM[13336] <= 32'b00000000010000010000000100010011;
ROM[13337] <= 32'b00000000000000001101001110110111;
ROM[13338] <= 32'b00001011000000111000001110010011;
ROM[13339] <= 32'b00000000111000111000001110110011;
ROM[13340] <= 32'b00000000011100010010000000100011;
ROM[13341] <= 32'b00000000010000010000000100010011;
ROM[13342] <= 32'b00000000001100010010000000100011;
ROM[13343] <= 32'b00000000010000010000000100010011;
ROM[13344] <= 32'b00000000010000010010000000100011;
ROM[13345] <= 32'b00000000010000010000000100010011;
ROM[13346] <= 32'b00000000010100010010000000100011;
ROM[13347] <= 32'b00000000010000010000000100010011;
ROM[13348] <= 32'b00000000011000010010000000100011;
ROM[13349] <= 32'b00000000010000010000000100010011;
ROM[13350] <= 32'b00000001010000000000001110010011;
ROM[13351] <= 32'b00000010010000111000001110010011;
ROM[13352] <= 32'b01000000011100010000001110110011;
ROM[13353] <= 32'b00000000011100000000001000110011;
ROM[13354] <= 32'b00000000001000000000000110110011;
ROM[13355] <= 32'b00111000110000000010000011101111;
ROM[13356] <= 32'b11111111110000010000000100010011;
ROM[13357] <= 32'b00000000000000010010001110000011;
ROM[13358] <= 32'b00000000011101100010000000100011;
ROM[13359] <= 32'b00000101000100000000001110010011;
ROM[13360] <= 32'b00000000011100010010000000100011;
ROM[13361] <= 32'b00000000010000010000000100010011;
ROM[13362] <= 32'b00000111100000000000001110010011;
ROM[13363] <= 32'b00000000011100010010000000100011;
ROM[13364] <= 32'b00000000010000010000000100010011;
ROM[13365] <= 32'b00001100110000000000001110010011;
ROM[13366] <= 32'b00000000011100010010000000100011;
ROM[13367] <= 32'b00000000010000010000000100010011;
ROM[13368] <= 32'b00001100110000000000001110010011;
ROM[13369] <= 32'b00000000011100010010000000100011;
ROM[13370] <= 32'b00000000010000010000000100010011;
ROM[13371] <= 32'b00001100110000000000001110010011;
ROM[13372] <= 32'b00000000011100010010000000100011;
ROM[13373] <= 32'b00000000010000010000000100010011;
ROM[13374] <= 32'b00001101110000000000001110010011;
ROM[13375] <= 32'b00000000011100010010000000100011;
ROM[13376] <= 32'b00000000010000010000000100010011;
ROM[13377] <= 32'b00000111100000000000001110010011;
ROM[13378] <= 32'b00000000011100010010000000100011;
ROM[13379] <= 32'b00000000010000010000000100010011;
ROM[13380] <= 32'b00000001110000000000001110010011;
ROM[13381] <= 32'b00000000011100010010000000100011;
ROM[13382] <= 32'b00000000010000010000000100010011;
ROM[13383] <= 32'b00000000000000000000001110010011;
ROM[13384] <= 32'b00000000011100010010000000100011;
ROM[13385] <= 32'b00000000010000010000000100010011;
ROM[13386] <= 32'b00000000000000001101001110110111;
ROM[13387] <= 32'b00010111010000111000001110010011;
ROM[13388] <= 32'b00000000111000111000001110110011;
ROM[13389] <= 32'b00000000011100010010000000100011;
ROM[13390] <= 32'b00000000010000010000000100010011;
ROM[13391] <= 32'b00000000001100010010000000100011;
ROM[13392] <= 32'b00000000010000010000000100010011;
ROM[13393] <= 32'b00000000010000010010000000100011;
ROM[13394] <= 32'b00000000010000010000000100010011;
ROM[13395] <= 32'b00000000010100010010000000100011;
ROM[13396] <= 32'b00000000010000010000000100010011;
ROM[13397] <= 32'b00000000011000010010000000100011;
ROM[13398] <= 32'b00000000010000010000000100010011;
ROM[13399] <= 32'b00000001010000000000001110010011;
ROM[13400] <= 32'b00000010010000111000001110010011;
ROM[13401] <= 32'b01000000011100010000001110110011;
ROM[13402] <= 32'b00000000011100000000001000110011;
ROM[13403] <= 32'b00000000001000000000000110110011;
ROM[13404] <= 32'b00101100100000000010000011101111;
ROM[13405] <= 32'b11111111110000010000000100010011;
ROM[13406] <= 32'b00000000000000010010001110000011;
ROM[13407] <= 32'b00000000011101100010000000100011;
ROM[13408] <= 32'b00000101001000000000001110010011;
ROM[13409] <= 32'b00000000011100010010000000100011;
ROM[13410] <= 32'b00000000010000010000000100010011;
ROM[13411] <= 32'b00001111110000000000001110010011;
ROM[13412] <= 32'b00000000011100010010000000100011;
ROM[13413] <= 32'b00000000010000010000000100010011;
ROM[13414] <= 32'b00000110011000000000001110010011;
ROM[13415] <= 32'b00000000011100010010000000100011;
ROM[13416] <= 32'b00000000010000010000000100010011;
ROM[13417] <= 32'b00000110011000000000001110010011;
ROM[13418] <= 32'b00000000011100010010000000100011;
ROM[13419] <= 32'b00000000010000010000000100010011;
ROM[13420] <= 32'b00000111110000000000001110010011;
ROM[13421] <= 32'b00000000011100010010000000100011;
ROM[13422] <= 32'b00000000010000010000000100010011;
ROM[13423] <= 32'b00000110110000000000001110010011;
ROM[13424] <= 32'b00000000011100010010000000100011;
ROM[13425] <= 32'b00000000010000010000000100010011;
ROM[13426] <= 32'b00000110011000000000001110010011;
ROM[13427] <= 32'b00000000011100010010000000100011;
ROM[13428] <= 32'b00000000010000010000000100010011;
ROM[13429] <= 32'b00001110011000000000001110010011;
ROM[13430] <= 32'b00000000011100010010000000100011;
ROM[13431] <= 32'b00000000010000010000000100010011;
ROM[13432] <= 32'b00000000000000000000001110010011;
ROM[13433] <= 32'b00000000011100010010000000100011;
ROM[13434] <= 32'b00000000010000010000000100010011;
ROM[13435] <= 32'b00000000000000001101001110110111;
ROM[13436] <= 32'b00100011100000111000001110010011;
ROM[13437] <= 32'b00000000111000111000001110110011;
ROM[13438] <= 32'b00000000011100010010000000100011;
ROM[13439] <= 32'b00000000010000010000000100010011;
ROM[13440] <= 32'b00000000001100010010000000100011;
ROM[13441] <= 32'b00000000010000010000000100010011;
ROM[13442] <= 32'b00000000010000010010000000100011;
ROM[13443] <= 32'b00000000010000010000000100010011;
ROM[13444] <= 32'b00000000010100010010000000100011;
ROM[13445] <= 32'b00000000010000010000000100010011;
ROM[13446] <= 32'b00000000011000010010000000100011;
ROM[13447] <= 32'b00000000010000010000000100010011;
ROM[13448] <= 32'b00000001010000000000001110010011;
ROM[13449] <= 32'b00000010010000111000001110010011;
ROM[13450] <= 32'b01000000011100010000001110110011;
ROM[13451] <= 32'b00000000011100000000001000110011;
ROM[13452] <= 32'b00000000001000000000000110110011;
ROM[13453] <= 32'b00100000010000000010000011101111;
ROM[13454] <= 32'b11111111110000010000000100010011;
ROM[13455] <= 32'b00000000000000010010001110000011;
ROM[13456] <= 32'b00000000011101100010000000100011;
ROM[13457] <= 32'b00000101001100000000001110010011;
ROM[13458] <= 32'b00000000011100010010000000100011;
ROM[13459] <= 32'b00000000010000010000000100010011;
ROM[13460] <= 32'b00000111100000000000001110010011;
ROM[13461] <= 32'b00000000011100010010000000100011;
ROM[13462] <= 32'b00000000010000010000000100010011;
ROM[13463] <= 32'b00001100110000000000001110010011;
ROM[13464] <= 32'b00000000011100010010000000100011;
ROM[13465] <= 32'b00000000010000010000000100010011;
ROM[13466] <= 32'b00001110000000000000001110010011;
ROM[13467] <= 32'b00000000011100010010000000100011;
ROM[13468] <= 32'b00000000010000010000000100010011;
ROM[13469] <= 32'b00000111000000000000001110010011;
ROM[13470] <= 32'b00000000011100010010000000100011;
ROM[13471] <= 32'b00000000010000010000000100010011;
ROM[13472] <= 32'b00000001110000000000001110010011;
ROM[13473] <= 32'b00000000011100010010000000100011;
ROM[13474] <= 32'b00000000010000010000000100010011;
ROM[13475] <= 32'b00001100110000000000001110010011;
ROM[13476] <= 32'b00000000011100010010000000100011;
ROM[13477] <= 32'b00000000010000010000000100010011;
ROM[13478] <= 32'b00000111100000000000001110010011;
ROM[13479] <= 32'b00000000011100010010000000100011;
ROM[13480] <= 32'b00000000010000010000000100010011;
ROM[13481] <= 32'b00000000000000000000001110010011;
ROM[13482] <= 32'b00000000011100010010000000100011;
ROM[13483] <= 32'b00000000010000010000000100010011;
ROM[13484] <= 32'b00000000000000001101001110110111;
ROM[13485] <= 32'b00101111110000111000001110010011;
ROM[13486] <= 32'b00000000111000111000001110110011;
ROM[13487] <= 32'b00000000011100010010000000100011;
ROM[13488] <= 32'b00000000010000010000000100010011;
ROM[13489] <= 32'b00000000001100010010000000100011;
ROM[13490] <= 32'b00000000010000010000000100010011;
ROM[13491] <= 32'b00000000010000010010000000100011;
ROM[13492] <= 32'b00000000010000010000000100010011;
ROM[13493] <= 32'b00000000010100010010000000100011;
ROM[13494] <= 32'b00000000010000010000000100010011;
ROM[13495] <= 32'b00000000011000010010000000100011;
ROM[13496] <= 32'b00000000010000010000000100010011;
ROM[13497] <= 32'b00000001010000000000001110010011;
ROM[13498] <= 32'b00000010010000111000001110010011;
ROM[13499] <= 32'b01000000011100010000001110110011;
ROM[13500] <= 32'b00000000011100000000001000110011;
ROM[13501] <= 32'b00000000001000000000000110110011;
ROM[13502] <= 32'b00010100000000000010000011101111;
ROM[13503] <= 32'b11111111110000010000000100010011;
ROM[13504] <= 32'b00000000000000010010001110000011;
ROM[13505] <= 32'b00000000011101100010000000100011;
ROM[13506] <= 32'b00000101010000000000001110010011;
ROM[13507] <= 32'b00000000011100010010000000100011;
ROM[13508] <= 32'b00000000010000010000000100010011;
ROM[13509] <= 32'b00001111110000000000001110010011;
ROM[13510] <= 32'b00000000011100010010000000100011;
ROM[13511] <= 32'b00000000010000010000000100010011;
ROM[13512] <= 32'b00001011010000000000001110010011;
ROM[13513] <= 32'b00000000011100010010000000100011;
ROM[13514] <= 32'b00000000010000010000000100010011;
ROM[13515] <= 32'b00000011000000000000001110010011;
ROM[13516] <= 32'b00000000011100010010000000100011;
ROM[13517] <= 32'b00000000010000010000000100010011;
ROM[13518] <= 32'b00000011000000000000001110010011;
ROM[13519] <= 32'b00000000011100010010000000100011;
ROM[13520] <= 32'b00000000010000010000000100010011;
ROM[13521] <= 32'b00000011000000000000001110010011;
ROM[13522] <= 32'b00000000011100010010000000100011;
ROM[13523] <= 32'b00000000010000010000000100010011;
ROM[13524] <= 32'b00000011000000000000001110010011;
ROM[13525] <= 32'b00000000011100010010000000100011;
ROM[13526] <= 32'b00000000010000010000000100010011;
ROM[13527] <= 32'b00000111100000000000001110010011;
ROM[13528] <= 32'b00000000011100010010000000100011;
ROM[13529] <= 32'b00000000010000010000000100010011;
ROM[13530] <= 32'b00000000000000000000001110010011;
ROM[13531] <= 32'b00000000011100010010000000100011;
ROM[13532] <= 32'b00000000010000010000000100010011;
ROM[13533] <= 32'b00000000000000001101001110110111;
ROM[13534] <= 32'b00111100000000111000001110010011;
ROM[13535] <= 32'b00000000111000111000001110110011;
ROM[13536] <= 32'b00000000011100010010000000100011;
ROM[13537] <= 32'b00000000010000010000000100010011;
ROM[13538] <= 32'b00000000001100010010000000100011;
ROM[13539] <= 32'b00000000010000010000000100010011;
ROM[13540] <= 32'b00000000010000010010000000100011;
ROM[13541] <= 32'b00000000010000010000000100010011;
ROM[13542] <= 32'b00000000010100010010000000100011;
ROM[13543] <= 32'b00000000010000010000000100010011;
ROM[13544] <= 32'b00000000011000010010000000100011;
ROM[13545] <= 32'b00000000010000010000000100010011;
ROM[13546] <= 32'b00000001010000000000001110010011;
ROM[13547] <= 32'b00000010010000111000001110010011;
ROM[13548] <= 32'b01000000011100010000001110110011;
ROM[13549] <= 32'b00000000011100000000001000110011;
ROM[13550] <= 32'b00000000001000000000000110110011;
ROM[13551] <= 32'b00000111110000000010000011101111;
ROM[13552] <= 32'b11111111110000010000000100010011;
ROM[13553] <= 32'b00000000000000010010001110000011;
ROM[13554] <= 32'b00000000011101100010000000100011;
ROM[13555] <= 32'b00000101010100000000001110010011;
ROM[13556] <= 32'b00000000011100010010000000100011;
ROM[13557] <= 32'b00000000010000010000000100010011;
ROM[13558] <= 32'b00001100110000000000001110010011;
ROM[13559] <= 32'b00000000011100010010000000100011;
ROM[13560] <= 32'b00000000010000010000000100010011;
ROM[13561] <= 32'b00001100110000000000001110010011;
ROM[13562] <= 32'b00000000011100010010000000100011;
ROM[13563] <= 32'b00000000010000010000000100010011;
ROM[13564] <= 32'b00001100110000000000001110010011;
ROM[13565] <= 32'b00000000011100010010000000100011;
ROM[13566] <= 32'b00000000010000010000000100010011;
ROM[13567] <= 32'b00001100110000000000001110010011;
ROM[13568] <= 32'b00000000011100010010000000100011;
ROM[13569] <= 32'b00000000010000010000000100010011;
ROM[13570] <= 32'b00001100110000000000001110010011;
ROM[13571] <= 32'b00000000011100010010000000100011;
ROM[13572] <= 32'b00000000010000010000000100010011;
ROM[13573] <= 32'b00001100110000000000001110010011;
ROM[13574] <= 32'b00000000011100010010000000100011;
ROM[13575] <= 32'b00000000010000010000000100010011;
ROM[13576] <= 32'b00001111110000000000001110010011;
ROM[13577] <= 32'b00000000011100010010000000100011;
ROM[13578] <= 32'b00000000010000010000000100010011;
ROM[13579] <= 32'b00000000000000000000001110010011;
ROM[13580] <= 32'b00000000011100010010000000100011;
ROM[13581] <= 32'b00000000010000010000000100010011;
ROM[13582] <= 32'b00000000000000001101001110110111;
ROM[13583] <= 32'b01001000010000111000001110010011;
ROM[13584] <= 32'b00000000111000111000001110110011;
ROM[13585] <= 32'b00000000011100010010000000100011;
ROM[13586] <= 32'b00000000010000010000000100010011;
ROM[13587] <= 32'b00000000001100010010000000100011;
ROM[13588] <= 32'b00000000010000010000000100010011;
ROM[13589] <= 32'b00000000010000010010000000100011;
ROM[13590] <= 32'b00000000010000010000000100010011;
ROM[13591] <= 32'b00000000010100010010000000100011;
ROM[13592] <= 32'b00000000010000010000000100010011;
ROM[13593] <= 32'b00000000011000010010000000100011;
ROM[13594] <= 32'b00000000010000010000000100010011;
ROM[13595] <= 32'b00000001010000000000001110010011;
ROM[13596] <= 32'b00000010010000111000001110010011;
ROM[13597] <= 32'b01000000011100010000001110110011;
ROM[13598] <= 32'b00000000011100000000001000110011;
ROM[13599] <= 32'b00000000001000000000000110110011;
ROM[13600] <= 32'b01111011100100000001000011101111;
ROM[13601] <= 32'b11111111110000010000000100010011;
ROM[13602] <= 32'b00000000000000010010001110000011;
ROM[13603] <= 32'b00000000011101100010000000100011;
ROM[13604] <= 32'b00000101011000000000001110010011;
ROM[13605] <= 32'b00000000011100010010000000100011;
ROM[13606] <= 32'b00000000010000010000000100010011;
ROM[13607] <= 32'b00001100110000000000001110010011;
ROM[13608] <= 32'b00000000011100010010000000100011;
ROM[13609] <= 32'b00000000010000010000000100010011;
ROM[13610] <= 32'b00001100110000000000001110010011;
ROM[13611] <= 32'b00000000011100010010000000100011;
ROM[13612] <= 32'b00000000010000010000000100010011;
ROM[13613] <= 32'b00001100110000000000001110010011;
ROM[13614] <= 32'b00000000011100010010000000100011;
ROM[13615] <= 32'b00000000010000010000000100010011;
ROM[13616] <= 32'b00001100110000000000001110010011;
ROM[13617] <= 32'b00000000011100010010000000100011;
ROM[13618] <= 32'b00000000010000010000000100010011;
ROM[13619] <= 32'b00001100110000000000001110010011;
ROM[13620] <= 32'b00000000011100010010000000100011;
ROM[13621] <= 32'b00000000010000010000000100010011;
ROM[13622] <= 32'b00000111100000000000001110010011;
ROM[13623] <= 32'b00000000011100010010000000100011;
ROM[13624] <= 32'b00000000010000010000000100010011;
ROM[13625] <= 32'b00000011000000000000001110010011;
ROM[13626] <= 32'b00000000011100010010000000100011;
ROM[13627] <= 32'b00000000010000010000000100010011;
ROM[13628] <= 32'b00000000000000000000001110010011;
ROM[13629] <= 32'b00000000011100010010000000100011;
ROM[13630] <= 32'b00000000010000010000000100010011;
ROM[13631] <= 32'b00000000000000001101001110110111;
ROM[13632] <= 32'b01010100100000111000001110010011;
ROM[13633] <= 32'b00000000111000111000001110110011;
ROM[13634] <= 32'b00000000011100010010000000100011;
ROM[13635] <= 32'b00000000010000010000000100010011;
ROM[13636] <= 32'b00000000001100010010000000100011;
ROM[13637] <= 32'b00000000010000010000000100010011;
ROM[13638] <= 32'b00000000010000010010000000100011;
ROM[13639] <= 32'b00000000010000010000000100010011;
ROM[13640] <= 32'b00000000010100010010000000100011;
ROM[13641] <= 32'b00000000010000010000000100010011;
ROM[13642] <= 32'b00000000011000010010000000100011;
ROM[13643] <= 32'b00000000010000010000000100010011;
ROM[13644] <= 32'b00000001010000000000001110010011;
ROM[13645] <= 32'b00000010010000111000001110010011;
ROM[13646] <= 32'b01000000011100010000001110110011;
ROM[13647] <= 32'b00000000011100000000001000110011;
ROM[13648] <= 32'b00000000001000000000000110110011;
ROM[13649] <= 32'b01101111010100000001000011101111;
ROM[13650] <= 32'b11111111110000010000000100010011;
ROM[13651] <= 32'b00000000000000010010001110000011;
ROM[13652] <= 32'b00000000011101100010000000100011;
ROM[13653] <= 32'b00000101011100000000001110010011;
ROM[13654] <= 32'b00000000011100010010000000100011;
ROM[13655] <= 32'b00000000010000010000000100010011;
ROM[13656] <= 32'b00001100011000000000001110010011;
ROM[13657] <= 32'b00000000011100010010000000100011;
ROM[13658] <= 32'b00000000010000010000000100010011;
ROM[13659] <= 32'b00001100011000000000001110010011;
ROM[13660] <= 32'b00000000011100010010000000100011;
ROM[13661] <= 32'b00000000010000010000000100010011;
ROM[13662] <= 32'b00001100011000000000001110010011;
ROM[13663] <= 32'b00000000011100010010000000100011;
ROM[13664] <= 32'b00000000010000010000000100010011;
ROM[13665] <= 32'b00001101011000000000001110010011;
ROM[13666] <= 32'b00000000011100010010000000100011;
ROM[13667] <= 32'b00000000010000010000000100010011;
ROM[13668] <= 32'b00001111111000000000001110010011;
ROM[13669] <= 32'b00000000011100010010000000100011;
ROM[13670] <= 32'b00000000010000010000000100010011;
ROM[13671] <= 32'b00001110111000000000001110010011;
ROM[13672] <= 32'b00000000011100010010000000100011;
ROM[13673] <= 32'b00000000010000010000000100010011;
ROM[13674] <= 32'b00001100011000000000001110010011;
ROM[13675] <= 32'b00000000011100010010000000100011;
ROM[13676] <= 32'b00000000010000010000000100010011;
ROM[13677] <= 32'b00000000000000000000001110010011;
ROM[13678] <= 32'b00000000011100010010000000100011;
ROM[13679] <= 32'b00000000010000010000000100010011;
ROM[13680] <= 32'b00000000000000001101001110110111;
ROM[13681] <= 32'b01100000110000111000001110010011;
ROM[13682] <= 32'b00000000111000111000001110110011;
ROM[13683] <= 32'b00000000011100010010000000100011;
ROM[13684] <= 32'b00000000010000010000000100010011;
ROM[13685] <= 32'b00000000001100010010000000100011;
ROM[13686] <= 32'b00000000010000010000000100010011;
ROM[13687] <= 32'b00000000010000010010000000100011;
ROM[13688] <= 32'b00000000010000010000000100010011;
ROM[13689] <= 32'b00000000010100010010000000100011;
ROM[13690] <= 32'b00000000010000010000000100010011;
ROM[13691] <= 32'b00000000011000010010000000100011;
ROM[13692] <= 32'b00000000010000010000000100010011;
ROM[13693] <= 32'b00000001010000000000001110010011;
ROM[13694] <= 32'b00000010010000111000001110010011;
ROM[13695] <= 32'b01000000011100010000001110110011;
ROM[13696] <= 32'b00000000011100000000001000110011;
ROM[13697] <= 32'b00000000001000000000000110110011;
ROM[13698] <= 32'b01100011000100000001000011101111;
ROM[13699] <= 32'b11111111110000010000000100010011;
ROM[13700] <= 32'b00000000000000010010001110000011;
ROM[13701] <= 32'b00000000011101100010000000100011;
ROM[13702] <= 32'b00000101100000000000001110010011;
ROM[13703] <= 32'b00000000011100010010000000100011;
ROM[13704] <= 32'b00000000010000010000000100010011;
ROM[13705] <= 32'b00001100011000000000001110010011;
ROM[13706] <= 32'b00000000011100010010000000100011;
ROM[13707] <= 32'b00000000010000010000000100010011;
ROM[13708] <= 32'b00001100011000000000001110010011;
ROM[13709] <= 32'b00000000011100010010000000100011;
ROM[13710] <= 32'b00000000010000010000000100010011;
ROM[13711] <= 32'b00000110110000000000001110010011;
ROM[13712] <= 32'b00000000011100010010000000100011;
ROM[13713] <= 32'b00000000010000010000000100010011;
ROM[13714] <= 32'b00000011100000000000001110010011;
ROM[13715] <= 32'b00000000011100010010000000100011;
ROM[13716] <= 32'b00000000010000010000000100010011;
ROM[13717] <= 32'b00000011100000000000001110010011;
ROM[13718] <= 32'b00000000011100010010000000100011;
ROM[13719] <= 32'b00000000010000010000000100010011;
ROM[13720] <= 32'b00000110110000000000001110010011;
ROM[13721] <= 32'b00000000011100010010000000100011;
ROM[13722] <= 32'b00000000010000010000000100010011;
ROM[13723] <= 32'b00001100011000000000001110010011;
ROM[13724] <= 32'b00000000011100010010000000100011;
ROM[13725] <= 32'b00000000010000010000000100010011;
ROM[13726] <= 32'b00000000000000000000001110010011;
ROM[13727] <= 32'b00000000011100010010000000100011;
ROM[13728] <= 32'b00000000010000010000000100010011;
ROM[13729] <= 32'b00000000000000001101001110110111;
ROM[13730] <= 32'b01101101000000111000001110010011;
ROM[13731] <= 32'b00000000111000111000001110110011;
ROM[13732] <= 32'b00000000011100010010000000100011;
ROM[13733] <= 32'b00000000010000010000000100010011;
ROM[13734] <= 32'b00000000001100010010000000100011;
ROM[13735] <= 32'b00000000010000010000000100010011;
ROM[13736] <= 32'b00000000010000010010000000100011;
ROM[13737] <= 32'b00000000010000010000000100010011;
ROM[13738] <= 32'b00000000010100010010000000100011;
ROM[13739] <= 32'b00000000010000010000000100010011;
ROM[13740] <= 32'b00000000011000010010000000100011;
ROM[13741] <= 32'b00000000010000010000000100010011;
ROM[13742] <= 32'b00000001010000000000001110010011;
ROM[13743] <= 32'b00000010010000111000001110010011;
ROM[13744] <= 32'b01000000011100010000001110110011;
ROM[13745] <= 32'b00000000011100000000001000110011;
ROM[13746] <= 32'b00000000001000000000000110110011;
ROM[13747] <= 32'b01010110110100000001000011101111;
ROM[13748] <= 32'b11111111110000010000000100010011;
ROM[13749] <= 32'b00000000000000010010001110000011;
ROM[13750] <= 32'b00000000011101100010000000100011;
ROM[13751] <= 32'b00000101100100000000001110010011;
ROM[13752] <= 32'b00000000011100010010000000100011;
ROM[13753] <= 32'b00000000010000010000000100010011;
ROM[13754] <= 32'b00001100110000000000001110010011;
ROM[13755] <= 32'b00000000011100010010000000100011;
ROM[13756] <= 32'b00000000010000010000000100010011;
ROM[13757] <= 32'b00001100110000000000001110010011;
ROM[13758] <= 32'b00000000011100010010000000100011;
ROM[13759] <= 32'b00000000010000010000000100010011;
ROM[13760] <= 32'b00001100110000000000001110010011;
ROM[13761] <= 32'b00000000011100010010000000100011;
ROM[13762] <= 32'b00000000010000010000000100010011;
ROM[13763] <= 32'b00000111100000000000001110010011;
ROM[13764] <= 32'b00000000011100010010000000100011;
ROM[13765] <= 32'b00000000010000010000000100010011;
ROM[13766] <= 32'b00000011000000000000001110010011;
ROM[13767] <= 32'b00000000011100010010000000100011;
ROM[13768] <= 32'b00000000010000010000000100010011;
ROM[13769] <= 32'b00000011000000000000001110010011;
ROM[13770] <= 32'b00000000011100010010000000100011;
ROM[13771] <= 32'b00000000010000010000000100010011;
ROM[13772] <= 32'b00000111100000000000001110010011;
ROM[13773] <= 32'b00000000011100010010000000100011;
ROM[13774] <= 32'b00000000010000010000000100010011;
ROM[13775] <= 32'b00000000000000000000001110010011;
ROM[13776] <= 32'b00000000011100010010000000100011;
ROM[13777] <= 32'b00000000010000010000000100010011;
ROM[13778] <= 32'b00000000000000001101001110110111;
ROM[13779] <= 32'b01111001010000111000001110010011;
ROM[13780] <= 32'b00000000111000111000001110110011;
ROM[13781] <= 32'b00000000011100010010000000100011;
ROM[13782] <= 32'b00000000010000010000000100010011;
ROM[13783] <= 32'b00000000001100010010000000100011;
ROM[13784] <= 32'b00000000010000010000000100010011;
ROM[13785] <= 32'b00000000010000010010000000100011;
ROM[13786] <= 32'b00000000010000010000000100010011;
ROM[13787] <= 32'b00000000010100010010000000100011;
ROM[13788] <= 32'b00000000010000010000000100010011;
ROM[13789] <= 32'b00000000011000010010000000100011;
ROM[13790] <= 32'b00000000010000010000000100010011;
ROM[13791] <= 32'b00000001010000000000001110010011;
ROM[13792] <= 32'b00000010010000111000001110010011;
ROM[13793] <= 32'b01000000011100010000001110110011;
ROM[13794] <= 32'b00000000011100000000001000110011;
ROM[13795] <= 32'b00000000001000000000000110110011;
ROM[13796] <= 32'b01001010100100000001000011101111;
ROM[13797] <= 32'b11111111110000010000000100010011;
ROM[13798] <= 32'b00000000000000010010001110000011;
ROM[13799] <= 32'b00000000011101100010000000100011;
ROM[13800] <= 32'b00000101101000000000001110010011;
ROM[13801] <= 32'b00000000011100010010000000100011;
ROM[13802] <= 32'b00000000010000010000000100010011;
ROM[13803] <= 32'b00001111111000000000001110010011;
ROM[13804] <= 32'b00000000011100010010000000100011;
ROM[13805] <= 32'b00000000010000010000000100010011;
ROM[13806] <= 32'b00001100011000000000001110010011;
ROM[13807] <= 32'b00000000011100010010000000100011;
ROM[13808] <= 32'b00000000010000010000000100010011;
ROM[13809] <= 32'b00001000110000000000001110010011;
ROM[13810] <= 32'b00000000011100010010000000100011;
ROM[13811] <= 32'b00000000010000010000000100010011;
ROM[13812] <= 32'b00000001100000000000001110010011;
ROM[13813] <= 32'b00000000011100010010000000100011;
ROM[13814] <= 32'b00000000010000010000000100010011;
ROM[13815] <= 32'b00000011001000000000001110010011;
ROM[13816] <= 32'b00000000011100010010000000100011;
ROM[13817] <= 32'b00000000010000010000000100010011;
ROM[13818] <= 32'b00000110011000000000001110010011;
ROM[13819] <= 32'b00000000011100010010000000100011;
ROM[13820] <= 32'b00000000010000010000000100010011;
ROM[13821] <= 32'b00001111111000000000001110010011;
ROM[13822] <= 32'b00000000011100010010000000100011;
ROM[13823] <= 32'b00000000010000010000000100010011;
ROM[13824] <= 32'b00000000000000000000001110010011;
ROM[13825] <= 32'b00000000011100010010000000100011;
ROM[13826] <= 32'b00000000010000010000000100010011;
ROM[13827] <= 32'b00000000000000001110001110110111;
ROM[13828] <= 32'b10000101100000111000001110010011;
ROM[13829] <= 32'b00000000111000111000001110110011;
ROM[13830] <= 32'b00000000011100010010000000100011;
ROM[13831] <= 32'b00000000010000010000000100010011;
ROM[13832] <= 32'b00000000001100010010000000100011;
ROM[13833] <= 32'b00000000010000010000000100010011;
ROM[13834] <= 32'b00000000010000010010000000100011;
ROM[13835] <= 32'b00000000010000010000000100010011;
ROM[13836] <= 32'b00000000010100010010000000100011;
ROM[13837] <= 32'b00000000010000010000000100010011;
ROM[13838] <= 32'b00000000011000010010000000100011;
ROM[13839] <= 32'b00000000010000010000000100010011;
ROM[13840] <= 32'b00000001010000000000001110010011;
ROM[13841] <= 32'b00000010010000111000001110010011;
ROM[13842] <= 32'b01000000011100010000001110110011;
ROM[13843] <= 32'b00000000011100000000001000110011;
ROM[13844] <= 32'b00000000001000000000000110110011;
ROM[13845] <= 32'b00111110010100000001000011101111;
ROM[13846] <= 32'b11111111110000010000000100010011;
ROM[13847] <= 32'b00000000000000010010001110000011;
ROM[13848] <= 32'b00000000011101100010000000100011;
ROM[13849] <= 32'b00000101101100000000001110010011;
ROM[13850] <= 32'b00000000011100010010000000100011;
ROM[13851] <= 32'b00000000010000010000000100010011;
ROM[13852] <= 32'b00000111100000000000001110010011;
ROM[13853] <= 32'b00000000011100010010000000100011;
ROM[13854] <= 32'b00000000010000010000000100010011;
ROM[13855] <= 32'b00000110000000000000001110010011;
ROM[13856] <= 32'b00000000011100010010000000100011;
ROM[13857] <= 32'b00000000010000010000000100010011;
ROM[13858] <= 32'b00000110000000000000001110010011;
ROM[13859] <= 32'b00000000011100010010000000100011;
ROM[13860] <= 32'b00000000010000010000000100010011;
ROM[13861] <= 32'b00000110000000000000001110010011;
ROM[13862] <= 32'b00000000011100010010000000100011;
ROM[13863] <= 32'b00000000010000010000000100010011;
ROM[13864] <= 32'b00000110000000000000001110010011;
ROM[13865] <= 32'b00000000011100010010000000100011;
ROM[13866] <= 32'b00000000010000010000000100010011;
ROM[13867] <= 32'b00000110000000000000001110010011;
ROM[13868] <= 32'b00000000011100010010000000100011;
ROM[13869] <= 32'b00000000010000010000000100010011;
ROM[13870] <= 32'b00000111100000000000001110010011;
ROM[13871] <= 32'b00000000011100010010000000100011;
ROM[13872] <= 32'b00000000010000010000000100010011;
ROM[13873] <= 32'b00000000000000000000001110010011;
ROM[13874] <= 32'b00000000011100010010000000100011;
ROM[13875] <= 32'b00000000010000010000000100010011;
ROM[13876] <= 32'b00000000000000001110001110110111;
ROM[13877] <= 32'b10010001110000111000001110010011;
ROM[13878] <= 32'b00000000111000111000001110110011;
ROM[13879] <= 32'b00000000011100010010000000100011;
ROM[13880] <= 32'b00000000010000010000000100010011;
ROM[13881] <= 32'b00000000001100010010000000100011;
ROM[13882] <= 32'b00000000010000010000000100010011;
ROM[13883] <= 32'b00000000010000010010000000100011;
ROM[13884] <= 32'b00000000010000010000000100010011;
ROM[13885] <= 32'b00000000010100010010000000100011;
ROM[13886] <= 32'b00000000010000010000000100010011;
ROM[13887] <= 32'b00000000011000010010000000100011;
ROM[13888] <= 32'b00000000010000010000000100010011;
ROM[13889] <= 32'b00000001010000000000001110010011;
ROM[13890] <= 32'b00000010010000111000001110010011;
ROM[13891] <= 32'b01000000011100010000001110110011;
ROM[13892] <= 32'b00000000011100000000001000110011;
ROM[13893] <= 32'b00000000001000000000000110110011;
ROM[13894] <= 32'b00110010000100000001000011101111;
ROM[13895] <= 32'b11111111110000010000000100010011;
ROM[13896] <= 32'b00000000000000010010001110000011;
ROM[13897] <= 32'b00000000011101100010000000100011;
ROM[13898] <= 32'b00000101110000000000001110010011;
ROM[13899] <= 32'b00000000011100010010000000100011;
ROM[13900] <= 32'b00000000010000010000000100010011;
ROM[13901] <= 32'b00001100000000000000001110010011;
ROM[13902] <= 32'b00000000011100010010000000100011;
ROM[13903] <= 32'b00000000010000010000000100010011;
ROM[13904] <= 32'b00000110000000000000001110010011;
ROM[13905] <= 32'b00000000011100010010000000100011;
ROM[13906] <= 32'b00000000010000010000000100010011;
ROM[13907] <= 32'b00000011000000000000001110010011;
ROM[13908] <= 32'b00000000011100010010000000100011;
ROM[13909] <= 32'b00000000010000010000000100010011;
ROM[13910] <= 32'b00000001100000000000001110010011;
ROM[13911] <= 32'b00000000011100010010000000100011;
ROM[13912] <= 32'b00000000010000010000000100010011;
ROM[13913] <= 32'b00000000110000000000001110010011;
ROM[13914] <= 32'b00000000011100010010000000100011;
ROM[13915] <= 32'b00000000010000010000000100010011;
ROM[13916] <= 32'b00000000011000000000001110010011;
ROM[13917] <= 32'b00000000011100010010000000100011;
ROM[13918] <= 32'b00000000010000010000000100010011;
ROM[13919] <= 32'b00000000001000000000001110010011;
ROM[13920] <= 32'b00000000011100010010000000100011;
ROM[13921] <= 32'b00000000010000010000000100010011;
ROM[13922] <= 32'b00000000000000000000001110010011;
ROM[13923] <= 32'b00000000011100010010000000100011;
ROM[13924] <= 32'b00000000010000010000000100010011;
ROM[13925] <= 32'b00000000000000001110001110110111;
ROM[13926] <= 32'b10011110000000111000001110010011;
ROM[13927] <= 32'b00000000111000111000001110110011;
ROM[13928] <= 32'b00000000011100010010000000100011;
ROM[13929] <= 32'b00000000010000010000000100010011;
ROM[13930] <= 32'b00000000001100010010000000100011;
ROM[13931] <= 32'b00000000010000010000000100010011;
ROM[13932] <= 32'b00000000010000010010000000100011;
ROM[13933] <= 32'b00000000010000010000000100010011;
ROM[13934] <= 32'b00000000010100010010000000100011;
ROM[13935] <= 32'b00000000010000010000000100010011;
ROM[13936] <= 32'b00000000011000010010000000100011;
ROM[13937] <= 32'b00000000010000010000000100010011;
ROM[13938] <= 32'b00000001010000000000001110010011;
ROM[13939] <= 32'b00000010010000111000001110010011;
ROM[13940] <= 32'b01000000011100010000001110110011;
ROM[13941] <= 32'b00000000011100000000001000110011;
ROM[13942] <= 32'b00000000001000000000000110110011;
ROM[13943] <= 32'b00100101110100000001000011101111;
ROM[13944] <= 32'b11111111110000010000000100010011;
ROM[13945] <= 32'b00000000000000010010001110000011;
ROM[13946] <= 32'b00000000011101100010000000100011;
ROM[13947] <= 32'b00000101110100000000001110010011;
ROM[13948] <= 32'b00000000011100010010000000100011;
ROM[13949] <= 32'b00000000010000010000000100010011;
ROM[13950] <= 32'b00000111100000000000001110010011;
ROM[13951] <= 32'b00000000011100010010000000100011;
ROM[13952] <= 32'b00000000010000010000000100010011;
ROM[13953] <= 32'b00000001100000000000001110010011;
ROM[13954] <= 32'b00000000011100010010000000100011;
ROM[13955] <= 32'b00000000010000010000000100010011;
ROM[13956] <= 32'b00000001100000000000001110010011;
ROM[13957] <= 32'b00000000011100010010000000100011;
ROM[13958] <= 32'b00000000010000010000000100010011;
ROM[13959] <= 32'b00000001100000000000001110010011;
ROM[13960] <= 32'b00000000011100010010000000100011;
ROM[13961] <= 32'b00000000010000010000000100010011;
ROM[13962] <= 32'b00000001100000000000001110010011;
ROM[13963] <= 32'b00000000011100010010000000100011;
ROM[13964] <= 32'b00000000010000010000000100010011;
ROM[13965] <= 32'b00000001100000000000001110010011;
ROM[13966] <= 32'b00000000011100010010000000100011;
ROM[13967] <= 32'b00000000010000010000000100010011;
ROM[13968] <= 32'b00000111100000000000001110010011;
ROM[13969] <= 32'b00000000011100010010000000100011;
ROM[13970] <= 32'b00000000010000010000000100010011;
ROM[13971] <= 32'b00000000000000000000001110010011;
ROM[13972] <= 32'b00000000011100010010000000100011;
ROM[13973] <= 32'b00000000010000010000000100010011;
ROM[13974] <= 32'b00000000000000001110001110110111;
ROM[13975] <= 32'b10101010010000111000001110010011;
ROM[13976] <= 32'b00000000111000111000001110110011;
ROM[13977] <= 32'b00000000011100010010000000100011;
ROM[13978] <= 32'b00000000010000010000000100010011;
ROM[13979] <= 32'b00000000001100010010000000100011;
ROM[13980] <= 32'b00000000010000010000000100010011;
ROM[13981] <= 32'b00000000010000010010000000100011;
ROM[13982] <= 32'b00000000010000010000000100010011;
ROM[13983] <= 32'b00000000010100010010000000100011;
ROM[13984] <= 32'b00000000010000010000000100010011;
ROM[13985] <= 32'b00000000011000010010000000100011;
ROM[13986] <= 32'b00000000010000010000000100010011;
ROM[13987] <= 32'b00000001010000000000001110010011;
ROM[13988] <= 32'b00000010010000111000001110010011;
ROM[13989] <= 32'b01000000011100010000001110110011;
ROM[13990] <= 32'b00000000011100000000001000110011;
ROM[13991] <= 32'b00000000001000000000000110110011;
ROM[13992] <= 32'b00011001100100000001000011101111;
ROM[13993] <= 32'b11111111110000010000000100010011;
ROM[13994] <= 32'b00000000000000010010001110000011;
ROM[13995] <= 32'b00000000011101100010000000100011;
ROM[13996] <= 32'b00000101111000000000001110010011;
ROM[13997] <= 32'b00000000011100010010000000100011;
ROM[13998] <= 32'b00000000010000010000000100010011;
ROM[13999] <= 32'b00000001000000000000001110010011;
ROM[14000] <= 32'b00000000011100010010000000100011;
ROM[14001] <= 32'b00000000010000010000000100010011;
ROM[14002] <= 32'b00000011100000000000001110010011;
ROM[14003] <= 32'b00000000011100010010000000100011;
ROM[14004] <= 32'b00000000010000010000000100010011;
ROM[14005] <= 32'b00000110110000000000001110010011;
ROM[14006] <= 32'b00000000011100010010000000100011;
ROM[14007] <= 32'b00000000010000010000000100010011;
ROM[14008] <= 32'b00001100011000000000001110010011;
ROM[14009] <= 32'b00000000011100010010000000100011;
ROM[14010] <= 32'b00000000010000010000000100010011;
ROM[14011] <= 32'b00000000000000000000001110010011;
ROM[14012] <= 32'b00000000011100010010000000100011;
ROM[14013] <= 32'b00000000010000010000000100010011;
ROM[14014] <= 32'b00000000000000000000001110010011;
ROM[14015] <= 32'b00000000011100010010000000100011;
ROM[14016] <= 32'b00000000010000010000000100010011;
ROM[14017] <= 32'b00000000000000000000001110010011;
ROM[14018] <= 32'b00000000011100010010000000100011;
ROM[14019] <= 32'b00000000010000010000000100010011;
ROM[14020] <= 32'b00000000000000000000001110010011;
ROM[14021] <= 32'b00000000011100010010000000100011;
ROM[14022] <= 32'b00000000010000010000000100010011;
ROM[14023] <= 32'b00000000000000001110001110110111;
ROM[14024] <= 32'b10110110100000111000001110010011;
ROM[14025] <= 32'b00000000111000111000001110110011;
ROM[14026] <= 32'b00000000011100010010000000100011;
ROM[14027] <= 32'b00000000010000010000000100010011;
ROM[14028] <= 32'b00000000001100010010000000100011;
ROM[14029] <= 32'b00000000010000010000000100010011;
ROM[14030] <= 32'b00000000010000010010000000100011;
ROM[14031] <= 32'b00000000010000010000000100010011;
ROM[14032] <= 32'b00000000010100010010000000100011;
ROM[14033] <= 32'b00000000010000010000000100010011;
ROM[14034] <= 32'b00000000011000010010000000100011;
ROM[14035] <= 32'b00000000010000010000000100010011;
ROM[14036] <= 32'b00000001010000000000001110010011;
ROM[14037] <= 32'b00000010010000111000001110010011;
ROM[14038] <= 32'b01000000011100010000001110110011;
ROM[14039] <= 32'b00000000011100000000001000110011;
ROM[14040] <= 32'b00000000001000000000000110110011;
ROM[14041] <= 32'b00001101010100000001000011101111;
ROM[14042] <= 32'b11111111110000010000000100010011;
ROM[14043] <= 32'b00000000000000010010001110000011;
ROM[14044] <= 32'b00000000011101100010000000100011;
ROM[14045] <= 32'b00000101111100000000001110010011;
ROM[14046] <= 32'b00000000011100010010000000100011;
ROM[14047] <= 32'b00000000010000010000000100010011;
ROM[14048] <= 32'b00000000000000000000001110010011;
ROM[14049] <= 32'b00000000011100010010000000100011;
ROM[14050] <= 32'b00000000010000010000000100010011;
ROM[14051] <= 32'b00000000000000000000001110010011;
ROM[14052] <= 32'b00000000011100010010000000100011;
ROM[14053] <= 32'b00000000010000010000000100010011;
ROM[14054] <= 32'b00000000000000000000001110010011;
ROM[14055] <= 32'b00000000011100010010000000100011;
ROM[14056] <= 32'b00000000010000010000000100010011;
ROM[14057] <= 32'b00000000000000000000001110010011;
ROM[14058] <= 32'b00000000011100010010000000100011;
ROM[14059] <= 32'b00000000010000010000000100010011;
ROM[14060] <= 32'b00000000000000000000001110010011;
ROM[14061] <= 32'b00000000011100010010000000100011;
ROM[14062] <= 32'b00000000010000010000000100010011;
ROM[14063] <= 32'b00000000000000000000001110010011;
ROM[14064] <= 32'b00000000011100010010000000100011;
ROM[14065] <= 32'b00000000010000010000000100010011;
ROM[14066] <= 32'b00000000000000000000001110010011;
ROM[14067] <= 32'b00000000011100010010000000100011;
ROM[14068] <= 32'b00000000010000010000000100010011;
ROM[14069] <= 32'b00001111111100000000001110010011;
ROM[14070] <= 32'b00000000011100010010000000100011;
ROM[14071] <= 32'b00000000010000010000000100010011;
ROM[14072] <= 32'b00000000000000001110001110110111;
ROM[14073] <= 32'b11000010110000111000001110010011;
ROM[14074] <= 32'b00000000111000111000001110110011;
ROM[14075] <= 32'b00000000011100010010000000100011;
ROM[14076] <= 32'b00000000010000010000000100010011;
ROM[14077] <= 32'b00000000001100010010000000100011;
ROM[14078] <= 32'b00000000010000010000000100010011;
ROM[14079] <= 32'b00000000010000010010000000100011;
ROM[14080] <= 32'b00000000010000010000000100010011;
ROM[14081] <= 32'b00000000010100010010000000100011;
ROM[14082] <= 32'b00000000010000010000000100010011;
ROM[14083] <= 32'b00000000011000010010000000100011;
ROM[14084] <= 32'b00000000010000010000000100010011;
ROM[14085] <= 32'b00000001010000000000001110010011;
ROM[14086] <= 32'b00000010010000111000001110010011;
ROM[14087] <= 32'b01000000011100010000001110110011;
ROM[14088] <= 32'b00000000011100000000001000110011;
ROM[14089] <= 32'b00000000001000000000000110110011;
ROM[14090] <= 32'b00000001000100000001000011101111;
ROM[14091] <= 32'b11111111110000010000000100010011;
ROM[14092] <= 32'b00000000000000010010001110000011;
ROM[14093] <= 32'b00000000011101100010000000100011;
ROM[14094] <= 32'b00000110000000000000001110010011;
ROM[14095] <= 32'b00000000011100010010000000100011;
ROM[14096] <= 32'b00000000010000010000000100010011;
ROM[14097] <= 32'b00000011000000000000001110010011;
ROM[14098] <= 32'b00000000011100010010000000100011;
ROM[14099] <= 32'b00000000010000010000000100010011;
ROM[14100] <= 32'b00000011000000000000001110010011;
ROM[14101] <= 32'b00000000011100010010000000100011;
ROM[14102] <= 32'b00000000010000010000000100010011;
ROM[14103] <= 32'b00000001100000000000001110010011;
ROM[14104] <= 32'b00000000011100010010000000100011;
ROM[14105] <= 32'b00000000010000010000000100010011;
ROM[14106] <= 32'b00000000000000000000001110010011;
ROM[14107] <= 32'b00000000011100010010000000100011;
ROM[14108] <= 32'b00000000010000010000000100010011;
ROM[14109] <= 32'b00000000000000000000001110010011;
ROM[14110] <= 32'b00000000011100010010000000100011;
ROM[14111] <= 32'b00000000010000010000000100010011;
ROM[14112] <= 32'b00000000000000000000001110010011;
ROM[14113] <= 32'b00000000011100010010000000100011;
ROM[14114] <= 32'b00000000010000010000000100010011;
ROM[14115] <= 32'b00000000000000000000001110010011;
ROM[14116] <= 32'b00000000011100010010000000100011;
ROM[14117] <= 32'b00000000010000010000000100010011;
ROM[14118] <= 32'b00000000000000000000001110010011;
ROM[14119] <= 32'b00000000011100010010000000100011;
ROM[14120] <= 32'b00000000010000010000000100010011;
ROM[14121] <= 32'b00000000000000001110001110110111;
ROM[14122] <= 32'b11001111000000111000001110010011;
ROM[14123] <= 32'b00000000111000111000001110110011;
ROM[14124] <= 32'b00000000011100010010000000100011;
ROM[14125] <= 32'b00000000010000010000000100010011;
ROM[14126] <= 32'b00000000001100010010000000100011;
ROM[14127] <= 32'b00000000010000010000000100010011;
ROM[14128] <= 32'b00000000010000010010000000100011;
ROM[14129] <= 32'b00000000010000010000000100010011;
ROM[14130] <= 32'b00000000010100010010000000100011;
ROM[14131] <= 32'b00000000010000010000000100010011;
ROM[14132] <= 32'b00000000011000010010000000100011;
ROM[14133] <= 32'b00000000010000010000000100010011;
ROM[14134] <= 32'b00000001010000000000001110010011;
ROM[14135] <= 32'b00000010010000111000001110010011;
ROM[14136] <= 32'b01000000011100010000001110110011;
ROM[14137] <= 32'b00000000011100000000001000110011;
ROM[14138] <= 32'b00000000001000000000000110110011;
ROM[14139] <= 32'b01110100110000000001000011101111;
ROM[14140] <= 32'b11111111110000010000000100010011;
ROM[14141] <= 32'b00000000000000010010001110000011;
ROM[14142] <= 32'b00000000011101100010000000100011;
ROM[14143] <= 32'b00000110000100000000001110010011;
ROM[14144] <= 32'b00000000011100010010000000100011;
ROM[14145] <= 32'b00000000010000010000000100010011;
ROM[14146] <= 32'b00000000000000000000001110010011;
ROM[14147] <= 32'b00000000011100010010000000100011;
ROM[14148] <= 32'b00000000010000010000000100010011;
ROM[14149] <= 32'b00000000000000000000001110010011;
ROM[14150] <= 32'b00000000011100010010000000100011;
ROM[14151] <= 32'b00000000010000010000000100010011;
ROM[14152] <= 32'b00000111100000000000001110010011;
ROM[14153] <= 32'b00000000011100010010000000100011;
ROM[14154] <= 32'b00000000010000010000000100010011;
ROM[14155] <= 32'b00000000110000000000001110010011;
ROM[14156] <= 32'b00000000011100010010000000100011;
ROM[14157] <= 32'b00000000010000010000000100010011;
ROM[14158] <= 32'b00000111110000000000001110010011;
ROM[14159] <= 32'b00000000011100010010000000100011;
ROM[14160] <= 32'b00000000010000010000000100010011;
ROM[14161] <= 32'b00001100110000000000001110010011;
ROM[14162] <= 32'b00000000011100010010000000100011;
ROM[14163] <= 32'b00000000010000010000000100010011;
ROM[14164] <= 32'b00000111011000000000001110010011;
ROM[14165] <= 32'b00000000011100010010000000100011;
ROM[14166] <= 32'b00000000010000010000000100010011;
ROM[14167] <= 32'b00000000000000000000001110010011;
ROM[14168] <= 32'b00000000011100010010000000100011;
ROM[14169] <= 32'b00000000010000010000000100010011;
ROM[14170] <= 32'b00000000000000001110001110110111;
ROM[14171] <= 32'b11011011010000111000001110010011;
ROM[14172] <= 32'b00000000111000111000001110110011;
ROM[14173] <= 32'b00000000011100010010000000100011;
ROM[14174] <= 32'b00000000010000010000000100010011;
ROM[14175] <= 32'b00000000001100010010000000100011;
ROM[14176] <= 32'b00000000010000010000000100010011;
ROM[14177] <= 32'b00000000010000010010000000100011;
ROM[14178] <= 32'b00000000010000010000000100010011;
ROM[14179] <= 32'b00000000010100010010000000100011;
ROM[14180] <= 32'b00000000010000010000000100010011;
ROM[14181] <= 32'b00000000011000010010000000100011;
ROM[14182] <= 32'b00000000010000010000000100010011;
ROM[14183] <= 32'b00000001010000000000001110010011;
ROM[14184] <= 32'b00000010010000111000001110010011;
ROM[14185] <= 32'b01000000011100010000001110110011;
ROM[14186] <= 32'b00000000011100000000001000110011;
ROM[14187] <= 32'b00000000001000000000000110110011;
ROM[14188] <= 32'b01101000100000000001000011101111;
ROM[14189] <= 32'b11111111110000010000000100010011;
ROM[14190] <= 32'b00000000000000010010001110000011;
ROM[14191] <= 32'b00000000011101100010000000100011;
ROM[14192] <= 32'b00000110001000000000001110010011;
ROM[14193] <= 32'b00000000011100010010000000100011;
ROM[14194] <= 32'b00000000010000010000000100010011;
ROM[14195] <= 32'b00001110000000000000001110010011;
ROM[14196] <= 32'b00000000011100010010000000100011;
ROM[14197] <= 32'b00000000010000010000000100010011;
ROM[14198] <= 32'b00000110000000000000001110010011;
ROM[14199] <= 32'b00000000011100010010000000100011;
ROM[14200] <= 32'b00000000010000010000000100010011;
ROM[14201] <= 32'b00000110000000000000001110010011;
ROM[14202] <= 32'b00000000011100010010000000100011;
ROM[14203] <= 32'b00000000010000010000000100010011;
ROM[14204] <= 32'b00000111110000000000001110010011;
ROM[14205] <= 32'b00000000011100010010000000100011;
ROM[14206] <= 32'b00000000010000010000000100010011;
ROM[14207] <= 32'b00000110011000000000001110010011;
ROM[14208] <= 32'b00000000011100010010000000100011;
ROM[14209] <= 32'b00000000010000010000000100010011;
ROM[14210] <= 32'b00000110011000000000001110010011;
ROM[14211] <= 32'b00000000011100010010000000100011;
ROM[14212] <= 32'b00000000010000010000000100010011;
ROM[14213] <= 32'b00001101110000000000001110010011;
ROM[14214] <= 32'b00000000011100010010000000100011;
ROM[14215] <= 32'b00000000010000010000000100010011;
ROM[14216] <= 32'b00000000000000000000001110010011;
ROM[14217] <= 32'b00000000011100010010000000100011;
ROM[14218] <= 32'b00000000010000010000000100010011;
ROM[14219] <= 32'b00000000000000001110001110110111;
ROM[14220] <= 32'b11100111100000111000001110010011;
ROM[14221] <= 32'b00000000111000111000001110110011;
ROM[14222] <= 32'b00000000011100010010000000100011;
ROM[14223] <= 32'b00000000010000010000000100010011;
ROM[14224] <= 32'b00000000001100010010000000100011;
ROM[14225] <= 32'b00000000010000010000000100010011;
ROM[14226] <= 32'b00000000010000010010000000100011;
ROM[14227] <= 32'b00000000010000010000000100010011;
ROM[14228] <= 32'b00000000010100010010000000100011;
ROM[14229] <= 32'b00000000010000010000000100010011;
ROM[14230] <= 32'b00000000011000010010000000100011;
ROM[14231] <= 32'b00000000010000010000000100010011;
ROM[14232] <= 32'b00000001010000000000001110010011;
ROM[14233] <= 32'b00000010010000111000001110010011;
ROM[14234] <= 32'b01000000011100010000001110110011;
ROM[14235] <= 32'b00000000011100000000001000110011;
ROM[14236] <= 32'b00000000001000000000000110110011;
ROM[14237] <= 32'b01011100010000000001000011101111;
ROM[14238] <= 32'b11111111110000010000000100010011;
ROM[14239] <= 32'b00000000000000010010001110000011;
ROM[14240] <= 32'b00000000011101100010000000100011;
ROM[14241] <= 32'b00000110001100000000001110010011;
ROM[14242] <= 32'b00000000011100010010000000100011;
ROM[14243] <= 32'b00000000010000010000000100010011;
ROM[14244] <= 32'b00000000000000000000001110010011;
ROM[14245] <= 32'b00000000011100010010000000100011;
ROM[14246] <= 32'b00000000010000010000000100010011;
ROM[14247] <= 32'b00000000000000000000001110010011;
ROM[14248] <= 32'b00000000011100010010000000100011;
ROM[14249] <= 32'b00000000010000010000000100010011;
ROM[14250] <= 32'b00000111100000000000001110010011;
ROM[14251] <= 32'b00000000011100010010000000100011;
ROM[14252] <= 32'b00000000010000010000000100010011;
ROM[14253] <= 32'b00001100110000000000001110010011;
ROM[14254] <= 32'b00000000011100010010000000100011;
ROM[14255] <= 32'b00000000010000010000000100010011;
ROM[14256] <= 32'b00001100000000000000001110010011;
ROM[14257] <= 32'b00000000011100010010000000100011;
ROM[14258] <= 32'b00000000010000010000000100010011;
ROM[14259] <= 32'b00001100110000000000001110010011;
ROM[14260] <= 32'b00000000011100010010000000100011;
ROM[14261] <= 32'b00000000010000010000000100010011;
ROM[14262] <= 32'b00000111100000000000001110010011;
ROM[14263] <= 32'b00000000011100010010000000100011;
ROM[14264] <= 32'b00000000010000010000000100010011;
ROM[14265] <= 32'b00000000000000000000001110010011;
ROM[14266] <= 32'b00000000011100010010000000100011;
ROM[14267] <= 32'b00000000010000010000000100010011;
ROM[14268] <= 32'b00000000000000001110001110110111;
ROM[14269] <= 32'b11110011110000111000001110010011;
ROM[14270] <= 32'b00000000111000111000001110110011;
ROM[14271] <= 32'b00000000011100010010000000100011;
ROM[14272] <= 32'b00000000010000010000000100010011;
ROM[14273] <= 32'b00000000001100010010000000100011;
ROM[14274] <= 32'b00000000010000010000000100010011;
ROM[14275] <= 32'b00000000010000010010000000100011;
ROM[14276] <= 32'b00000000010000010000000100010011;
ROM[14277] <= 32'b00000000010100010010000000100011;
ROM[14278] <= 32'b00000000010000010000000100010011;
ROM[14279] <= 32'b00000000011000010010000000100011;
ROM[14280] <= 32'b00000000010000010000000100010011;
ROM[14281] <= 32'b00000001010000000000001110010011;
ROM[14282] <= 32'b00000010010000111000001110010011;
ROM[14283] <= 32'b01000000011100010000001110110011;
ROM[14284] <= 32'b00000000011100000000001000110011;
ROM[14285] <= 32'b00000000001000000000000110110011;
ROM[14286] <= 32'b01010000000000000001000011101111;
ROM[14287] <= 32'b11111111110000010000000100010011;
ROM[14288] <= 32'b00000000000000010010001110000011;
ROM[14289] <= 32'b00000000011101100010000000100011;
ROM[14290] <= 32'b00000110010000000000001110010011;
ROM[14291] <= 32'b00000000011100010010000000100011;
ROM[14292] <= 32'b00000000010000010000000100010011;
ROM[14293] <= 32'b00000001110000000000001110010011;
ROM[14294] <= 32'b00000000011100010010000000100011;
ROM[14295] <= 32'b00000000010000010000000100010011;
ROM[14296] <= 32'b00000000110000000000001110010011;
ROM[14297] <= 32'b00000000011100010010000000100011;
ROM[14298] <= 32'b00000000010000010000000100010011;
ROM[14299] <= 32'b00000000110000000000001110010011;
ROM[14300] <= 32'b00000000011100010010000000100011;
ROM[14301] <= 32'b00000000010000010000000100010011;
ROM[14302] <= 32'b00000111110000000000001110010011;
ROM[14303] <= 32'b00000000011100010010000000100011;
ROM[14304] <= 32'b00000000010000010000000100010011;
ROM[14305] <= 32'b00001100110000000000001110010011;
ROM[14306] <= 32'b00000000011100010010000000100011;
ROM[14307] <= 32'b00000000010000010000000100010011;
ROM[14308] <= 32'b00001100110000000000001110010011;
ROM[14309] <= 32'b00000000011100010010000000100011;
ROM[14310] <= 32'b00000000010000010000000100010011;
ROM[14311] <= 32'b00000111011000000000001110010011;
ROM[14312] <= 32'b00000000011100010010000000100011;
ROM[14313] <= 32'b00000000010000010000000100010011;
ROM[14314] <= 32'b00000000000000000000001110010011;
ROM[14315] <= 32'b00000000011100010010000000100011;
ROM[14316] <= 32'b00000000010000010000000100010011;
ROM[14317] <= 32'b00000000000000001110001110110111;
ROM[14318] <= 32'b00000000000000111000001110010011;
ROM[14319] <= 32'b00000000111000111000001110110011;
ROM[14320] <= 32'b00000000011100010010000000100011;
ROM[14321] <= 32'b00000000010000010000000100010011;
ROM[14322] <= 32'b00000000001100010010000000100011;
ROM[14323] <= 32'b00000000010000010000000100010011;
ROM[14324] <= 32'b00000000010000010010000000100011;
ROM[14325] <= 32'b00000000010000010000000100010011;
ROM[14326] <= 32'b00000000010100010010000000100011;
ROM[14327] <= 32'b00000000010000010000000100010011;
ROM[14328] <= 32'b00000000011000010010000000100011;
ROM[14329] <= 32'b00000000010000010000000100010011;
ROM[14330] <= 32'b00000001010000000000001110010011;
ROM[14331] <= 32'b00000010010000111000001110010011;
ROM[14332] <= 32'b01000000011100010000001110110011;
ROM[14333] <= 32'b00000000011100000000001000110011;
ROM[14334] <= 32'b00000000001000000000000110110011;
ROM[14335] <= 32'b01000011110000000001000011101111;
ROM[14336] <= 32'b11111111110000010000000100010011;
ROM[14337] <= 32'b00000000000000010010001110000011;
ROM[14338] <= 32'b00000000011101100010000000100011;
ROM[14339] <= 32'b00000110010100000000001110010011;
ROM[14340] <= 32'b00000000011100010010000000100011;
ROM[14341] <= 32'b00000000010000010000000100010011;
ROM[14342] <= 32'b00000000000000000000001110010011;
ROM[14343] <= 32'b00000000011100010010000000100011;
ROM[14344] <= 32'b00000000010000010000000100010011;
ROM[14345] <= 32'b00000000000000000000001110010011;
ROM[14346] <= 32'b00000000011100010010000000100011;
ROM[14347] <= 32'b00000000010000010000000100010011;
ROM[14348] <= 32'b00000111100000000000001110010011;
ROM[14349] <= 32'b00000000011100010010000000100011;
ROM[14350] <= 32'b00000000010000010000000100010011;
ROM[14351] <= 32'b00001100110000000000001110010011;
ROM[14352] <= 32'b00000000011100010010000000100011;
ROM[14353] <= 32'b00000000010000010000000100010011;
ROM[14354] <= 32'b00001111110000000000001110010011;
ROM[14355] <= 32'b00000000011100010010000000100011;
ROM[14356] <= 32'b00000000010000010000000100010011;
ROM[14357] <= 32'b00001100000000000000001110010011;
ROM[14358] <= 32'b00000000011100010010000000100011;
ROM[14359] <= 32'b00000000010000010000000100010011;
ROM[14360] <= 32'b00000111100000000000001110010011;
ROM[14361] <= 32'b00000000011100010010000000100011;
ROM[14362] <= 32'b00000000010000010000000100010011;
ROM[14363] <= 32'b00000000000000000000001110010011;
ROM[14364] <= 32'b00000000011100010010000000100011;
ROM[14365] <= 32'b00000000010000010000000100010011;
ROM[14366] <= 32'b00000000000000001110001110110111;
ROM[14367] <= 32'b00001100010000111000001110010011;
ROM[14368] <= 32'b00000000111000111000001110110011;
ROM[14369] <= 32'b00000000011100010010000000100011;
ROM[14370] <= 32'b00000000010000010000000100010011;
ROM[14371] <= 32'b00000000001100010010000000100011;
ROM[14372] <= 32'b00000000010000010000000100010011;
ROM[14373] <= 32'b00000000010000010010000000100011;
ROM[14374] <= 32'b00000000010000010000000100010011;
ROM[14375] <= 32'b00000000010100010010000000100011;
ROM[14376] <= 32'b00000000010000010000000100010011;
ROM[14377] <= 32'b00000000011000010010000000100011;
ROM[14378] <= 32'b00000000010000010000000100010011;
ROM[14379] <= 32'b00000001010000000000001110010011;
ROM[14380] <= 32'b00000010010000111000001110010011;
ROM[14381] <= 32'b01000000011100010000001110110011;
ROM[14382] <= 32'b00000000011100000000001000110011;
ROM[14383] <= 32'b00000000001000000000000110110011;
ROM[14384] <= 32'b00110111100000000001000011101111;
ROM[14385] <= 32'b11111111110000010000000100010011;
ROM[14386] <= 32'b00000000000000010010001110000011;
ROM[14387] <= 32'b00000000011101100010000000100011;
ROM[14388] <= 32'b00000110011000000000001110010011;
ROM[14389] <= 32'b00000000011100010010000000100011;
ROM[14390] <= 32'b00000000010000010000000100010011;
ROM[14391] <= 32'b00000011100000000000001110010011;
ROM[14392] <= 32'b00000000011100010010000000100011;
ROM[14393] <= 32'b00000000010000010000000100010011;
ROM[14394] <= 32'b00000110110000000000001110010011;
ROM[14395] <= 32'b00000000011100010010000000100011;
ROM[14396] <= 32'b00000000010000010000000100010011;
ROM[14397] <= 32'b00000110000000000000001110010011;
ROM[14398] <= 32'b00000000011100010010000000100011;
ROM[14399] <= 32'b00000000010000010000000100010011;
ROM[14400] <= 32'b00001111000000000000001110010011;
ROM[14401] <= 32'b00000000011100010010000000100011;
ROM[14402] <= 32'b00000000010000010000000100010011;
ROM[14403] <= 32'b00000110000000000000001110010011;
ROM[14404] <= 32'b00000000011100010010000000100011;
ROM[14405] <= 32'b00000000010000010000000100010011;
ROM[14406] <= 32'b00000110000000000000001110010011;
ROM[14407] <= 32'b00000000011100010010000000100011;
ROM[14408] <= 32'b00000000010000010000000100010011;
ROM[14409] <= 32'b00001111000000000000001110010011;
ROM[14410] <= 32'b00000000011100010010000000100011;
ROM[14411] <= 32'b00000000010000010000000100010011;
ROM[14412] <= 32'b00000000000000000000001110010011;
ROM[14413] <= 32'b00000000011100010010000000100011;
ROM[14414] <= 32'b00000000010000010000000100010011;
ROM[14415] <= 32'b00000000000000001110001110110111;
ROM[14416] <= 32'b00011000100000111000001110010011;
ROM[14417] <= 32'b00000000111000111000001110110011;
ROM[14418] <= 32'b00000000011100010010000000100011;
ROM[14419] <= 32'b00000000010000010000000100010011;
ROM[14420] <= 32'b00000000001100010010000000100011;
ROM[14421] <= 32'b00000000010000010000000100010011;
ROM[14422] <= 32'b00000000010000010010000000100011;
ROM[14423] <= 32'b00000000010000010000000100010011;
ROM[14424] <= 32'b00000000010100010010000000100011;
ROM[14425] <= 32'b00000000010000010000000100010011;
ROM[14426] <= 32'b00000000011000010010000000100011;
ROM[14427] <= 32'b00000000010000010000000100010011;
ROM[14428] <= 32'b00000001010000000000001110010011;
ROM[14429] <= 32'b00000010010000111000001110010011;
ROM[14430] <= 32'b01000000011100010000001110110011;
ROM[14431] <= 32'b00000000011100000000001000110011;
ROM[14432] <= 32'b00000000001000000000000110110011;
ROM[14433] <= 32'b00101011010000000001000011101111;
ROM[14434] <= 32'b11111111110000010000000100010011;
ROM[14435] <= 32'b00000000000000010010001110000011;
ROM[14436] <= 32'b00000000011101100010000000100011;
ROM[14437] <= 32'b00000110011100000000001110010011;
ROM[14438] <= 32'b00000000011100010010000000100011;
ROM[14439] <= 32'b00000000010000010000000100010011;
ROM[14440] <= 32'b00000000000000000000001110010011;
ROM[14441] <= 32'b00000000011100010010000000100011;
ROM[14442] <= 32'b00000000010000010000000100010011;
ROM[14443] <= 32'b00000000000000000000001110010011;
ROM[14444] <= 32'b00000000011100010010000000100011;
ROM[14445] <= 32'b00000000010000010000000100010011;
ROM[14446] <= 32'b00000111011000000000001110010011;
ROM[14447] <= 32'b00000000011100010010000000100011;
ROM[14448] <= 32'b00000000010000010000000100010011;
ROM[14449] <= 32'b00001100110000000000001110010011;
ROM[14450] <= 32'b00000000011100010010000000100011;
ROM[14451] <= 32'b00000000010000010000000100010011;
ROM[14452] <= 32'b00001100110000000000001110010011;
ROM[14453] <= 32'b00000000011100010010000000100011;
ROM[14454] <= 32'b00000000010000010000000100010011;
ROM[14455] <= 32'b00000111110000000000001110010011;
ROM[14456] <= 32'b00000000011100010010000000100011;
ROM[14457] <= 32'b00000000010000010000000100010011;
ROM[14458] <= 32'b00000000110000000000001110010011;
ROM[14459] <= 32'b00000000011100010010000000100011;
ROM[14460] <= 32'b00000000010000010000000100010011;
ROM[14461] <= 32'b00001111100000000000001110010011;
ROM[14462] <= 32'b00000000011100010010000000100011;
ROM[14463] <= 32'b00000000010000010000000100010011;
ROM[14464] <= 32'b00000000000000001110001110110111;
ROM[14465] <= 32'b00100100110000111000001110010011;
ROM[14466] <= 32'b00000000111000111000001110110011;
ROM[14467] <= 32'b00000000011100010010000000100011;
ROM[14468] <= 32'b00000000010000010000000100010011;
ROM[14469] <= 32'b00000000001100010010000000100011;
ROM[14470] <= 32'b00000000010000010000000100010011;
ROM[14471] <= 32'b00000000010000010010000000100011;
ROM[14472] <= 32'b00000000010000010000000100010011;
ROM[14473] <= 32'b00000000010100010010000000100011;
ROM[14474] <= 32'b00000000010000010000000100010011;
ROM[14475] <= 32'b00000000011000010010000000100011;
ROM[14476] <= 32'b00000000010000010000000100010011;
ROM[14477] <= 32'b00000001010000000000001110010011;
ROM[14478] <= 32'b00000010010000111000001110010011;
ROM[14479] <= 32'b01000000011100010000001110110011;
ROM[14480] <= 32'b00000000011100000000001000110011;
ROM[14481] <= 32'b00000000001000000000000110110011;
ROM[14482] <= 32'b00011111000000000001000011101111;
ROM[14483] <= 32'b11111111110000010000000100010011;
ROM[14484] <= 32'b00000000000000010010001110000011;
ROM[14485] <= 32'b00000000011101100010000000100011;
ROM[14486] <= 32'b00000110100000000000001110010011;
ROM[14487] <= 32'b00000000011100010010000000100011;
ROM[14488] <= 32'b00000000010000010000000100010011;
ROM[14489] <= 32'b00001110000000000000001110010011;
ROM[14490] <= 32'b00000000011100010010000000100011;
ROM[14491] <= 32'b00000000010000010000000100010011;
ROM[14492] <= 32'b00000110000000000000001110010011;
ROM[14493] <= 32'b00000000011100010010000000100011;
ROM[14494] <= 32'b00000000010000010000000100010011;
ROM[14495] <= 32'b00000110110000000000001110010011;
ROM[14496] <= 32'b00000000011100010010000000100011;
ROM[14497] <= 32'b00000000010000010000000100010011;
ROM[14498] <= 32'b00000111011000000000001110010011;
ROM[14499] <= 32'b00000000011100010010000000100011;
ROM[14500] <= 32'b00000000010000010000000100010011;
ROM[14501] <= 32'b00000110011000000000001110010011;
ROM[14502] <= 32'b00000000011100010010000000100011;
ROM[14503] <= 32'b00000000010000010000000100010011;
ROM[14504] <= 32'b00000110011000000000001110010011;
ROM[14505] <= 32'b00000000011100010010000000100011;
ROM[14506] <= 32'b00000000010000010000000100010011;
ROM[14507] <= 32'b00001110011000000000001110010011;
ROM[14508] <= 32'b00000000011100010010000000100011;
ROM[14509] <= 32'b00000000010000010000000100010011;
ROM[14510] <= 32'b00000000000000000000001110010011;
ROM[14511] <= 32'b00000000011100010010000000100011;
ROM[14512] <= 32'b00000000010000010000000100010011;
ROM[14513] <= 32'b00000000000000001110001110110111;
ROM[14514] <= 32'b00110001000000111000001110010011;
ROM[14515] <= 32'b00000000111000111000001110110011;
ROM[14516] <= 32'b00000000011100010010000000100011;
ROM[14517] <= 32'b00000000010000010000000100010011;
ROM[14518] <= 32'b00000000001100010010000000100011;
ROM[14519] <= 32'b00000000010000010000000100010011;
ROM[14520] <= 32'b00000000010000010010000000100011;
ROM[14521] <= 32'b00000000010000010000000100010011;
ROM[14522] <= 32'b00000000010100010010000000100011;
ROM[14523] <= 32'b00000000010000010000000100010011;
ROM[14524] <= 32'b00000000011000010010000000100011;
ROM[14525] <= 32'b00000000010000010000000100010011;
ROM[14526] <= 32'b00000001010000000000001110010011;
ROM[14527] <= 32'b00000010010000111000001110010011;
ROM[14528] <= 32'b01000000011100010000001110110011;
ROM[14529] <= 32'b00000000011100000000001000110011;
ROM[14530] <= 32'b00000000001000000000000110110011;
ROM[14531] <= 32'b00010010110000000001000011101111;
ROM[14532] <= 32'b11111111110000010000000100010011;
ROM[14533] <= 32'b00000000000000010010001110000011;
ROM[14534] <= 32'b00000000011101100010000000100011;
ROM[14535] <= 32'b00000110100100000000001110010011;
ROM[14536] <= 32'b00000000011100010010000000100011;
ROM[14537] <= 32'b00000000010000010000000100010011;
ROM[14538] <= 32'b00000011000000000000001110010011;
ROM[14539] <= 32'b00000000011100010010000000100011;
ROM[14540] <= 32'b00000000010000010000000100010011;
ROM[14541] <= 32'b00000000000000000000001110010011;
ROM[14542] <= 32'b00000000011100010010000000100011;
ROM[14543] <= 32'b00000000010000010000000100010011;
ROM[14544] <= 32'b00000111000000000000001110010011;
ROM[14545] <= 32'b00000000011100010010000000100011;
ROM[14546] <= 32'b00000000010000010000000100010011;
ROM[14547] <= 32'b00000011000000000000001110010011;
ROM[14548] <= 32'b00000000011100010010000000100011;
ROM[14549] <= 32'b00000000010000010000000100010011;
ROM[14550] <= 32'b00000011000000000000001110010011;
ROM[14551] <= 32'b00000000011100010010000000100011;
ROM[14552] <= 32'b00000000010000010000000100010011;
ROM[14553] <= 32'b00000011000000000000001110010011;
ROM[14554] <= 32'b00000000011100010010000000100011;
ROM[14555] <= 32'b00000000010000010000000100010011;
ROM[14556] <= 32'b00000111100000000000001110010011;
ROM[14557] <= 32'b00000000011100010010000000100011;
ROM[14558] <= 32'b00000000010000010000000100010011;
ROM[14559] <= 32'b00000000000000000000001110010011;
ROM[14560] <= 32'b00000000011100010010000000100011;
ROM[14561] <= 32'b00000000010000010000000100010011;
ROM[14562] <= 32'b00000000000000001110001110110111;
ROM[14563] <= 32'b00111101010000111000001110010011;
ROM[14564] <= 32'b00000000111000111000001110110011;
ROM[14565] <= 32'b00000000011100010010000000100011;
ROM[14566] <= 32'b00000000010000010000000100010011;
ROM[14567] <= 32'b00000000001100010010000000100011;
ROM[14568] <= 32'b00000000010000010000000100010011;
ROM[14569] <= 32'b00000000010000010010000000100011;
ROM[14570] <= 32'b00000000010000010000000100010011;
ROM[14571] <= 32'b00000000010100010010000000100011;
ROM[14572] <= 32'b00000000010000010000000100010011;
ROM[14573] <= 32'b00000000011000010010000000100011;
ROM[14574] <= 32'b00000000010000010000000100010011;
ROM[14575] <= 32'b00000001010000000000001110010011;
ROM[14576] <= 32'b00000010010000111000001110010011;
ROM[14577] <= 32'b01000000011100010000001110110011;
ROM[14578] <= 32'b00000000011100000000001000110011;
ROM[14579] <= 32'b00000000001000000000000110110011;
ROM[14580] <= 32'b00000110100000000001000011101111;
ROM[14581] <= 32'b11111111110000010000000100010011;
ROM[14582] <= 32'b00000000000000010010001110000011;
ROM[14583] <= 32'b00000000011101100010000000100011;
ROM[14584] <= 32'b00000110101000000000001110010011;
ROM[14585] <= 32'b00000000011100010010000000100011;
ROM[14586] <= 32'b00000000010000010000000100010011;
ROM[14587] <= 32'b00000000110000000000001110010011;
ROM[14588] <= 32'b00000000011100010010000000100011;
ROM[14589] <= 32'b00000000010000010000000100010011;
ROM[14590] <= 32'b00000000000000000000001110010011;
ROM[14591] <= 32'b00000000011100010010000000100011;
ROM[14592] <= 32'b00000000010000010000000100010011;
ROM[14593] <= 32'b00000000110000000000001110010011;
ROM[14594] <= 32'b00000000011100010010000000100011;
ROM[14595] <= 32'b00000000010000010000000100010011;
ROM[14596] <= 32'b00000000110000000000001110010011;
ROM[14597] <= 32'b00000000011100010010000000100011;
ROM[14598] <= 32'b00000000010000010000000100010011;
ROM[14599] <= 32'b00000000110000000000001110010011;
ROM[14600] <= 32'b00000000011100010010000000100011;
ROM[14601] <= 32'b00000000010000010000000100010011;
ROM[14602] <= 32'b00001100110000000000001110010011;
ROM[14603] <= 32'b00000000011100010010000000100011;
ROM[14604] <= 32'b00000000010000010000000100010011;
ROM[14605] <= 32'b00001100110000000000001110010011;
ROM[14606] <= 32'b00000000011100010010000000100011;
ROM[14607] <= 32'b00000000010000010000000100010011;
ROM[14608] <= 32'b00000111100000000000001110010011;
ROM[14609] <= 32'b00000000011100010010000000100011;
ROM[14610] <= 32'b00000000010000010000000100010011;
ROM[14611] <= 32'b00000000000000001110001110110111;
ROM[14612] <= 32'b01001001100000111000001110010011;
ROM[14613] <= 32'b00000000111000111000001110110011;
ROM[14614] <= 32'b00000000011100010010000000100011;
ROM[14615] <= 32'b00000000010000010000000100010011;
ROM[14616] <= 32'b00000000001100010010000000100011;
ROM[14617] <= 32'b00000000010000010000000100010011;
ROM[14618] <= 32'b00000000010000010010000000100011;
ROM[14619] <= 32'b00000000010000010000000100010011;
ROM[14620] <= 32'b00000000010100010010000000100011;
ROM[14621] <= 32'b00000000010000010000000100010011;
ROM[14622] <= 32'b00000000011000010010000000100011;
ROM[14623] <= 32'b00000000010000010000000100010011;
ROM[14624] <= 32'b00000001010000000000001110010011;
ROM[14625] <= 32'b00000010010000111000001110010011;
ROM[14626] <= 32'b01000000011100010000001110110011;
ROM[14627] <= 32'b00000000011100000000001000110011;
ROM[14628] <= 32'b00000000001000000000000110110011;
ROM[14629] <= 32'b01111010010100000000000011101111;
ROM[14630] <= 32'b11111111110000010000000100010011;
ROM[14631] <= 32'b00000000000000010010001110000011;
ROM[14632] <= 32'b00000000011101100010000000100011;
ROM[14633] <= 32'b00000110101100000000001110010011;
ROM[14634] <= 32'b00000000011100010010000000100011;
ROM[14635] <= 32'b00000000010000010000000100010011;
ROM[14636] <= 32'b00001110000000000000001110010011;
ROM[14637] <= 32'b00000000011100010010000000100011;
ROM[14638] <= 32'b00000000010000010000000100010011;
ROM[14639] <= 32'b00000110000000000000001110010011;
ROM[14640] <= 32'b00000000011100010010000000100011;
ROM[14641] <= 32'b00000000010000010000000100010011;
ROM[14642] <= 32'b00000110011000000000001110010011;
ROM[14643] <= 32'b00000000011100010010000000100011;
ROM[14644] <= 32'b00000000010000010000000100010011;
ROM[14645] <= 32'b00000110110000000000001110010011;
ROM[14646] <= 32'b00000000011100010010000000100011;
ROM[14647] <= 32'b00000000010000010000000100010011;
ROM[14648] <= 32'b00000111100000000000001110010011;
ROM[14649] <= 32'b00000000011100010010000000100011;
ROM[14650] <= 32'b00000000010000010000000100010011;
ROM[14651] <= 32'b00000110110000000000001110010011;
ROM[14652] <= 32'b00000000011100010010000000100011;
ROM[14653] <= 32'b00000000010000010000000100010011;
ROM[14654] <= 32'b00001110011000000000001110010011;
ROM[14655] <= 32'b00000000011100010010000000100011;
ROM[14656] <= 32'b00000000010000010000000100010011;
ROM[14657] <= 32'b00000000000000000000001110010011;
ROM[14658] <= 32'b00000000011100010010000000100011;
ROM[14659] <= 32'b00000000010000010000000100010011;
ROM[14660] <= 32'b00000000000000001110001110110111;
ROM[14661] <= 32'b01010101110000111000001110010011;
ROM[14662] <= 32'b00000000111000111000001110110011;
ROM[14663] <= 32'b00000000011100010010000000100011;
ROM[14664] <= 32'b00000000010000010000000100010011;
ROM[14665] <= 32'b00000000001100010010000000100011;
ROM[14666] <= 32'b00000000010000010000000100010011;
ROM[14667] <= 32'b00000000010000010010000000100011;
ROM[14668] <= 32'b00000000010000010000000100010011;
ROM[14669] <= 32'b00000000010100010010000000100011;
ROM[14670] <= 32'b00000000010000010000000100010011;
ROM[14671] <= 32'b00000000011000010010000000100011;
ROM[14672] <= 32'b00000000010000010000000100010011;
ROM[14673] <= 32'b00000001010000000000001110010011;
ROM[14674] <= 32'b00000010010000111000001110010011;
ROM[14675] <= 32'b01000000011100010000001110110011;
ROM[14676] <= 32'b00000000011100000000001000110011;
ROM[14677] <= 32'b00000000001000000000000110110011;
ROM[14678] <= 32'b01101110000100000000000011101111;
ROM[14679] <= 32'b11111111110000010000000100010011;
ROM[14680] <= 32'b00000000000000010010001110000011;
ROM[14681] <= 32'b00000000011101100010000000100011;
ROM[14682] <= 32'b00000110110000000000001110010011;
ROM[14683] <= 32'b00000000011100010010000000100011;
ROM[14684] <= 32'b00000000010000010000000100010011;
ROM[14685] <= 32'b00000111000000000000001110010011;
ROM[14686] <= 32'b00000000011100010010000000100011;
ROM[14687] <= 32'b00000000010000010000000100010011;
ROM[14688] <= 32'b00000011000000000000001110010011;
ROM[14689] <= 32'b00000000011100010010000000100011;
ROM[14690] <= 32'b00000000010000010000000100010011;
ROM[14691] <= 32'b00000011000000000000001110010011;
ROM[14692] <= 32'b00000000011100010010000000100011;
ROM[14693] <= 32'b00000000010000010000000100010011;
ROM[14694] <= 32'b00000011000000000000001110010011;
ROM[14695] <= 32'b00000000011100010010000000100011;
ROM[14696] <= 32'b00000000010000010000000100010011;
ROM[14697] <= 32'b00000011000000000000001110010011;
ROM[14698] <= 32'b00000000011100010010000000100011;
ROM[14699] <= 32'b00000000010000010000000100010011;
ROM[14700] <= 32'b00000011000000000000001110010011;
ROM[14701] <= 32'b00000000011100010010000000100011;
ROM[14702] <= 32'b00000000010000010000000100010011;
ROM[14703] <= 32'b00000111100000000000001110010011;
ROM[14704] <= 32'b00000000011100010010000000100011;
ROM[14705] <= 32'b00000000010000010000000100010011;
ROM[14706] <= 32'b00000000000000000000001110010011;
ROM[14707] <= 32'b00000000011100010010000000100011;
ROM[14708] <= 32'b00000000010000010000000100010011;
ROM[14709] <= 32'b00000000000000001110001110110111;
ROM[14710] <= 32'b01100010000000111000001110010011;
ROM[14711] <= 32'b00000000111000111000001110110011;
ROM[14712] <= 32'b00000000011100010010000000100011;
ROM[14713] <= 32'b00000000010000010000000100010011;
ROM[14714] <= 32'b00000000001100010010000000100011;
ROM[14715] <= 32'b00000000010000010000000100010011;
ROM[14716] <= 32'b00000000010000010010000000100011;
ROM[14717] <= 32'b00000000010000010000000100010011;
ROM[14718] <= 32'b00000000010100010010000000100011;
ROM[14719] <= 32'b00000000010000010000000100010011;
ROM[14720] <= 32'b00000000011000010010000000100011;
ROM[14721] <= 32'b00000000010000010000000100010011;
ROM[14722] <= 32'b00000001010000000000001110010011;
ROM[14723] <= 32'b00000010010000111000001110010011;
ROM[14724] <= 32'b01000000011100010000001110110011;
ROM[14725] <= 32'b00000000011100000000001000110011;
ROM[14726] <= 32'b00000000001000000000000110110011;
ROM[14727] <= 32'b01100001110100000000000011101111;
ROM[14728] <= 32'b11111111110000010000000100010011;
ROM[14729] <= 32'b00000000000000010010001110000011;
ROM[14730] <= 32'b00000000011101100010000000100011;
ROM[14731] <= 32'b00000110110100000000001110010011;
ROM[14732] <= 32'b00000000011100010010000000100011;
ROM[14733] <= 32'b00000000010000010000000100010011;
ROM[14734] <= 32'b00000000000000000000001110010011;
ROM[14735] <= 32'b00000000011100010010000000100011;
ROM[14736] <= 32'b00000000010000010000000100010011;
ROM[14737] <= 32'b00000000000000000000001110010011;
ROM[14738] <= 32'b00000000011100010010000000100011;
ROM[14739] <= 32'b00000000010000010000000100010011;
ROM[14740] <= 32'b00001100110000000000001110010011;
ROM[14741] <= 32'b00000000011100010010000000100011;
ROM[14742] <= 32'b00000000010000010000000100010011;
ROM[14743] <= 32'b00001111111000000000001110010011;
ROM[14744] <= 32'b00000000011100010010000000100011;
ROM[14745] <= 32'b00000000010000010000000100010011;
ROM[14746] <= 32'b00001111111000000000001110010011;
ROM[14747] <= 32'b00000000011100010010000000100011;
ROM[14748] <= 32'b00000000010000010000000100010011;
ROM[14749] <= 32'b00001101011000000000001110010011;
ROM[14750] <= 32'b00000000011100010010000000100011;
ROM[14751] <= 32'b00000000010000010000000100010011;
ROM[14752] <= 32'b00001100011000000000001110010011;
ROM[14753] <= 32'b00000000011100010010000000100011;
ROM[14754] <= 32'b00000000010000010000000100010011;
ROM[14755] <= 32'b00000000000000000000001110010011;
ROM[14756] <= 32'b00000000011100010010000000100011;
ROM[14757] <= 32'b00000000010000010000000100010011;
ROM[14758] <= 32'b00000000000000001110001110110111;
ROM[14759] <= 32'b01101110010000111000001110010011;
ROM[14760] <= 32'b00000000111000111000001110110011;
ROM[14761] <= 32'b00000000011100010010000000100011;
ROM[14762] <= 32'b00000000010000010000000100010011;
ROM[14763] <= 32'b00000000001100010010000000100011;
ROM[14764] <= 32'b00000000010000010000000100010011;
ROM[14765] <= 32'b00000000010000010010000000100011;
ROM[14766] <= 32'b00000000010000010000000100010011;
ROM[14767] <= 32'b00000000010100010010000000100011;
ROM[14768] <= 32'b00000000010000010000000100010011;
ROM[14769] <= 32'b00000000011000010010000000100011;
ROM[14770] <= 32'b00000000010000010000000100010011;
ROM[14771] <= 32'b00000001010000000000001110010011;
ROM[14772] <= 32'b00000010010000111000001110010011;
ROM[14773] <= 32'b01000000011100010000001110110011;
ROM[14774] <= 32'b00000000011100000000001000110011;
ROM[14775] <= 32'b00000000001000000000000110110011;
ROM[14776] <= 32'b01010101100100000000000011101111;
ROM[14777] <= 32'b11111111110000010000000100010011;
ROM[14778] <= 32'b00000000000000010010001110000011;
ROM[14779] <= 32'b00000000011101100010000000100011;
ROM[14780] <= 32'b00000110111000000000001110010011;
ROM[14781] <= 32'b00000000011100010010000000100011;
ROM[14782] <= 32'b00000000010000010000000100010011;
ROM[14783] <= 32'b00000000000000000000001110010011;
ROM[14784] <= 32'b00000000011100010010000000100011;
ROM[14785] <= 32'b00000000010000010000000100010011;
ROM[14786] <= 32'b00000000000000000000001110010011;
ROM[14787] <= 32'b00000000011100010010000000100011;
ROM[14788] <= 32'b00000000010000010000000100010011;
ROM[14789] <= 32'b00001111100000000000001110010011;
ROM[14790] <= 32'b00000000011100010010000000100011;
ROM[14791] <= 32'b00000000010000010000000100010011;
ROM[14792] <= 32'b00001100110000000000001110010011;
ROM[14793] <= 32'b00000000011100010010000000100011;
ROM[14794] <= 32'b00000000010000010000000100010011;
ROM[14795] <= 32'b00001100110000000000001110010011;
ROM[14796] <= 32'b00000000011100010010000000100011;
ROM[14797] <= 32'b00000000010000010000000100010011;
ROM[14798] <= 32'b00001100110000000000001110010011;
ROM[14799] <= 32'b00000000011100010010000000100011;
ROM[14800] <= 32'b00000000010000010000000100010011;
ROM[14801] <= 32'b00001100110000000000001110010011;
ROM[14802] <= 32'b00000000011100010010000000100011;
ROM[14803] <= 32'b00000000010000010000000100010011;
ROM[14804] <= 32'b00000000000000000000001110010011;
ROM[14805] <= 32'b00000000011100010010000000100011;
ROM[14806] <= 32'b00000000010000010000000100010011;
ROM[14807] <= 32'b00000000000000001110001110110111;
ROM[14808] <= 32'b01111010100000111000001110010011;
ROM[14809] <= 32'b00000000111000111000001110110011;
ROM[14810] <= 32'b00000000011100010010000000100011;
ROM[14811] <= 32'b00000000010000010000000100010011;
ROM[14812] <= 32'b00000000001100010010000000100011;
ROM[14813] <= 32'b00000000010000010000000100010011;
ROM[14814] <= 32'b00000000010000010010000000100011;
ROM[14815] <= 32'b00000000010000010000000100010011;
ROM[14816] <= 32'b00000000010100010010000000100011;
ROM[14817] <= 32'b00000000010000010000000100010011;
ROM[14818] <= 32'b00000000011000010010000000100011;
ROM[14819] <= 32'b00000000010000010000000100010011;
ROM[14820] <= 32'b00000001010000000000001110010011;
ROM[14821] <= 32'b00000010010000111000001110010011;
ROM[14822] <= 32'b01000000011100010000001110110011;
ROM[14823] <= 32'b00000000011100000000001000110011;
ROM[14824] <= 32'b00000000001000000000000110110011;
ROM[14825] <= 32'b01001001010100000000000011101111;
ROM[14826] <= 32'b11111111110000010000000100010011;
ROM[14827] <= 32'b00000000000000010010001110000011;
ROM[14828] <= 32'b00000000011101100010000000100011;
ROM[14829] <= 32'b00000110111100000000001110010011;
ROM[14830] <= 32'b00000000011100010010000000100011;
ROM[14831] <= 32'b00000000010000010000000100010011;
ROM[14832] <= 32'b00000000000000000000001110010011;
ROM[14833] <= 32'b00000000011100010010000000100011;
ROM[14834] <= 32'b00000000010000010000000100010011;
ROM[14835] <= 32'b00000000000000000000001110010011;
ROM[14836] <= 32'b00000000011100010010000000100011;
ROM[14837] <= 32'b00000000010000010000000100010011;
ROM[14838] <= 32'b00000111100000000000001110010011;
ROM[14839] <= 32'b00000000011100010010000000100011;
ROM[14840] <= 32'b00000000010000010000000100010011;
ROM[14841] <= 32'b00001100110000000000001110010011;
ROM[14842] <= 32'b00000000011100010010000000100011;
ROM[14843] <= 32'b00000000010000010000000100010011;
ROM[14844] <= 32'b00001100110000000000001110010011;
ROM[14845] <= 32'b00000000011100010010000000100011;
ROM[14846] <= 32'b00000000010000010000000100010011;
ROM[14847] <= 32'b00001100110000000000001110010011;
ROM[14848] <= 32'b00000000011100010010000000100011;
ROM[14849] <= 32'b00000000010000010000000100010011;
ROM[14850] <= 32'b00000111100000000000001110010011;
ROM[14851] <= 32'b00000000011100010010000000100011;
ROM[14852] <= 32'b00000000010000010000000100010011;
ROM[14853] <= 32'b00000000000000000000001110010011;
ROM[14854] <= 32'b00000000011100010010000000100011;
ROM[14855] <= 32'b00000000010000010000000100010011;
ROM[14856] <= 32'b00000000000000001111001110110111;
ROM[14857] <= 32'b10000110110000111000001110010011;
ROM[14858] <= 32'b00000000111000111000001110110011;
ROM[14859] <= 32'b00000000011100010010000000100011;
ROM[14860] <= 32'b00000000010000010000000100010011;
ROM[14861] <= 32'b00000000001100010010000000100011;
ROM[14862] <= 32'b00000000010000010000000100010011;
ROM[14863] <= 32'b00000000010000010010000000100011;
ROM[14864] <= 32'b00000000010000010000000100010011;
ROM[14865] <= 32'b00000000010100010010000000100011;
ROM[14866] <= 32'b00000000010000010000000100010011;
ROM[14867] <= 32'b00000000011000010010000000100011;
ROM[14868] <= 32'b00000000010000010000000100010011;
ROM[14869] <= 32'b00000001010000000000001110010011;
ROM[14870] <= 32'b00000010010000111000001110010011;
ROM[14871] <= 32'b01000000011100010000001110110011;
ROM[14872] <= 32'b00000000011100000000001000110011;
ROM[14873] <= 32'b00000000001000000000000110110011;
ROM[14874] <= 32'b00111101000100000000000011101111;
ROM[14875] <= 32'b11111111110000010000000100010011;
ROM[14876] <= 32'b00000000000000010010001110000011;
ROM[14877] <= 32'b00000000011101100010000000100011;
ROM[14878] <= 32'b00000111000000000000001110010011;
ROM[14879] <= 32'b00000000011100010010000000100011;
ROM[14880] <= 32'b00000000010000010000000100010011;
ROM[14881] <= 32'b00000000000000000000001110010011;
ROM[14882] <= 32'b00000000011100010010000000100011;
ROM[14883] <= 32'b00000000010000010000000100010011;
ROM[14884] <= 32'b00000000000000000000001110010011;
ROM[14885] <= 32'b00000000011100010010000000100011;
ROM[14886] <= 32'b00000000010000010000000100010011;
ROM[14887] <= 32'b00001101110000000000001110010011;
ROM[14888] <= 32'b00000000011100010010000000100011;
ROM[14889] <= 32'b00000000010000010000000100010011;
ROM[14890] <= 32'b00000110011000000000001110010011;
ROM[14891] <= 32'b00000000011100010010000000100011;
ROM[14892] <= 32'b00000000010000010000000100010011;
ROM[14893] <= 32'b00000110011000000000001110010011;
ROM[14894] <= 32'b00000000011100010010000000100011;
ROM[14895] <= 32'b00000000010000010000000100010011;
ROM[14896] <= 32'b00000111110000000000001110010011;
ROM[14897] <= 32'b00000000011100010010000000100011;
ROM[14898] <= 32'b00000000010000010000000100010011;
ROM[14899] <= 32'b00000110000000000000001110010011;
ROM[14900] <= 32'b00000000011100010010000000100011;
ROM[14901] <= 32'b00000000010000010000000100010011;
ROM[14902] <= 32'b00001111000000000000001110010011;
ROM[14903] <= 32'b00000000011100010010000000100011;
ROM[14904] <= 32'b00000000010000010000000100010011;
ROM[14905] <= 32'b00000000000000001111001110110111;
ROM[14906] <= 32'b10010011000000111000001110010011;
ROM[14907] <= 32'b00000000111000111000001110110011;
ROM[14908] <= 32'b00000000011100010010000000100011;
ROM[14909] <= 32'b00000000010000010000000100010011;
ROM[14910] <= 32'b00000000001100010010000000100011;
ROM[14911] <= 32'b00000000010000010000000100010011;
ROM[14912] <= 32'b00000000010000010010000000100011;
ROM[14913] <= 32'b00000000010000010000000100010011;
ROM[14914] <= 32'b00000000010100010010000000100011;
ROM[14915] <= 32'b00000000010000010000000100010011;
ROM[14916] <= 32'b00000000011000010010000000100011;
ROM[14917] <= 32'b00000000010000010000000100010011;
ROM[14918] <= 32'b00000001010000000000001110010011;
ROM[14919] <= 32'b00000010010000111000001110010011;
ROM[14920] <= 32'b01000000011100010000001110110011;
ROM[14921] <= 32'b00000000011100000000001000110011;
ROM[14922] <= 32'b00000000001000000000000110110011;
ROM[14923] <= 32'b00110000110100000000000011101111;
ROM[14924] <= 32'b11111111110000010000000100010011;
ROM[14925] <= 32'b00000000000000010010001110000011;
ROM[14926] <= 32'b00000000011101100010000000100011;
ROM[14927] <= 32'b00000111000100000000001110010011;
ROM[14928] <= 32'b00000000011100010010000000100011;
ROM[14929] <= 32'b00000000010000010000000100010011;
ROM[14930] <= 32'b00000000000000000000001110010011;
ROM[14931] <= 32'b00000000011100010010000000100011;
ROM[14932] <= 32'b00000000010000010000000100010011;
ROM[14933] <= 32'b00000000000000000000001110010011;
ROM[14934] <= 32'b00000000011100010010000000100011;
ROM[14935] <= 32'b00000000010000010000000100010011;
ROM[14936] <= 32'b00000111011000000000001110010011;
ROM[14937] <= 32'b00000000011100010010000000100011;
ROM[14938] <= 32'b00000000010000010000000100010011;
ROM[14939] <= 32'b00001100110000000000001110010011;
ROM[14940] <= 32'b00000000011100010010000000100011;
ROM[14941] <= 32'b00000000010000010000000100010011;
ROM[14942] <= 32'b00001100110000000000001110010011;
ROM[14943] <= 32'b00000000011100010010000000100011;
ROM[14944] <= 32'b00000000010000010000000100010011;
ROM[14945] <= 32'b00000111110000000000001110010011;
ROM[14946] <= 32'b00000000011100010010000000100011;
ROM[14947] <= 32'b00000000010000010000000100010011;
ROM[14948] <= 32'b00000000110000000000001110010011;
ROM[14949] <= 32'b00000000011100010010000000100011;
ROM[14950] <= 32'b00000000010000010000000100010011;
ROM[14951] <= 32'b00000001111000000000001110010011;
ROM[14952] <= 32'b00000000011100010010000000100011;
ROM[14953] <= 32'b00000000010000010000000100010011;
ROM[14954] <= 32'b00000000000000001111001110110111;
ROM[14955] <= 32'b10011111010000111000001110010011;
ROM[14956] <= 32'b00000000111000111000001110110011;
ROM[14957] <= 32'b00000000011100010010000000100011;
ROM[14958] <= 32'b00000000010000010000000100010011;
ROM[14959] <= 32'b00000000001100010010000000100011;
ROM[14960] <= 32'b00000000010000010000000100010011;
ROM[14961] <= 32'b00000000010000010010000000100011;
ROM[14962] <= 32'b00000000010000010000000100010011;
ROM[14963] <= 32'b00000000010100010010000000100011;
ROM[14964] <= 32'b00000000010000010000000100010011;
ROM[14965] <= 32'b00000000011000010010000000100011;
ROM[14966] <= 32'b00000000010000010000000100010011;
ROM[14967] <= 32'b00000001010000000000001110010011;
ROM[14968] <= 32'b00000010010000111000001110010011;
ROM[14969] <= 32'b01000000011100010000001110110011;
ROM[14970] <= 32'b00000000011100000000001000110011;
ROM[14971] <= 32'b00000000001000000000000110110011;
ROM[14972] <= 32'b00100100100100000000000011101111;
ROM[14973] <= 32'b11111111110000010000000100010011;
ROM[14974] <= 32'b00000000000000010010001110000011;
ROM[14975] <= 32'b00000000011101100010000000100011;
ROM[14976] <= 32'b00000111001000000000001110010011;
ROM[14977] <= 32'b00000000011100010010000000100011;
ROM[14978] <= 32'b00000000010000010000000100010011;
ROM[14979] <= 32'b00000000000000000000001110010011;
ROM[14980] <= 32'b00000000011100010010000000100011;
ROM[14981] <= 32'b00000000010000010000000100010011;
ROM[14982] <= 32'b00000000000000000000001110010011;
ROM[14983] <= 32'b00000000011100010010000000100011;
ROM[14984] <= 32'b00000000010000010000000100010011;
ROM[14985] <= 32'b00001101110000000000001110010011;
ROM[14986] <= 32'b00000000011100010010000000100011;
ROM[14987] <= 32'b00000000010000010000000100010011;
ROM[14988] <= 32'b00000111011000000000001110010011;
ROM[14989] <= 32'b00000000011100010010000000100011;
ROM[14990] <= 32'b00000000010000010000000100010011;
ROM[14991] <= 32'b00000110011000000000001110010011;
ROM[14992] <= 32'b00000000011100010010000000100011;
ROM[14993] <= 32'b00000000010000010000000100010011;
ROM[14994] <= 32'b00000110000000000000001110010011;
ROM[14995] <= 32'b00000000011100010010000000100011;
ROM[14996] <= 32'b00000000010000010000000100010011;
ROM[14997] <= 32'b00001111000000000000001110010011;
ROM[14998] <= 32'b00000000011100010010000000100011;
ROM[14999] <= 32'b00000000010000010000000100010011;
ROM[15000] <= 32'b00000000000000000000001110010011;
ROM[15001] <= 32'b00000000011100010010000000100011;
ROM[15002] <= 32'b00000000010000010000000100010011;
ROM[15003] <= 32'b00000000000000001111001110110111;
ROM[15004] <= 32'b10101011100000111000001110010011;
ROM[15005] <= 32'b00000000111000111000001110110011;
ROM[15006] <= 32'b00000000011100010010000000100011;
ROM[15007] <= 32'b00000000010000010000000100010011;
ROM[15008] <= 32'b00000000001100010010000000100011;
ROM[15009] <= 32'b00000000010000010000000100010011;
ROM[15010] <= 32'b00000000010000010010000000100011;
ROM[15011] <= 32'b00000000010000010000000100010011;
ROM[15012] <= 32'b00000000010100010010000000100011;
ROM[15013] <= 32'b00000000010000010000000100010011;
ROM[15014] <= 32'b00000000011000010010000000100011;
ROM[15015] <= 32'b00000000010000010000000100010011;
ROM[15016] <= 32'b00000001010000000000001110010011;
ROM[15017] <= 32'b00000010010000111000001110010011;
ROM[15018] <= 32'b01000000011100010000001110110011;
ROM[15019] <= 32'b00000000011100000000001000110011;
ROM[15020] <= 32'b00000000001000000000000110110011;
ROM[15021] <= 32'b00011000010100000000000011101111;
ROM[15022] <= 32'b11111111110000010000000100010011;
ROM[15023] <= 32'b00000000000000010010001110000011;
ROM[15024] <= 32'b00000000011101100010000000100011;
ROM[15025] <= 32'b00000111001100000000001110010011;
ROM[15026] <= 32'b00000000011100010010000000100011;
ROM[15027] <= 32'b00000000010000010000000100010011;
ROM[15028] <= 32'b00000000000000000000001110010011;
ROM[15029] <= 32'b00000000011100010010000000100011;
ROM[15030] <= 32'b00000000010000010000000100010011;
ROM[15031] <= 32'b00000000000000000000001110010011;
ROM[15032] <= 32'b00000000011100010010000000100011;
ROM[15033] <= 32'b00000000010000010000000100010011;
ROM[15034] <= 32'b00000111110000000000001110010011;
ROM[15035] <= 32'b00000000011100010010000000100011;
ROM[15036] <= 32'b00000000010000010000000100010011;
ROM[15037] <= 32'b00001100000000000000001110010011;
ROM[15038] <= 32'b00000000011100010010000000100011;
ROM[15039] <= 32'b00000000010000010000000100010011;
ROM[15040] <= 32'b00000111100000000000001110010011;
ROM[15041] <= 32'b00000000011100010010000000100011;
ROM[15042] <= 32'b00000000010000010000000100010011;
ROM[15043] <= 32'b00000000110000000000001110010011;
ROM[15044] <= 32'b00000000011100010010000000100011;
ROM[15045] <= 32'b00000000010000010000000100010011;
ROM[15046] <= 32'b00001111100000000000001110010011;
ROM[15047] <= 32'b00000000011100010010000000100011;
ROM[15048] <= 32'b00000000010000010000000100010011;
ROM[15049] <= 32'b00000000000000000000001110010011;
ROM[15050] <= 32'b00000000011100010010000000100011;
ROM[15051] <= 32'b00000000010000010000000100010011;
ROM[15052] <= 32'b00000000000000001111001110110111;
ROM[15053] <= 32'b10110111110000111000001110010011;
ROM[15054] <= 32'b00000000111000111000001110110011;
ROM[15055] <= 32'b00000000011100010010000000100011;
ROM[15056] <= 32'b00000000010000010000000100010011;
ROM[15057] <= 32'b00000000001100010010000000100011;
ROM[15058] <= 32'b00000000010000010000000100010011;
ROM[15059] <= 32'b00000000010000010010000000100011;
ROM[15060] <= 32'b00000000010000010000000100010011;
ROM[15061] <= 32'b00000000010100010010000000100011;
ROM[15062] <= 32'b00000000010000010000000100010011;
ROM[15063] <= 32'b00000000011000010010000000100011;
ROM[15064] <= 32'b00000000010000010000000100010011;
ROM[15065] <= 32'b00000001010000000000001110010011;
ROM[15066] <= 32'b00000010010000111000001110010011;
ROM[15067] <= 32'b01000000011100010000001110110011;
ROM[15068] <= 32'b00000000011100000000001000110011;
ROM[15069] <= 32'b00000000001000000000000110110011;
ROM[15070] <= 32'b00001100000100000000000011101111;
ROM[15071] <= 32'b11111111110000010000000100010011;
ROM[15072] <= 32'b00000000000000010010001110000011;
ROM[15073] <= 32'b00000000011101100010000000100011;
ROM[15074] <= 32'b00000111010000000000001110010011;
ROM[15075] <= 32'b00000000011100010010000000100011;
ROM[15076] <= 32'b00000000010000010000000100010011;
ROM[15077] <= 32'b00000001000000000000001110010011;
ROM[15078] <= 32'b00000000011100010010000000100011;
ROM[15079] <= 32'b00000000010000010000000100010011;
ROM[15080] <= 32'b00000011000000000000001110010011;
ROM[15081] <= 32'b00000000011100010010000000100011;
ROM[15082] <= 32'b00000000010000010000000100010011;
ROM[15083] <= 32'b00000111110000000000001110010011;
ROM[15084] <= 32'b00000000011100010010000000100011;
ROM[15085] <= 32'b00000000010000010000000100010011;
ROM[15086] <= 32'b00000011000000000000001110010011;
ROM[15087] <= 32'b00000000011100010010000000100011;
ROM[15088] <= 32'b00000000010000010000000100010011;
ROM[15089] <= 32'b00000011000000000000001110010011;
ROM[15090] <= 32'b00000000011100010010000000100011;
ROM[15091] <= 32'b00000000010000010000000100010011;
ROM[15092] <= 32'b00000011010000000000001110010011;
ROM[15093] <= 32'b00000000011100010010000000100011;
ROM[15094] <= 32'b00000000010000010000000100010011;
ROM[15095] <= 32'b00000001100000000000001110010011;
ROM[15096] <= 32'b00000000011100010010000000100011;
ROM[15097] <= 32'b00000000010000010000000100010011;
ROM[15098] <= 32'b00000000000000000000001110010011;
ROM[15099] <= 32'b00000000011100010010000000100011;
ROM[15100] <= 32'b00000000010000010000000100010011;
ROM[15101] <= 32'b00000000000000001111001110110111;
ROM[15102] <= 32'b11000100000000111000001110010011;
ROM[15103] <= 32'b00000000111000111000001110110011;
ROM[15104] <= 32'b00000000011100010010000000100011;
ROM[15105] <= 32'b00000000010000010000000100010011;
ROM[15106] <= 32'b00000000001100010010000000100011;
ROM[15107] <= 32'b00000000010000010000000100010011;
ROM[15108] <= 32'b00000000010000010010000000100011;
ROM[15109] <= 32'b00000000010000010000000100010011;
ROM[15110] <= 32'b00000000010100010010000000100011;
ROM[15111] <= 32'b00000000010000010000000100010011;
ROM[15112] <= 32'b00000000011000010010000000100011;
ROM[15113] <= 32'b00000000010000010000000100010011;
ROM[15114] <= 32'b00000001010000000000001110010011;
ROM[15115] <= 32'b00000010010000111000001110010011;
ROM[15116] <= 32'b01000000011100010000001110110011;
ROM[15117] <= 32'b00000000011100000000001000110011;
ROM[15118] <= 32'b00000000001000000000000110110011;
ROM[15119] <= 32'b01111111110000000000000011101111;
ROM[15120] <= 32'b11111111110000010000000100010011;
ROM[15121] <= 32'b00000000000000010010001110000011;
ROM[15122] <= 32'b00000000011101100010000000100011;
ROM[15123] <= 32'b00000111010100000000001110010011;
ROM[15124] <= 32'b00000000011100010010000000100011;
ROM[15125] <= 32'b00000000010000010000000100010011;
ROM[15126] <= 32'b00000000000000000000001110010011;
ROM[15127] <= 32'b00000000011100010010000000100011;
ROM[15128] <= 32'b00000000010000010000000100010011;
ROM[15129] <= 32'b00000000000000000000001110010011;
ROM[15130] <= 32'b00000000011100010010000000100011;
ROM[15131] <= 32'b00000000010000010000000100010011;
ROM[15132] <= 32'b00001100110000000000001110010011;
ROM[15133] <= 32'b00000000011100010010000000100011;
ROM[15134] <= 32'b00000000010000010000000100010011;
ROM[15135] <= 32'b00001100110000000000001110010011;
ROM[15136] <= 32'b00000000011100010010000000100011;
ROM[15137] <= 32'b00000000010000010000000100010011;
ROM[15138] <= 32'b00001100110000000000001110010011;
ROM[15139] <= 32'b00000000011100010010000000100011;
ROM[15140] <= 32'b00000000010000010000000100010011;
ROM[15141] <= 32'b00001100110000000000001110010011;
ROM[15142] <= 32'b00000000011100010010000000100011;
ROM[15143] <= 32'b00000000010000010000000100010011;
ROM[15144] <= 32'b00000111011000000000001110010011;
ROM[15145] <= 32'b00000000011100010010000000100011;
ROM[15146] <= 32'b00000000010000010000000100010011;
ROM[15147] <= 32'b00000000000000000000001110010011;
ROM[15148] <= 32'b00000000011100010010000000100011;
ROM[15149] <= 32'b00000000010000010000000100010011;
ROM[15150] <= 32'b00000000000000001111001110110111;
ROM[15151] <= 32'b11010000010000111000001110010011;
ROM[15152] <= 32'b00000000111000111000001110110011;
ROM[15153] <= 32'b00000000011100010010000000100011;
ROM[15154] <= 32'b00000000010000010000000100010011;
ROM[15155] <= 32'b00000000001100010010000000100011;
ROM[15156] <= 32'b00000000010000010000000100010011;
ROM[15157] <= 32'b00000000010000010010000000100011;
ROM[15158] <= 32'b00000000010000010000000100010011;
ROM[15159] <= 32'b00000000010100010010000000100011;
ROM[15160] <= 32'b00000000010000010000000100010011;
ROM[15161] <= 32'b00000000011000010010000000100011;
ROM[15162] <= 32'b00000000010000010000000100010011;
ROM[15163] <= 32'b00000001010000000000001110010011;
ROM[15164] <= 32'b00000010010000111000001110010011;
ROM[15165] <= 32'b01000000011100010000001110110011;
ROM[15166] <= 32'b00000000011100000000001000110011;
ROM[15167] <= 32'b00000000001000000000000110110011;
ROM[15168] <= 32'b01110011100000000000000011101111;
ROM[15169] <= 32'b11111111110000010000000100010011;
ROM[15170] <= 32'b00000000000000010010001110000011;
ROM[15171] <= 32'b00000000011101100010000000100011;
ROM[15172] <= 32'b00000111011000000000001110010011;
ROM[15173] <= 32'b00000000011100010010000000100011;
ROM[15174] <= 32'b00000000010000010000000100010011;
ROM[15175] <= 32'b00000000000000000000001110010011;
ROM[15176] <= 32'b00000000011100010010000000100011;
ROM[15177] <= 32'b00000000010000010000000100010011;
ROM[15178] <= 32'b00000000000000000000001110010011;
ROM[15179] <= 32'b00000000011100010010000000100011;
ROM[15180] <= 32'b00000000010000010000000100010011;
ROM[15181] <= 32'b00001100110000000000001110010011;
ROM[15182] <= 32'b00000000011100010010000000100011;
ROM[15183] <= 32'b00000000010000010000000100010011;
ROM[15184] <= 32'b00001100110000000000001110010011;
ROM[15185] <= 32'b00000000011100010010000000100011;
ROM[15186] <= 32'b00000000010000010000000100010011;
ROM[15187] <= 32'b00001100110000000000001110010011;
ROM[15188] <= 32'b00000000011100010010000000100011;
ROM[15189] <= 32'b00000000010000010000000100010011;
ROM[15190] <= 32'b00000111100000000000001110010011;
ROM[15191] <= 32'b00000000011100010010000000100011;
ROM[15192] <= 32'b00000000010000010000000100010011;
ROM[15193] <= 32'b00000011000000000000001110010011;
ROM[15194] <= 32'b00000000011100010010000000100011;
ROM[15195] <= 32'b00000000010000010000000100010011;
ROM[15196] <= 32'b00000000000000000000001110010011;
ROM[15197] <= 32'b00000000011100010010000000100011;
ROM[15198] <= 32'b00000000010000010000000100010011;
ROM[15199] <= 32'b00000000000000001111001110110111;
ROM[15200] <= 32'b11011100100000111000001110010011;
ROM[15201] <= 32'b00000000111000111000001110110011;
ROM[15202] <= 32'b00000000011100010010000000100011;
ROM[15203] <= 32'b00000000010000010000000100010011;
ROM[15204] <= 32'b00000000001100010010000000100011;
ROM[15205] <= 32'b00000000010000010000000100010011;
ROM[15206] <= 32'b00000000010000010010000000100011;
ROM[15207] <= 32'b00000000010000010000000100010011;
ROM[15208] <= 32'b00000000010100010010000000100011;
ROM[15209] <= 32'b00000000010000010000000100010011;
ROM[15210] <= 32'b00000000011000010010000000100011;
ROM[15211] <= 32'b00000000010000010000000100010011;
ROM[15212] <= 32'b00000001010000000000001110010011;
ROM[15213] <= 32'b00000010010000111000001110010011;
ROM[15214] <= 32'b01000000011100010000001110110011;
ROM[15215] <= 32'b00000000011100000000001000110011;
ROM[15216] <= 32'b00000000001000000000000110110011;
ROM[15217] <= 32'b01100111010000000000000011101111;
ROM[15218] <= 32'b11111111110000010000000100010011;
ROM[15219] <= 32'b00000000000000010010001110000011;
ROM[15220] <= 32'b00000000011101100010000000100011;
ROM[15221] <= 32'b00000111011100000000001110010011;
ROM[15222] <= 32'b00000000011100010010000000100011;
ROM[15223] <= 32'b00000000010000010000000100010011;
ROM[15224] <= 32'b00000000000000000000001110010011;
ROM[15225] <= 32'b00000000011100010010000000100011;
ROM[15226] <= 32'b00000000010000010000000100010011;
ROM[15227] <= 32'b00000000000000000000001110010011;
ROM[15228] <= 32'b00000000011100010010000000100011;
ROM[15229] <= 32'b00000000010000010000000100010011;
ROM[15230] <= 32'b00001100011000000000001110010011;
ROM[15231] <= 32'b00000000011100010010000000100011;
ROM[15232] <= 32'b00000000010000010000000100010011;
ROM[15233] <= 32'b00001101011000000000001110010011;
ROM[15234] <= 32'b00000000011100010010000000100011;
ROM[15235] <= 32'b00000000010000010000000100010011;
ROM[15236] <= 32'b00001111111000000000001110010011;
ROM[15237] <= 32'b00000000011100010010000000100011;
ROM[15238] <= 32'b00000000010000010000000100010011;
ROM[15239] <= 32'b00001111111000000000001110010011;
ROM[15240] <= 32'b00000000011100010010000000100011;
ROM[15241] <= 32'b00000000010000010000000100010011;
ROM[15242] <= 32'b00000110110000000000001110010011;
ROM[15243] <= 32'b00000000011100010010000000100011;
ROM[15244] <= 32'b00000000010000010000000100010011;
ROM[15245] <= 32'b00000000000000000000001110010011;
ROM[15246] <= 32'b00000000011100010010000000100011;
ROM[15247] <= 32'b00000000010000010000000100010011;
ROM[15248] <= 32'b00000000000000001111001110110111;
ROM[15249] <= 32'b11101000110000111000001110010011;
ROM[15250] <= 32'b00000000111000111000001110110011;
ROM[15251] <= 32'b00000000011100010010000000100011;
ROM[15252] <= 32'b00000000010000010000000100010011;
ROM[15253] <= 32'b00000000001100010010000000100011;
ROM[15254] <= 32'b00000000010000010000000100010011;
ROM[15255] <= 32'b00000000010000010010000000100011;
ROM[15256] <= 32'b00000000010000010000000100010011;
ROM[15257] <= 32'b00000000010100010010000000100011;
ROM[15258] <= 32'b00000000010000010000000100010011;
ROM[15259] <= 32'b00000000011000010010000000100011;
ROM[15260] <= 32'b00000000010000010000000100010011;
ROM[15261] <= 32'b00000001010000000000001110010011;
ROM[15262] <= 32'b00000010010000111000001110010011;
ROM[15263] <= 32'b01000000011100010000001110110011;
ROM[15264] <= 32'b00000000011100000000001000110011;
ROM[15265] <= 32'b00000000001000000000000110110011;
ROM[15266] <= 32'b01011011000000000000000011101111;
ROM[15267] <= 32'b11111111110000010000000100010011;
ROM[15268] <= 32'b00000000000000010010001110000011;
ROM[15269] <= 32'b00000000011101100010000000100011;
ROM[15270] <= 32'b00000111100000000000001110010011;
ROM[15271] <= 32'b00000000011100010010000000100011;
ROM[15272] <= 32'b00000000010000010000000100010011;
ROM[15273] <= 32'b00000000000000000000001110010011;
ROM[15274] <= 32'b00000000011100010010000000100011;
ROM[15275] <= 32'b00000000010000010000000100010011;
ROM[15276] <= 32'b00000000000000000000001110010011;
ROM[15277] <= 32'b00000000011100010010000000100011;
ROM[15278] <= 32'b00000000010000010000000100010011;
ROM[15279] <= 32'b00001100011000000000001110010011;
ROM[15280] <= 32'b00000000011100010010000000100011;
ROM[15281] <= 32'b00000000010000010000000100010011;
ROM[15282] <= 32'b00000110110000000000001110010011;
ROM[15283] <= 32'b00000000011100010010000000100011;
ROM[15284] <= 32'b00000000010000010000000100010011;
ROM[15285] <= 32'b00000011100000000000001110010011;
ROM[15286] <= 32'b00000000011100010010000000100011;
ROM[15287] <= 32'b00000000010000010000000100010011;
ROM[15288] <= 32'b00000110110000000000001110010011;
ROM[15289] <= 32'b00000000011100010010000000100011;
ROM[15290] <= 32'b00000000010000010000000100010011;
ROM[15291] <= 32'b00001100011000000000001110010011;
ROM[15292] <= 32'b00000000011100010010000000100011;
ROM[15293] <= 32'b00000000010000010000000100010011;
ROM[15294] <= 32'b00000000000000000000001110010011;
ROM[15295] <= 32'b00000000011100010010000000100011;
ROM[15296] <= 32'b00000000010000010000000100010011;
ROM[15297] <= 32'b00000000000000001111001110110111;
ROM[15298] <= 32'b11110101000000111000001110010011;
ROM[15299] <= 32'b00000000111000111000001110110011;
ROM[15300] <= 32'b00000000011100010010000000100011;
ROM[15301] <= 32'b00000000010000010000000100010011;
ROM[15302] <= 32'b00000000001100010010000000100011;
ROM[15303] <= 32'b00000000010000010000000100010011;
ROM[15304] <= 32'b00000000010000010010000000100011;
ROM[15305] <= 32'b00000000010000010000000100010011;
ROM[15306] <= 32'b00000000010100010010000000100011;
ROM[15307] <= 32'b00000000010000010000000100010011;
ROM[15308] <= 32'b00000000011000010010000000100011;
ROM[15309] <= 32'b00000000010000010000000100010011;
ROM[15310] <= 32'b00000001010000000000001110010011;
ROM[15311] <= 32'b00000010010000111000001110010011;
ROM[15312] <= 32'b01000000011100010000001110110011;
ROM[15313] <= 32'b00000000011100000000001000110011;
ROM[15314] <= 32'b00000000001000000000000110110011;
ROM[15315] <= 32'b01001110110000000000000011101111;
ROM[15316] <= 32'b11111111110000010000000100010011;
ROM[15317] <= 32'b00000000000000010010001110000011;
ROM[15318] <= 32'b00000000011101100010000000100011;
ROM[15319] <= 32'b00000111100100000000001110010011;
ROM[15320] <= 32'b00000000011100010010000000100011;
ROM[15321] <= 32'b00000000010000010000000100010011;
ROM[15322] <= 32'b00000000000000000000001110010011;
ROM[15323] <= 32'b00000000011100010010000000100011;
ROM[15324] <= 32'b00000000010000010000000100010011;
ROM[15325] <= 32'b00000000000000000000001110010011;
ROM[15326] <= 32'b00000000011100010010000000100011;
ROM[15327] <= 32'b00000000010000010000000100010011;
ROM[15328] <= 32'b00001100110000000000001110010011;
ROM[15329] <= 32'b00000000011100010010000000100011;
ROM[15330] <= 32'b00000000010000010000000100010011;
ROM[15331] <= 32'b00001100110000000000001110010011;
ROM[15332] <= 32'b00000000011100010010000000100011;
ROM[15333] <= 32'b00000000010000010000000100010011;
ROM[15334] <= 32'b00001100110000000000001110010011;
ROM[15335] <= 32'b00000000011100010010000000100011;
ROM[15336] <= 32'b00000000010000010000000100010011;
ROM[15337] <= 32'b00000111110000000000001110010011;
ROM[15338] <= 32'b00000000011100010010000000100011;
ROM[15339] <= 32'b00000000010000010000000100010011;
ROM[15340] <= 32'b00000000110000000000001110010011;
ROM[15341] <= 32'b00000000011100010010000000100011;
ROM[15342] <= 32'b00000000010000010000000100010011;
ROM[15343] <= 32'b00001111100000000000001110010011;
ROM[15344] <= 32'b00000000011100010010000000100011;
ROM[15345] <= 32'b00000000010000010000000100010011;
ROM[15346] <= 32'b00000000000000001111001110110111;
ROM[15347] <= 32'b00000001010000111000001110010011;
ROM[15348] <= 32'b00000000111000111000001110110011;
ROM[15349] <= 32'b00000000011100010010000000100011;
ROM[15350] <= 32'b00000000010000010000000100010011;
ROM[15351] <= 32'b00000000001100010010000000100011;
ROM[15352] <= 32'b00000000010000010000000100010011;
ROM[15353] <= 32'b00000000010000010010000000100011;
ROM[15354] <= 32'b00000000010000010000000100010011;
ROM[15355] <= 32'b00000000010100010010000000100011;
ROM[15356] <= 32'b00000000010000010000000100010011;
ROM[15357] <= 32'b00000000011000010010000000100011;
ROM[15358] <= 32'b00000000010000010000000100010011;
ROM[15359] <= 32'b00000001010000000000001110010011;
ROM[15360] <= 32'b00000010010000111000001110010011;
ROM[15361] <= 32'b01000000011100010000001110110011;
ROM[15362] <= 32'b00000000011100000000001000110011;
ROM[15363] <= 32'b00000000001000000000000110110011;
ROM[15364] <= 32'b01000010100000000000000011101111;
ROM[15365] <= 32'b11111111110000010000000100010011;
ROM[15366] <= 32'b00000000000000010010001110000011;
ROM[15367] <= 32'b00000000011101100010000000100011;
ROM[15368] <= 32'b00000111101000000000001110010011;
ROM[15369] <= 32'b00000000011100010010000000100011;
ROM[15370] <= 32'b00000000010000010000000100010011;
ROM[15371] <= 32'b00000000000000000000001110010011;
ROM[15372] <= 32'b00000000011100010010000000100011;
ROM[15373] <= 32'b00000000010000010000000100010011;
ROM[15374] <= 32'b00000000000000000000001110010011;
ROM[15375] <= 32'b00000000011100010010000000100011;
ROM[15376] <= 32'b00000000010000010000000100010011;
ROM[15377] <= 32'b00001111110000000000001110010011;
ROM[15378] <= 32'b00000000011100010010000000100011;
ROM[15379] <= 32'b00000000010000010000000100010011;
ROM[15380] <= 32'b00001001100000000000001110010011;
ROM[15381] <= 32'b00000000011100010010000000100011;
ROM[15382] <= 32'b00000000010000010000000100010011;
ROM[15383] <= 32'b00000011000000000000001110010011;
ROM[15384] <= 32'b00000000011100010010000000100011;
ROM[15385] <= 32'b00000000010000010000000100010011;
ROM[15386] <= 32'b00000110010000000000001110010011;
ROM[15387] <= 32'b00000000011100010010000000100011;
ROM[15388] <= 32'b00000000010000010000000100010011;
ROM[15389] <= 32'b00001111110000000000001110010011;
ROM[15390] <= 32'b00000000011100010010000000100011;
ROM[15391] <= 32'b00000000010000010000000100010011;
ROM[15392] <= 32'b00000000000000000000001110010011;
ROM[15393] <= 32'b00000000011100010010000000100011;
ROM[15394] <= 32'b00000000010000010000000100010011;
ROM[15395] <= 32'b00000000000000001111001110110111;
ROM[15396] <= 32'b00001101100000111000001110010011;
ROM[15397] <= 32'b00000000111000111000001110110011;
ROM[15398] <= 32'b00000000011100010010000000100011;
ROM[15399] <= 32'b00000000010000010000000100010011;
ROM[15400] <= 32'b00000000001100010010000000100011;
ROM[15401] <= 32'b00000000010000010000000100010011;
ROM[15402] <= 32'b00000000010000010010000000100011;
ROM[15403] <= 32'b00000000010000010000000100010011;
ROM[15404] <= 32'b00000000010100010010000000100011;
ROM[15405] <= 32'b00000000010000010000000100010011;
ROM[15406] <= 32'b00000000011000010010000000100011;
ROM[15407] <= 32'b00000000010000010000000100010011;
ROM[15408] <= 32'b00000001010000000000001110010011;
ROM[15409] <= 32'b00000010010000111000001110010011;
ROM[15410] <= 32'b01000000011100010000001110110011;
ROM[15411] <= 32'b00000000011100000000001000110011;
ROM[15412] <= 32'b00000000001000000000000110110011;
ROM[15413] <= 32'b00110110010000000000000011101111;
ROM[15414] <= 32'b11111111110000010000000100010011;
ROM[15415] <= 32'b00000000000000010010001110000011;
ROM[15416] <= 32'b00000000011101100010000000100011;
ROM[15417] <= 32'b00000111101100000000001110010011;
ROM[15418] <= 32'b00000000011100010010000000100011;
ROM[15419] <= 32'b00000000010000010000000100010011;
ROM[15420] <= 32'b00000001110000000000001110010011;
ROM[15421] <= 32'b00000000011100010010000000100011;
ROM[15422] <= 32'b00000000010000010000000100010011;
ROM[15423] <= 32'b00000011000000000000001110010011;
ROM[15424] <= 32'b00000000011100010010000000100011;
ROM[15425] <= 32'b00000000010000010000000100010011;
ROM[15426] <= 32'b00000011000000000000001110010011;
ROM[15427] <= 32'b00000000011100010010000000100011;
ROM[15428] <= 32'b00000000010000010000000100010011;
ROM[15429] <= 32'b00001110000000000000001110010011;
ROM[15430] <= 32'b00000000011100010010000000100011;
ROM[15431] <= 32'b00000000010000010000000100010011;
ROM[15432] <= 32'b00000011000000000000001110010011;
ROM[15433] <= 32'b00000000011100010010000000100011;
ROM[15434] <= 32'b00000000010000010000000100010011;
ROM[15435] <= 32'b00000011000000000000001110010011;
ROM[15436] <= 32'b00000000011100010010000000100011;
ROM[15437] <= 32'b00000000010000010000000100010011;
ROM[15438] <= 32'b00000001110000000000001110010011;
ROM[15439] <= 32'b00000000011100010010000000100011;
ROM[15440] <= 32'b00000000010000010000000100010011;
ROM[15441] <= 32'b00000000000000000000001110010011;
ROM[15442] <= 32'b00000000011100010010000000100011;
ROM[15443] <= 32'b00000000010000010000000100010011;
ROM[15444] <= 32'b00000000000000001111001110110111;
ROM[15445] <= 32'b00011001110000111000001110010011;
ROM[15446] <= 32'b00000000111000111000001110110011;
ROM[15447] <= 32'b00000000011100010010000000100011;
ROM[15448] <= 32'b00000000010000010000000100010011;
ROM[15449] <= 32'b00000000001100010010000000100011;
ROM[15450] <= 32'b00000000010000010000000100010011;
ROM[15451] <= 32'b00000000010000010010000000100011;
ROM[15452] <= 32'b00000000010000010000000100010011;
ROM[15453] <= 32'b00000000010100010010000000100011;
ROM[15454] <= 32'b00000000010000010000000100010011;
ROM[15455] <= 32'b00000000011000010010000000100011;
ROM[15456] <= 32'b00000000010000010000000100010011;
ROM[15457] <= 32'b00000001010000000000001110010011;
ROM[15458] <= 32'b00000010010000111000001110010011;
ROM[15459] <= 32'b01000000011100010000001110110011;
ROM[15460] <= 32'b00000000011100000000001000110011;
ROM[15461] <= 32'b00000000001000000000000110110011;
ROM[15462] <= 32'b00101010000000000000000011101111;
ROM[15463] <= 32'b11111111110000010000000100010011;
ROM[15464] <= 32'b00000000000000010010001110000011;
ROM[15465] <= 32'b00000000011101100010000000100011;
ROM[15466] <= 32'b00000111110000000000001110010011;
ROM[15467] <= 32'b00000000011100010010000000100011;
ROM[15468] <= 32'b00000000010000010000000100010011;
ROM[15469] <= 32'b00000001100000000000001110010011;
ROM[15470] <= 32'b00000000011100010010000000100011;
ROM[15471] <= 32'b00000000010000010000000100010011;
ROM[15472] <= 32'b00000001100000000000001110010011;
ROM[15473] <= 32'b00000000011100010010000000100011;
ROM[15474] <= 32'b00000000010000010000000100010011;
ROM[15475] <= 32'b00000001100000000000001110010011;
ROM[15476] <= 32'b00000000011100010010000000100011;
ROM[15477] <= 32'b00000000010000010000000100010011;
ROM[15478] <= 32'b00000000000000000000001110010011;
ROM[15479] <= 32'b00000000011100010010000000100011;
ROM[15480] <= 32'b00000000010000010000000100010011;
ROM[15481] <= 32'b00000001100000000000001110010011;
ROM[15482] <= 32'b00000000011100010010000000100011;
ROM[15483] <= 32'b00000000010000010000000100010011;
ROM[15484] <= 32'b00000001100000000000001110010011;
ROM[15485] <= 32'b00000000011100010010000000100011;
ROM[15486] <= 32'b00000000010000010000000100010011;
ROM[15487] <= 32'b00000001100000000000001110010011;
ROM[15488] <= 32'b00000000011100010010000000100011;
ROM[15489] <= 32'b00000000010000010000000100010011;
ROM[15490] <= 32'b00000000000000000000001110010011;
ROM[15491] <= 32'b00000000011100010010000000100011;
ROM[15492] <= 32'b00000000010000010000000100010011;
ROM[15493] <= 32'b00000000000000001111001110110111;
ROM[15494] <= 32'b00100110000000111000001110010011;
ROM[15495] <= 32'b00000000111000111000001110110011;
ROM[15496] <= 32'b00000000011100010010000000100011;
ROM[15497] <= 32'b00000000010000010000000100010011;
ROM[15498] <= 32'b00000000001100010010000000100011;
ROM[15499] <= 32'b00000000010000010000000100010011;
ROM[15500] <= 32'b00000000010000010010000000100011;
ROM[15501] <= 32'b00000000010000010000000100010011;
ROM[15502] <= 32'b00000000010100010010000000100011;
ROM[15503] <= 32'b00000000010000010000000100010011;
ROM[15504] <= 32'b00000000011000010010000000100011;
ROM[15505] <= 32'b00000000010000010000000100010011;
ROM[15506] <= 32'b00000001010000000000001110010011;
ROM[15507] <= 32'b00000010010000111000001110010011;
ROM[15508] <= 32'b01000000011100010000001110110011;
ROM[15509] <= 32'b00000000011100000000001000110011;
ROM[15510] <= 32'b00000000001000000000000110110011;
ROM[15511] <= 32'b00011101110000000000000011101111;
ROM[15512] <= 32'b11111111110000010000000100010011;
ROM[15513] <= 32'b00000000000000010010001110000011;
ROM[15514] <= 32'b00000000011101100010000000100011;
ROM[15515] <= 32'b00000111110100000000001110010011;
ROM[15516] <= 32'b00000000011100010010000000100011;
ROM[15517] <= 32'b00000000010000010000000100010011;
ROM[15518] <= 32'b00001110000000000000001110010011;
ROM[15519] <= 32'b00000000011100010010000000100011;
ROM[15520] <= 32'b00000000010000010000000100010011;
ROM[15521] <= 32'b00000011000000000000001110010011;
ROM[15522] <= 32'b00000000011100010010000000100011;
ROM[15523] <= 32'b00000000010000010000000100010011;
ROM[15524] <= 32'b00000011000000000000001110010011;
ROM[15525] <= 32'b00000000011100010010000000100011;
ROM[15526] <= 32'b00000000010000010000000100010011;
ROM[15527] <= 32'b00000001110000000000001110010011;
ROM[15528] <= 32'b00000000011100010010000000100011;
ROM[15529] <= 32'b00000000010000010000000100010011;
ROM[15530] <= 32'b00000011000000000000001110010011;
ROM[15531] <= 32'b00000000011100010010000000100011;
ROM[15532] <= 32'b00000000010000010000000100010011;
ROM[15533] <= 32'b00000011000000000000001110010011;
ROM[15534] <= 32'b00000000011100010010000000100011;
ROM[15535] <= 32'b00000000010000010000000100010011;
ROM[15536] <= 32'b00001110000000000000001110010011;
ROM[15537] <= 32'b00000000011100010010000000100011;
ROM[15538] <= 32'b00000000010000010000000100010011;
ROM[15539] <= 32'b00000000000000000000001110010011;
ROM[15540] <= 32'b00000000011100010010000000100011;
ROM[15541] <= 32'b00000000010000010000000100010011;
ROM[15542] <= 32'b00000000000000001111001110110111;
ROM[15543] <= 32'b00110010010000111000001110010011;
ROM[15544] <= 32'b00000000111000111000001110110011;
ROM[15545] <= 32'b00000000011100010010000000100011;
ROM[15546] <= 32'b00000000010000010000000100010011;
ROM[15547] <= 32'b00000000001100010010000000100011;
ROM[15548] <= 32'b00000000010000010000000100010011;
ROM[15549] <= 32'b00000000010000010010000000100011;
ROM[15550] <= 32'b00000000010000010000000100010011;
ROM[15551] <= 32'b00000000010100010010000000100011;
ROM[15552] <= 32'b00000000010000010000000100010011;
ROM[15553] <= 32'b00000000011000010010000000100011;
ROM[15554] <= 32'b00000000010000010000000100010011;
ROM[15555] <= 32'b00000001010000000000001110010011;
ROM[15556] <= 32'b00000010010000111000001110010011;
ROM[15557] <= 32'b01000000011100010000001110110011;
ROM[15558] <= 32'b00000000011100000000001000110011;
ROM[15559] <= 32'b00000000001000000000000110110011;
ROM[15560] <= 32'b00010001100000000000000011101111;
ROM[15561] <= 32'b11111111110000010000000100010011;
ROM[15562] <= 32'b00000000000000010010001110000011;
ROM[15563] <= 32'b00000000011101100010000000100011;
ROM[15564] <= 32'b00000111111000000000001110010011;
ROM[15565] <= 32'b00000000011100010010000000100011;
ROM[15566] <= 32'b00000000010000010000000100010011;
ROM[15567] <= 32'b00000111011000000000001110010011;
ROM[15568] <= 32'b00000000011100010010000000100011;
ROM[15569] <= 32'b00000000010000010000000100010011;
ROM[15570] <= 32'b00001101110000000000001110010011;
ROM[15571] <= 32'b00000000011100010010000000100011;
ROM[15572] <= 32'b00000000010000010000000100010011;
ROM[15573] <= 32'b00000000000000000000001110010011;
ROM[15574] <= 32'b00000000011100010010000000100011;
ROM[15575] <= 32'b00000000010000010000000100010011;
ROM[15576] <= 32'b00000000000000000000001110010011;
ROM[15577] <= 32'b00000000011100010010000000100011;
ROM[15578] <= 32'b00000000010000010000000100010011;
ROM[15579] <= 32'b00000000000000000000001110010011;
ROM[15580] <= 32'b00000000011100010010000000100011;
ROM[15581] <= 32'b00000000010000010000000100010011;
ROM[15582] <= 32'b00000000000000000000001110010011;
ROM[15583] <= 32'b00000000011100010010000000100011;
ROM[15584] <= 32'b00000000010000010000000100010011;
ROM[15585] <= 32'b00000000000000000000001110010011;
ROM[15586] <= 32'b00000000011100010010000000100011;
ROM[15587] <= 32'b00000000010000010000000100010011;
ROM[15588] <= 32'b00000000000000000000001110010011;
ROM[15589] <= 32'b00000000011100010010000000100011;
ROM[15590] <= 32'b00000000010000010000000100010011;
ROM[15591] <= 32'b00000000000000001111001110110111;
ROM[15592] <= 32'b00111110100000111000001110010011;
ROM[15593] <= 32'b00000000111000111000001110110011;
ROM[15594] <= 32'b00000000011100010010000000100011;
ROM[15595] <= 32'b00000000010000010000000100010011;
ROM[15596] <= 32'b00000000001100010010000000100011;
ROM[15597] <= 32'b00000000010000010000000100010011;
ROM[15598] <= 32'b00000000010000010010000000100011;
ROM[15599] <= 32'b00000000010000010000000100010011;
ROM[15600] <= 32'b00000000010100010010000000100011;
ROM[15601] <= 32'b00000000010000010000000100010011;
ROM[15602] <= 32'b00000000011000010010000000100011;
ROM[15603] <= 32'b00000000010000010000000100010011;
ROM[15604] <= 32'b00000001010000000000001110010011;
ROM[15605] <= 32'b00000010010000111000001110010011;
ROM[15606] <= 32'b01000000011100010000001110110011;
ROM[15607] <= 32'b00000000011100000000001000110011;
ROM[15608] <= 32'b00000000001000000000000110110011;
ROM[15609] <= 32'b00000101010000000000000011101111;
ROM[15610] <= 32'b11111111110000010000000100010011;
ROM[15611] <= 32'b00000000000000010010001110000011;
ROM[15612] <= 32'b00000000011101100010000000100011;
ROM[15613] <= 32'b00000000000000000000001110010011;
ROM[15614] <= 32'b00000000011100010010000000100011;
ROM[15615] <= 32'b00000000010000010000000100010011;
ROM[15616] <= 32'b00000001010000000000001110010011;
ROM[15617] <= 32'b01000000011100011000001110110011;
ROM[15618] <= 32'b00000000000000111010000010000011;
ROM[15619] <= 32'b11111111110000010000000100010011;
ROM[15620] <= 32'b00000000000000010010001110000011;
ROM[15621] <= 32'b00000000011100100010000000100011;
ROM[15622] <= 32'b00000000010000100000000100010011;
ROM[15623] <= 32'b00000001010000000000001110010011;
ROM[15624] <= 32'b01000000011100011000001110110011;
ROM[15625] <= 32'b00000000010000111010000110000011;
ROM[15626] <= 32'b00000000100000111010001000000011;
ROM[15627] <= 32'b00000000110000111010001010000011;
ROM[15628] <= 32'b00000001000000111010001100000011;
ROM[15629] <= 32'b00000000000000001000000011100111;
ROM[15630] <= 32'b00000000000000010010000000100011;
ROM[15631] <= 32'b00000000010000010000000100010011;
ROM[15632] <= 32'b00000000100000000000001110010011;
ROM[15633] <= 32'b00000000011100010010000000100011;
ROM[15634] <= 32'b00000000010000010000000100010011;
ROM[15635] <= 32'b00000000000000001111001110110111;
ROM[15636] <= 32'b01001001100000111000001110010011;
ROM[15637] <= 32'b00000000111000111000001110110011;
ROM[15638] <= 32'b00000000011100010010000000100011;
ROM[15639] <= 32'b00000000010000010000000100010011;
ROM[15640] <= 32'b00000000001100010010000000100011;
ROM[15641] <= 32'b00000000010000010000000100010011;
ROM[15642] <= 32'b00000000010000010010000000100011;
ROM[15643] <= 32'b00000000010000010000000100010011;
ROM[15644] <= 32'b00000000010100010010000000100011;
ROM[15645] <= 32'b00000000010000010000000100010011;
ROM[15646] <= 32'b00000000011000010010000000100011;
ROM[15647] <= 32'b00000000010000010000000100010011;
ROM[15648] <= 32'b00000001010000000000001110010011;
ROM[15649] <= 32'b00000000010000111000001110010011;
ROM[15650] <= 32'b01000000011100010000001110110011;
ROM[15651] <= 32'b00000000011100000000001000110011;
ROM[15652] <= 32'b00000000001000000000000110110011;
ROM[15653] <= 32'b11111010110111110000000011101111;
ROM[15654] <= 32'b11111111110000010000000100010011;
ROM[15655] <= 32'b00000000000000010010001110000011;
ROM[15656] <= 32'b00000000011100011010000000100011;
ROM[15657] <= 32'b00000000000000100010001110000011;
ROM[15658] <= 32'b00000000011100010010000000100011;
ROM[15659] <= 32'b00000000010000010000000100010011;
ROM[15660] <= 32'b00000000010000000000001110010011;
ROM[15661] <= 32'b00000000011100010010000000100011;
ROM[15662] <= 32'b00000000010000010000000100010011;
ROM[15663] <= 32'b00000000000000001111001110110111;
ROM[15664] <= 32'b01010000100000111000001110010011;
ROM[15665] <= 32'b00000000111000111000001110110011;
ROM[15666] <= 32'b00000000011100010010000000100011;
ROM[15667] <= 32'b00000000010000010000000100010011;
ROM[15668] <= 32'b00000000001100010010000000100011;
ROM[15669] <= 32'b00000000010000010000000100010011;
ROM[15670] <= 32'b00000000010000010010000000100011;
ROM[15671] <= 32'b00000000010000010000000100010011;
ROM[15672] <= 32'b00000000010100010010000000100011;
ROM[15673] <= 32'b00000000010000010000000100010011;
ROM[15674] <= 32'b00000000011000010010000000100011;
ROM[15675] <= 32'b00000000010000010000000100010011;
ROM[15676] <= 32'b00000001010000000000001110010011;
ROM[15677] <= 32'b00000000100000111000001110010011;
ROM[15678] <= 32'b01000000011100010000001110110011;
ROM[15679] <= 32'b00000000011100000000001000110011;
ROM[15680] <= 32'b00000000001000000000000110110011;
ROM[15681] <= 32'b10111101000111111001000011101111;
ROM[15682] <= 32'b11111111110000010000000100010011;
ROM[15683] <= 32'b00000000000000010010001110000011;
ROM[15684] <= 32'b00000000011100100010000000100011;
ROM[15685] <= 32'b00000000000000100010001110000011;
ROM[15686] <= 32'b00000000011100010010000000100011;
ROM[15687] <= 32'b00000000010000010000000100010011;
ROM[15688] <= 32'b00001000100001101010001110000011;
ROM[15689] <= 32'b11111111110000010000000100010011;
ROM[15690] <= 32'b00000000000000010010010000000011;
ROM[15691] <= 32'b00000000011101000000001110110011;
ROM[15692] <= 32'b00000000011100010010000000100011;
ROM[15693] <= 32'b00000000010000010000000100010011;
ROM[15694] <= 32'b00000000000000011010001110000011;
ROM[15695] <= 32'b00000000011101100010000000100011;
ROM[15696] <= 32'b11111111110000010000000100010011;
ROM[15697] <= 32'b00000000000000010010001110000011;
ROM[15698] <= 32'b00000000000000111000001100010011;
ROM[15699] <= 32'b00000000000001100010001110000011;
ROM[15700] <= 32'b00000000110100110000010000110011;
ROM[15701] <= 32'b00000000011101000010000000100011;
ROM[15702] <= 32'b00000000000000000000001110010011;
ROM[15703] <= 32'b00000000011100010010000000100011;
ROM[15704] <= 32'b00000000010000010000000100010011;
ROM[15705] <= 32'b00000000000000011010001110000011;
ROM[15706] <= 32'b11111111110000010000000100010011;
ROM[15707] <= 32'b00000000000000010010010000000011;
ROM[15708] <= 32'b00000000011101000000001110110011;
ROM[15709] <= 32'b00000000011100010010000000100011;
ROM[15710] <= 32'b00000000010000010000000100010011;
ROM[15711] <= 32'b00000000010000100010001110000011;
ROM[15712] <= 32'b00000000011101100010000000100011;
ROM[15713] <= 32'b11111111110000010000000100010011;
ROM[15714] <= 32'b00000000000000010010001110000011;
ROM[15715] <= 32'b00000000000000111000001100010011;
ROM[15716] <= 32'b00000000000001100010001110000011;
ROM[15717] <= 32'b00000000110100110000010000110011;
ROM[15718] <= 32'b00000000011101000010000000100011;
ROM[15719] <= 32'b00000000010000000000001110010011;
ROM[15720] <= 32'b00000000011100010010000000100011;
ROM[15721] <= 32'b00000000010000010000000100010011;
ROM[15722] <= 32'b00000000000000011010001110000011;
ROM[15723] <= 32'b11111111110000010000000100010011;
ROM[15724] <= 32'b00000000000000010010010000000011;
ROM[15725] <= 32'b00000000011101000000001110110011;
ROM[15726] <= 32'b00000000011100010010000000100011;
ROM[15727] <= 32'b00000000010000010000000100010011;
ROM[15728] <= 32'b00000000100000100010001110000011;
ROM[15729] <= 32'b00000000011101100010000000100011;
ROM[15730] <= 32'b11111111110000010000000100010011;
ROM[15731] <= 32'b00000000000000010010001110000011;
ROM[15732] <= 32'b00000000000000111000001100010011;
ROM[15733] <= 32'b00000000000001100010001110000011;
ROM[15734] <= 32'b00000000110100110000010000110011;
ROM[15735] <= 32'b00000000011101000010000000100011;
ROM[15736] <= 32'b00000000100000000000001110010011;
ROM[15737] <= 32'b00000000011100010010000000100011;
ROM[15738] <= 32'b00000000010000010000000100010011;
ROM[15739] <= 32'b00000000000000011010001110000011;
ROM[15740] <= 32'b11111111110000010000000100010011;
ROM[15741] <= 32'b00000000000000010010010000000011;
ROM[15742] <= 32'b00000000011101000000001110110011;
ROM[15743] <= 32'b00000000011100010010000000100011;
ROM[15744] <= 32'b00000000010000010000000100010011;
ROM[15745] <= 32'b00000000110000100010001110000011;
ROM[15746] <= 32'b00000000011101100010000000100011;
ROM[15747] <= 32'b11111111110000010000000100010011;
ROM[15748] <= 32'b00000000000000010010001110000011;
ROM[15749] <= 32'b00000000000000111000001100010011;
ROM[15750] <= 32'b00000000000001100010001110000011;
ROM[15751] <= 32'b00000000110100110000010000110011;
ROM[15752] <= 32'b00000000011101000010000000100011;
ROM[15753] <= 32'b00000000110000000000001110010011;
ROM[15754] <= 32'b00000000011100010010000000100011;
ROM[15755] <= 32'b00000000010000010000000100010011;
ROM[15756] <= 32'b00000000000000011010001110000011;
ROM[15757] <= 32'b11111111110000010000000100010011;
ROM[15758] <= 32'b00000000000000010010010000000011;
ROM[15759] <= 32'b00000000011101000000001110110011;
ROM[15760] <= 32'b00000000011100010010000000100011;
ROM[15761] <= 32'b00000000010000010000000100010011;
ROM[15762] <= 32'b00000001000000100010001110000011;
ROM[15763] <= 32'b00000000011101100010000000100011;
ROM[15764] <= 32'b11111111110000010000000100010011;
ROM[15765] <= 32'b00000000000000010010001110000011;
ROM[15766] <= 32'b00000000000000111000001100010011;
ROM[15767] <= 32'b00000000000001100010001110000011;
ROM[15768] <= 32'b00000000110100110000010000110011;
ROM[15769] <= 32'b00000000011101000010000000100011;
ROM[15770] <= 32'b00000001000000000000001110010011;
ROM[15771] <= 32'b00000000011100010010000000100011;
ROM[15772] <= 32'b00000000010000010000000100010011;
ROM[15773] <= 32'b00000000000000011010001110000011;
ROM[15774] <= 32'b11111111110000010000000100010011;
ROM[15775] <= 32'b00000000000000010010010000000011;
ROM[15776] <= 32'b00000000011101000000001110110011;
ROM[15777] <= 32'b00000000011100010010000000100011;
ROM[15778] <= 32'b00000000010000010000000100010011;
ROM[15779] <= 32'b00000001010000100010001110000011;
ROM[15780] <= 32'b00000000011101100010000000100011;
ROM[15781] <= 32'b11111111110000010000000100010011;
ROM[15782] <= 32'b00000000000000010010001110000011;
ROM[15783] <= 32'b00000000000000111000001100010011;
ROM[15784] <= 32'b00000000000001100010001110000011;
ROM[15785] <= 32'b00000000110100110000010000110011;
ROM[15786] <= 32'b00000000011101000010000000100011;
ROM[15787] <= 32'b00000001010000000000001110010011;
ROM[15788] <= 32'b00000000011100010010000000100011;
ROM[15789] <= 32'b00000000010000010000000100010011;
ROM[15790] <= 32'b00000000000000011010001110000011;
ROM[15791] <= 32'b11111111110000010000000100010011;
ROM[15792] <= 32'b00000000000000010010010000000011;
ROM[15793] <= 32'b00000000011101000000001110110011;
ROM[15794] <= 32'b00000000011100010010000000100011;
ROM[15795] <= 32'b00000000010000010000000100010011;
ROM[15796] <= 32'b00000001100000100010001110000011;
ROM[15797] <= 32'b00000000011101100010000000100011;
ROM[15798] <= 32'b11111111110000010000000100010011;
ROM[15799] <= 32'b00000000000000010010001110000011;
ROM[15800] <= 32'b00000000000000111000001100010011;
ROM[15801] <= 32'b00000000000001100010001110000011;
ROM[15802] <= 32'b00000000110100110000010000110011;
ROM[15803] <= 32'b00000000011101000010000000100011;
ROM[15804] <= 32'b00000001100000000000001110010011;
ROM[15805] <= 32'b00000000011100010010000000100011;
ROM[15806] <= 32'b00000000010000010000000100010011;
ROM[15807] <= 32'b00000000000000011010001110000011;
ROM[15808] <= 32'b11111111110000010000000100010011;
ROM[15809] <= 32'b00000000000000010010010000000011;
ROM[15810] <= 32'b00000000011101000000001110110011;
ROM[15811] <= 32'b00000000011100010010000000100011;
ROM[15812] <= 32'b00000000010000010000000100010011;
ROM[15813] <= 32'b00000001110000100010001110000011;
ROM[15814] <= 32'b00000000011101100010000000100011;
ROM[15815] <= 32'b11111111110000010000000100010011;
ROM[15816] <= 32'b00000000000000010010001110000011;
ROM[15817] <= 32'b00000000000000111000001100010011;
ROM[15818] <= 32'b00000000000001100010001110000011;
ROM[15819] <= 32'b00000000110100110000010000110011;
ROM[15820] <= 32'b00000000011101000010000000100011;
ROM[15821] <= 32'b00000001110000000000001110010011;
ROM[15822] <= 32'b00000000011100010010000000100011;
ROM[15823] <= 32'b00000000010000010000000100010011;
ROM[15824] <= 32'b00000000000000011010001110000011;
ROM[15825] <= 32'b11111111110000010000000100010011;
ROM[15826] <= 32'b00000000000000010010010000000011;
ROM[15827] <= 32'b00000000011101000000001110110011;
ROM[15828] <= 32'b00000000011100010010000000100011;
ROM[15829] <= 32'b00000000010000010000000100010011;
ROM[15830] <= 32'b00000010000000100010001110000011;
ROM[15831] <= 32'b00000000011101100010000000100011;
ROM[15832] <= 32'b11111111110000010000000100010011;
ROM[15833] <= 32'b00000000000000010010001110000011;
ROM[15834] <= 32'b00000000000000111000001100010011;
ROM[15835] <= 32'b00000000000001100010001110000011;
ROM[15836] <= 32'b00000000110100110000010000110011;
ROM[15837] <= 32'b00000000011101000010000000100011;
ROM[15838] <= 32'b00000000000000000000001110010011;
ROM[15839] <= 32'b00000000011100010010000000100011;
ROM[15840] <= 32'b00000000010000010000000100010011;
ROM[15841] <= 32'b00000001010000000000001110010011;
ROM[15842] <= 32'b01000000011100011000001110110011;
ROM[15843] <= 32'b00000000000000111010000010000011;
ROM[15844] <= 32'b11111111110000010000000100010011;
ROM[15845] <= 32'b00000000000000010010001110000011;
ROM[15846] <= 32'b00000000011100100010000000100011;
ROM[15847] <= 32'b00000000010000100000000100010011;
ROM[15848] <= 32'b00000001010000000000001110010011;
ROM[15849] <= 32'b01000000011100011000001110110011;
ROM[15850] <= 32'b00000000010000111010000110000011;
ROM[15851] <= 32'b00000000100000111010001000000011;
ROM[15852] <= 32'b00000000110000111010001010000011;
ROM[15853] <= 32'b00000001000000111010001100000011;
ROM[15854] <= 32'b00000000000000001000000011100111;
ROM[15855] <= 32'b00000000000000010010000000100011;
ROM[15856] <= 32'b00000000010000010000000100010011;
ROM[15857] <= 32'b00000000000000100010001110000011;
ROM[15858] <= 32'b00000000011100010010000000100011;
ROM[15859] <= 32'b00000000010000010000000100010011;
ROM[15860] <= 32'b00000010000000000000001110010011;
ROM[15861] <= 32'b11111111110000010000000100010011;
ROM[15862] <= 32'b00000000000000010010010000000011;
ROM[15863] <= 32'b00000000011101000010001110110011;
ROM[15864] <= 32'b00000000011100010010000000100011;
ROM[15865] <= 32'b00000000010000010000000100010011;
ROM[15866] <= 32'b00000000000000100010001110000011;
ROM[15867] <= 32'b00000000011100010010000000100011;
ROM[15868] <= 32'b00000000010000010000000100010011;
ROM[15869] <= 32'b00000111111000000000001110010011;
ROM[15870] <= 32'b11111111110000010000000100010011;
ROM[15871] <= 32'b00000000000000010010010000000011;
ROM[15872] <= 32'b00000000100000111010001110110011;
ROM[15873] <= 32'b11111111110000010000000100010011;
ROM[15874] <= 32'b00000000000000010010010000000011;
ROM[15875] <= 32'b00000000011101000110001110110011;
ROM[15876] <= 32'b00000000000000111000101001100011;
ROM[15877] <= 32'b00000000000000010000001110110111;
ROM[15878] <= 32'b10000010100000111000001110010011;
ROM[15879] <= 32'b00000000111000111000001110110011;
ROM[15880] <= 32'b00000000000000111000000011100111;
ROM[15881] <= 32'b00000001000000000000000011101111;
ROM[15882] <= 32'b00000000000000000000001110010011;
ROM[15883] <= 32'b00000000011100100010000000100011;
ROM[15884] <= 32'b00000000010000000000000011101111;
ROM[15885] <= 32'b00000000000000100010001110000011;
ROM[15886] <= 32'b00000000011100010010000000100011;
ROM[15887] <= 32'b00000000010000010000000100010011;
ROM[15888] <= 32'b00000000000000100010001110000011;
ROM[15889] <= 32'b11111111110000010000000100010011;
ROM[15890] <= 32'b00000000000000010010010000000011;
ROM[15891] <= 32'b00000000011101000000001110110011;
ROM[15892] <= 32'b00000000011100010010000000100011;
ROM[15893] <= 32'b00000000010000010000000100010011;
ROM[15894] <= 32'b00000000000000100010001110000011;
ROM[15895] <= 32'b11111111110000010000000100010011;
ROM[15896] <= 32'b00000000000000010010010000000011;
ROM[15897] <= 32'b00000000011101000000001110110011;
ROM[15898] <= 32'b00000000011100010010000000100011;
ROM[15899] <= 32'b00000000010000010000000100010011;
ROM[15900] <= 32'b00000000000000100010001110000011;
ROM[15901] <= 32'b11111111110000010000000100010011;
ROM[15902] <= 32'b00000000000000010010010000000011;
ROM[15903] <= 32'b00000000011101000000001110110011;
ROM[15904] <= 32'b00000000011100011010000000100011;
ROM[15905] <= 32'b00000000000000011010001110000011;
ROM[15906] <= 32'b00000000011100010010000000100011;
ROM[15907] <= 32'b00000000010000010000000100010011;
ROM[15908] <= 32'b00001000100001101010001110000011;
ROM[15909] <= 32'b11111111110000010000000100010011;
ROM[15910] <= 32'b00000000000000010010010000000011;
ROM[15911] <= 32'b00000000011101000000001110110011;
ROM[15912] <= 32'b00000000000000111000001100010011;
ROM[15913] <= 32'b00000000110100110000010000110011;
ROM[15914] <= 32'b00000000000001000010001110000011;
ROM[15915] <= 32'b00000000011100010010000000100011;
ROM[15916] <= 32'b00000000010000010000000100010011;
ROM[15917] <= 32'b00000001010000000000001110010011;
ROM[15918] <= 32'b01000000011100011000001110110011;
ROM[15919] <= 32'b00000000000000111010000010000011;
ROM[15920] <= 32'b11111111110000010000000100010011;
ROM[15921] <= 32'b00000000000000010010001110000011;
ROM[15922] <= 32'b00000000011100100010000000100011;
ROM[15923] <= 32'b00000000010000100000000100010011;
ROM[15924] <= 32'b00000001010000000000001110010011;
ROM[15925] <= 32'b01000000011100011000001110110011;
ROM[15926] <= 32'b00000000010000111010000110000011;
ROM[15927] <= 32'b00000000100000111010001000000011;
ROM[15928] <= 32'b00000000110000111010001010000011;
ROM[15929] <= 32'b00000001000000111010001100000011;
ROM[15930] <= 32'b00000000000000001000000011100111;
ROM[15931] <= 32'b00000000010000100010001110000011;
ROM[15932] <= 32'b00001000011101101010000000100011;
ROM[15933] <= 32'b00000000000000100010001110000011;
ROM[15934] <= 32'b00001000011101101010001000100011;
ROM[15935] <= 32'b00000000000000000000001110010011;
ROM[15936] <= 32'b00000000011100010010000000100011;
ROM[15937] <= 32'b00000000010000010000000100010011;
ROM[15938] <= 32'b00000001010000000000001110010011;
ROM[15939] <= 32'b01000000011100011000001110110011;
ROM[15940] <= 32'b00000000000000111010000010000011;
ROM[15941] <= 32'b11111111110000010000000100010011;
ROM[15942] <= 32'b00000000000000010010001110000011;
ROM[15943] <= 32'b00000000011100100010000000100011;
ROM[15944] <= 32'b00000000010000100000000100010011;
ROM[15945] <= 32'b00000001010000000000001110010011;
ROM[15946] <= 32'b01000000011100011000001110110011;
ROM[15947] <= 32'b00000000010000111010000110000011;
ROM[15948] <= 32'b00000000100000111010001000000011;
ROM[15949] <= 32'b00000000110000111010001010000011;
ROM[15950] <= 32'b00000001000000111010001100000011;
ROM[15951] <= 32'b00000000000000001000000011100111;
ROM[15952] <= 32'b00000000000000010010000000100011;
ROM[15953] <= 32'b00000000010000010000000100010011;
ROM[15954] <= 32'b00000000000000010010000000100011;
ROM[15955] <= 32'b00000000010000010000000100010011;
ROM[15956] <= 32'b00000000000000010010000000100011;
ROM[15957] <= 32'b00000000010000010000000100010011;
ROM[15958] <= 32'b00000000000000010010000000100011;
ROM[15959] <= 32'b00000000010000010000000100010011;
ROM[15960] <= 32'b00000000000000010010000000100011;
ROM[15961] <= 32'b00000000010000010000000100010011;
ROM[15962] <= 32'b00000000000000010010000000100011;
ROM[15963] <= 32'b00000000010000010000000100010011;
ROM[15964] <= 32'b00000000000000010010000000100011;
ROM[15965] <= 32'b00000000010000010000000100010011;
ROM[15966] <= 32'b00000000000000010010000000100011;
ROM[15967] <= 32'b00000000010000010000000100010011;
ROM[15968] <= 32'b00000000000000010010000000100011;
ROM[15969] <= 32'b00000000010000010000000100010011;
ROM[15970] <= 32'b00000000000000010010000000100011;
ROM[15971] <= 32'b00000000010000010000000100010011;
ROM[15972] <= 32'b00000000000000010010000000100011;
ROM[15973] <= 32'b00000000010000010000000100010011;
ROM[15974] <= 32'b00000000000000100010001110000011;
ROM[15975] <= 32'b00000000011100010010000000100011;
ROM[15976] <= 32'b00000000010000010000000100010011;
ROM[15977] <= 32'b00000000000000010000001110110111;
ROM[15978] <= 32'b10011111000000111000001110010011;
ROM[15979] <= 32'b00000000111000111000001110110011;
ROM[15980] <= 32'b00000000011100010010000000100011;
ROM[15981] <= 32'b00000000010000010000000100010011;
ROM[15982] <= 32'b00000000001100010010000000100011;
ROM[15983] <= 32'b00000000010000010000000100010011;
ROM[15984] <= 32'b00000000010000010010000000100011;
ROM[15985] <= 32'b00000000010000010000000100010011;
ROM[15986] <= 32'b00000000010100010010000000100011;
ROM[15987] <= 32'b00000000010000010000000100010011;
ROM[15988] <= 32'b00000000011000010010000000100011;
ROM[15989] <= 32'b00000000010000010000000100010011;
ROM[15990] <= 32'b00000001010000000000001110010011;
ROM[15991] <= 32'b00000000010000111000001110010011;
ROM[15992] <= 32'b01000000011100010000001110110011;
ROM[15993] <= 32'b00000000011100000000001000110011;
ROM[15994] <= 32'b00000000001000000000000110110011;
ROM[15995] <= 32'b11011101000111111111000011101111;
ROM[15996] <= 32'b11111111110000010000000100010011;
ROM[15997] <= 32'b00000000000000010010001110000011;
ROM[15998] <= 32'b00000000011100011010000000100011;
ROM[15999] <= 32'b00001000010001101010001110000011;
ROM[16000] <= 32'b00000000011100010010000000100011;
ROM[16001] <= 32'b00000000010000010000000100010011;
ROM[16002] <= 32'b00000000101000000000001110010011;
ROM[16003] <= 32'b00000000011100010010000000100011;
ROM[16004] <= 32'b00000000010000010000000100010011;
ROM[16005] <= 32'b00000000000000010000001110110111;
ROM[16006] <= 32'b10100110000000111000001110010011;
ROM[16007] <= 32'b00000000111000111000001110110011;
ROM[16008] <= 32'b00000000011100010010000000100011;
ROM[16009] <= 32'b00000000010000010000000100010011;
ROM[16010] <= 32'b00000000001100010010000000100011;
ROM[16011] <= 32'b00000000010000010000000100010011;
ROM[16012] <= 32'b00000000010000010010000000100011;
ROM[16013] <= 32'b00000000010000010000000100010011;
ROM[16014] <= 32'b00000000010100010010000000100011;
ROM[16015] <= 32'b00000000010000010000000100010011;
ROM[16016] <= 32'b00000000011000010010000000100011;
ROM[16017] <= 32'b00000000010000010000000100010011;
ROM[16018] <= 32'b00000001010000000000001110010011;
ROM[16019] <= 32'b00000000100000111000001110010011;
ROM[16020] <= 32'b01000000011100010000001110110011;
ROM[16021] <= 32'b00000000011100000000001000110011;
ROM[16022] <= 32'b00000000001000000000000110110011;
ROM[16023] <= 32'b11100111100011111001000011101111;
ROM[16024] <= 32'b00000000100000000000001110010011;
ROM[16025] <= 32'b00000000011100010010000000100011;
ROM[16026] <= 32'b00000000010000010000000100010011;
ROM[16027] <= 32'b00000000000000010000001110110111;
ROM[16028] <= 32'b10101011100000111000001110010011;
ROM[16029] <= 32'b00000000111000111000001110110011;
ROM[16030] <= 32'b00000000011100010010000000100011;
ROM[16031] <= 32'b00000000010000010000000100010011;
ROM[16032] <= 32'b00000000001100010010000000100011;
ROM[16033] <= 32'b00000000010000010000000100010011;
ROM[16034] <= 32'b00000000010000010010000000100011;
ROM[16035] <= 32'b00000000010000010000000100010011;
ROM[16036] <= 32'b00000000010100010010000000100011;
ROM[16037] <= 32'b00000000010000010000000100010011;
ROM[16038] <= 32'b00000000011000010010000000100011;
ROM[16039] <= 32'b00000000010000010000000100010011;
ROM[16040] <= 32'b00000001010000000000001110010011;
ROM[16041] <= 32'b00000000100000111000001110010011;
ROM[16042] <= 32'b01000000011100010000001110110011;
ROM[16043] <= 32'b00000000011100000000001000110011;
ROM[16044] <= 32'b00000000001000000000000110110011;
ROM[16045] <= 32'b11100010000011111001000011101111;
ROM[16046] <= 32'b00001000000001101010001110000011;
ROM[16047] <= 32'b00000000011100010010000000100011;
ROM[16048] <= 32'b00000000010000010000000100010011;
ROM[16049] <= 32'b00000000010000000000001110010011;
ROM[16050] <= 32'b00000000011100010010000000100011;
ROM[16051] <= 32'b00000000010000010000000100010011;
ROM[16052] <= 32'b00000000000000010000001110110111;
ROM[16053] <= 32'b10110001110000111000001110010011;
ROM[16054] <= 32'b00000000111000111000001110110011;
ROM[16055] <= 32'b00000000011100010010000000100011;
ROM[16056] <= 32'b00000000010000010000000100010011;
ROM[16057] <= 32'b00000000001100010010000000100011;
ROM[16058] <= 32'b00000000010000010000000100010011;
ROM[16059] <= 32'b00000000010000010010000000100011;
ROM[16060] <= 32'b00000000010000010000000100010011;
ROM[16061] <= 32'b00000000010100010010000000100011;
ROM[16062] <= 32'b00000000010000010000000100010011;
ROM[16063] <= 32'b00000000011000010010000000100011;
ROM[16064] <= 32'b00000000010000010000000100010011;
ROM[16065] <= 32'b00000001010000000000001110010011;
ROM[16066] <= 32'b00000000100000111000001110010011;
ROM[16067] <= 32'b01000000011100010000001110110011;
ROM[16068] <= 32'b00000000011100000000001000110011;
ROM[16069] <= 32'b00000000001000000000000110110011;
ROM[16070] <= 32'b11111110000011111001000011101111;
ROM[16071] <= 32'b11111111110000010000000100010011;
ROM[16072] <= 32'b00000000000000010010001110000011;
ROM[16073] <= 32'b11111111110000010000000100010011;
ROM[16074] <= 32'b00000000000000010010010000000011;
ROM[16075] <= 32'b00000000011101000000001110110011;
ROM[16076] <= 32'b00000000011100011010001000100011;
ROM[16077] <= 32'b00001000000001101010001110000011;
ROM[16078] <= 32'b00000000011100010010000000100011;
ROM[16079] <= 32'b00000000010000010000000100010011;
ROM[16080] <= 32'b00000000001100000000001110010011;
ROM[16081] <= 32'b11111111110000010000000100010011;
ROM[16082] <= 32'b00000000000000010010010000000011;
ROM[16083] <= 32'b00000000011101000111001110110011;
ROM[16084] <= 32'b00000000011100011010010000100011;
ROM[16085] <= 32'b00000000000000000000001110010011;
ROM[16086] <= 32'b00000000011100011010100000100011;
ROM[16087] <= 32'b00000001000000011010001110000011;
ROM[16088] <= 32'b00000000011100010010000000100011;
ROM[16089] <= 32'b00000000010000010000000100010011;
ROM[16090] <= 32'b00000000100000000000001110010011;
ROM[16091] <= 32'b11111111110000010000000100010011;
ROM[16092] <= 32'b00000000000000010010010000000011;
ROM[16093] <= 32'b00000000011101000010001110110011;
ROM[16094] <= 32'b01000000011100000000001110110011;
ROM[16095] <= 32'b00000000000100111000001110010011;
ROM[16096] <= 32'b00000000000000111000101001100011;
ROM[16097] <= 32'b00000000000000010000001110110111;
ROM[16098] <= 32'b01010100100000111000001110010011;
ROM[16099] <= 32'b00000000111000111000001110110011;
ROM[16100] <= 32'b00000000000000111000000011100111;
ROM[16101] <= 32'b00000001000000011010001110000011;
ROM[16102] <= 32'b00000000011100010010000000100011;
ROM[16103] <= 32'b00000000010000010000000100010011;
ROM[16104] <= 32'b00000000010000000000001110010011;
ROM[16105] <= 32'b00000000011100010010000000100011;
ROM[16106] <= 32'b00000000010000010000000100010011;
ROM[16107] <= 32'b00000000000000010000001110110111;
ROM[16108] <= 32'b10111111100000111000001110010011;
ROM[16109] <= 32'b00000000111000111000001110110011;
ROM[16110] <= 32'b00000000011100010010000000100011;
ROM[16111] <= 32'b00000000010000010000000100010011;
ROM[16112] <= 32'b00000000001100010010000000100011;
ROM[16113] <= 32'b00000000010000010000000100010011;
ROM[16114] <= 32'b00000000010000010010000000100011;
ROM[16115] <= 32'b00000000010000010000000100010011;
ROM[16116] <= 32'b00000000010100010010000000100011;
ROM[16117] <= 32'b00000000010000010000000100010011;
ROM[16118] <= 32'b00000000011000010010000000100011;
ROM[16119] <= 32'b00000000010000010000000100010011;
ROM[16120] <= 32'b00000001010000000000001110010011;
ROM[16121] <= 32'b00000000100000111000001110010011;
ROM[16122] <= 32'b01000000011100010000001110110011;
ROM[16123] <= 32'b00000000011100000000001000110011;
ROM[16124] <= 32'b00000000001000000000000110110011;
ROM[16125] <= 32'b11001110000011111001000011101111;
ROM[16126] <= 32'b11111111110000010000000100010011;
ROM[16127] <= 32'b00000000000000010010001110000011;
ROM[16128] <= 32'b00000000011100011010101000100011;
ROM[16129] <= 32'b00000001010000011010001110000011;
ROM[16130] <= 32'b00000000011100010010000000100011;
ROM[16131] <= 32'b00000000010000010000000100010011;
ROM[16132] <= 32'b00000000000000011010001110000011;
ROM[16133] <= 32'b11111111110000010000000100010011;
ROM[16134] <= 32'b00000000000000010010010000000011;
ROM[16135] <= 32'b00000000011101000000001110110011;
ROM[16136] <= 32'b00000000000000111000001100010011;
ROM[16137] <= 32'b00000000110100110000010000110011;
ROM[16138] <= 32'b00000000000001000010001110000011;
ROM[16139] <= 32'b00000000011100011010011000100011;
ROM[16140] <= 32'b00000000010000011010001110000011;
ROM[16141] <= 32'b00000000011100010010000000100011;
ROM[16142] <= 32'b00000000010000010000000100010011;
ROM[16143] <= 32'b00000000010000000000001110010011;
ROM[16144] <= 32'b00000000011100010010000000100011;
ROM[16145] <= 32'b00000000010000010000000100010011;
ROM[16146] <= 32'b00000000000000010000001110110111;
ROM[16147] <= 32'b11001001010000111000001110010011;
ROM[16148] <= 32'b00000000111000111000001110110011;
ROM[16149] <= 32'b00000000011100010010000000100011;
ROM[16150] <= 32'b00000000010000010000000100010011;
ROM[16151] <= 32'b00000000001100010010000000100011;
ROM[16152] <= 32'b00000000010000010000000100010011;
ROM[16153] <= 32'b00000000010000010010000000100011;
ROM[16154] <= 32'b00000000010000010000000100010011;
ROM[16155] <= 32'b00000000010100010010000000100011;
ROM[16156] <= 32'b00000000010000010000000100010011;
ROM[16157] <= 32'b00000000011000010010000000100011;
ROM[16158] <= 32'b00000000010000010000000100010011;
ROM[16159] <= 32'b00000001010000000000001110010011;
ROM[16160] <= 32'b00000000100000111000001110010011;
ROM[16161] <= 32'b01000000011100010000001110110011;
ROM[16162] <= 32'b00000000011100000000001000110011;
ROM[16163] <= 32'b00000000001000000000000110110011;
ROM[16164] <= 32'b11000100010011111001000011101111;
ROM[16165] <= 32'b11111111110000010000000100010011;
ROM[16166] <= 32'b00000000000000010010001110000011;
ROM[16167] <= 32'b00000000011100011010110000100011;
ROM[16168] <= 32'b00000000100000011010001110000011;
ROM[16169] <= 32'b00000000011100010010000000100011;
ROM[16170] <= 32'b00000000010000010000000100010011;
ROM[16171] <= 32'b00000000000000000000001110010011;
ROM[16172] <= 32'b11111111110000010000000100010011;
ROM[16173] <= 32'b00000000000000010010010000000011;
ROM[16174] <= 32'b00000000011101000010010010110011;
ROM[16175] <= 32'b00000000100000111010010100110011;
ROM[16176] <= 32'b00000000101001001000001110110011;
ROM[16177] <= 32'b00000000000100111000001110010011;
ROM[16178] <= 32'b00000000000100111111001110010011;
ROM[16179] <= 32'b00000000000000111000101001100011;
ROM[16180] <= 32'b00000000000000010000001110110111;
ROM[16181] <= 32'b11001110010000111000001110010011;
ROM[16182] <= 32'b00000000111000111000001110110011;
ROM[16183] <= 32'b00000000000000111000000011100111;
ROM[16184] <= 32'b00011110100000000000000011101111;
ROM[16185] <= 32'b00000001100000000000001110010011;
ROM[16186] <= 32'b00000000011100010010000000100011;
ROM[16187] <= 32'b00000000010000010000000100010011;
ROM[16188] <= 32'b00000000000000010000001110110111;
ROM[16189] <= 32'b11010011110000111000001110010011;
ROM[16190] <= 32'b00000000111000111000001110110011;
ROM[16191] <= 32'b00000000011100010010000000100011;
ROM[16192] <= 32'b00000000010000010000000100010011;
ROM[16193] <= 32'b00000000001100010010000000100011;
ROM[16194] <= 32'b00000000010000010000000100010011;
ROM[16195] <= 32'b00000000010000010010000000100011;
ROM[16196] <= 32'b00000000010000010000000100010011;
ROM[16197] <= 32'b00000000010100010010000000100011;
ROM[16198] <= 32'b00000000010000010000000100010011;
ROM[16199] <= 32'b00000000011000010010000000100011;
ROM[16200] <= 32'b00000000010000010000000100010011;
ROM[16201] <= 32'b00000001010000000000001110010011;
ROM[16202] <= 32'b00000000010000111000001110010011;
ROM[16203] <= 32'b01000000011100010000001110110011;
ROM[16204] <= 32'b00000000011100000000001000110011;
ROM[16205] <= 32'b00000000001000000000000110110011;
ROM[16206] <= 32'b10001100010111111001000011101111;
ROM[16207] <= 32'b11111111110000010000000100010011;
ROM[16208] <= 32'b00000000000000010010001110000011;
ROM[16209] <= 32'b00000010011100011010001000100011;
ROM[16210] <= 32'b00000000110000011010001110000011;
ROM[16211] <= 32'b00000000011100010010000000100011;
ROM[16212] <= 32'b00000000010000010000000100010011;
ROM[16213] <= 32'b00000001100000000000001110010011;
ROM[16214] <= 32'b00000000011100010010000000100011;
ROM[16215] <= 32'b00000000010000010000000100010011;
ROM[16216] <= 32'b00000000000000010000001110110111;
ROM[16217] <= 32'b11011010110000111000001110010011;
ROM[16218] <= 32'b00000000111000111000001110110011;
ROM[16219] <= 32'b00000000011100010010000000100011;
ROM[16220] <= 32'b00000000010000010000000100010011;
ROM[16221] <= 32'b00000000001100010010000000100011;
ROM[16222] <= 32'b00000000010000010000000100010011;
ROM[16223] <= 32'b00000000010000010010000000100011;
ROM[16224] <= 32'b00000000010000010000000100010011;
ROM[16225] <= 32'b00000000010100010010000000100011;
ROM[16226] <= 32'b00000000010000010000000100010011;
ROM[16227] <= 32'b00000000011000010010000000100011;
ROM[16228] <= 32'b00000000010000010000000100010011;
ROM[16229] <= 32'b00000001010000000000001110010011;
ROM[16230] <= 32'b00000000010000111000001110010011;
ROM[16231] <= 32'b01000000011100010000001110110011;
ROM[16232] <= 32'b00000000011100000000001000110011;
ROM[16233] <= 32'b00000000001000000000000110110011;
ROM[16234] <= 32'b10000101010111111001000011101111;
ROM[16235] <= 32'b00000000000000010000001110110111;
ROM[16236] <= 32'b11011111100000111000001110010011;
ROM[16237] <= 32'b00000000111000111000001110110011;
ROM[16238] <= 32'b00000000011100010010000000100011;
ROM[16239] <= 32'b00000000010000010000000100010011;
ROM[16240] <= 32'b00000000001100010010000000100011;
ROM[16241] <= 32'b00000000010000010000000100010011;
ROM[16242] <= 32'b00000000010000010010000000100011;
ROM[16243] <= 32'b00000000010000010000000100010011;
ROM[16244] <= 32'b00000000010100010010000000100011;
ROM[16245] <= 32'b00000000010000010000000100010011;
ROM[16246] <= 32'b00000000011000010010000000100011;
ROM[16247] <= 32'b00000000010000010000000100010011;
ROM[16248] <= 32'b00000001010000000000001110010011;
ROM[16249] <= 32'b00000000100000111000001110010011;
ROM[16250] <= 32'b01000000011100010000001110110011;
ROM[16251] <= 32'b00000000011100000000001000110011;
ROM[16252] <= 32'b00000000001000000000000110110011;
ROM[16253] <= 32'b10101110000011111001000011101111;
ROM[16254] <= 32'b11111111110000010000000100010011;
ROM[16255] <= 32'b00000000000000010010001110000011;
ROM[16256] <= 32'b00000000011100011010011000100011;
ROM[16257] <= 32'b00000010010000011010001110000011;
ROM[16258] <= 32'b00000000011100010010000000100011;
ROM[16259] <= 32'b00000000010000010000000100010011;
ROM[16260] <= 32'b00000000000100000000001110010011;
ROM[16261] <= 32'b11111111110000010000000100010011;
ROM[16262] <= 32'b00000000000000010010010000000011;
ROM[16263] <= 32'b01000000011101000000001110110011;
ROM[16264] <= 32'b00000010011100011010001000100011;
ROM[16265] <= 32'b00000001100000011010001110000011;
ROM[16266] <= 32'b00000000011100010010000000100011;
ROM[16267] <= 32'b00000000010000010000000100010011;
ROM[16268] <= 32'b00000111110001101010001110000011;
ROM[16269] <= 32'b11111111110000010000000100010011;
ROM[16270] <= 32'b00000000000000010010010000000011;
ROM[16271] <= 32'b00000000011101000000001110110011;
ROM[16272] <= 32'b00000000000000111000001100010011;
ROM[16273] <= 32'b00000000110100110000010000110011;
ROM[16274] <= 32'b00000000000001000010001110000011;
ROM[16275] <= 32'b00000000011100010010000000100011;
ROM[16276] <= 32'b00000000010000010000000100010011;
ROM[16277] <= 32'b00000010010000011010001110000011;
ROM[16278] <= 32'b11111111110000010000000100010011;
ROM[16279] <= 32'b00000000000000010010010000000011;
ROM[16280] <= 32'b00000000011101000111001110110011;
ROM[16281] <= 32'b00000000011100010010000000100011;
ROM[16282] <= 32'b00000000010000010000000100010011;
ROM[16283] <= 32'b00000000110000011010001110000011;
ROM[16284] <= 32'b11111111110000010000000100010011;
ROM[16285] <= 32'b00000000000000010010010000000011;
ROM[16286] <= 32'b00000000011101000110001110110011;
ROM[16287] <= 32'b00000010011100011010010000100011;
ROM[16288] <= 32'b00000001100000011010001110000011;
ROM[16289] <= 32'b00000000011100010010000000100011;
ROM[16290] <= 32'b00000000010000010000000100010011;
ROM[16291] <= 32'b00000111110001101010001110000011;
ROM[16292] <= 32'b11111111110000010000000100010011;
ROM[16293] <= 32'b00000000000000010010010000000011;
ROM[16294] <= 32'b00000000011101000000001110110011;
ROM[16295] <= 32'b00000000011100010010000000100011;
ROM[16296] <= 32'b00000000010000010000000100010011;
ROM[16297] <= 32'b00000010100000011010001110000011;
ROM[16298] <= 32'b00000000011101100010000000100011;
ROM[16299] <= 32'b11111111110000010000000100010011;
ROM[16300] <= 32'b00000000000000010010001110000011;
ROM[16301] <= 32'b00000000000000111000001100010011;
ROM[16302] <= 32'b00000000000001100010001110000011;
ROM[16303] <= 32'b00000000110100110000010000110011;
ROM[16304] <= 32'b00000000011101000010000000100011;
ROM[16305] <= 32'b01100100000000000000000011101111;
ROM[16306] <= 32'b00000000100000011010001110000011;
ROM[16307] <= 32'b00000000011100010010000000100011;
ROM[16308] <= 32'b00000000010000010000000100010011;
ROM[16309] <= 32'b00000000000100000000001110010011;
ROM[16310] <= 32'b11111111110000010000000100010011;
ROM[16311] <= 32'b00000000000000010010010000000011;
ROM[16312] <= 32'b00000000011101000010010010110011;
ROM[16313] <= 32'b00000000100000111010010100110011;
ROM[16314] <= 32'b00000000101001001000001110110011;
ROM[16315] <= 32'b00000000000100111000001110010011;
ROM[16316] <= 32'b00000000000100111111001110010011;
ROM[16317] <= 32'b00000000000000111000101001100011;
ROM[16318] <= 32'b00000000000000010000001110110111;
ROM[16319] <= 32'b11110000110000111000001110010011;
ROM[16320] <= 32'b00000000111000111000001110110011;
ROM[16321] <= 32'b00000000000000111000000011100111;
ROM[16322] <= 32'b00101000110000000000000011101111;
ROM[16323] <= 32'b00000001100000000000001110010011;
ROM[16324] <= 32'b00000000011100010010000000100011;
ROM[16325] <= 32'b00000000010000010000000100010011;
ROM[16326] <= 32'b00000000000000010000001110110111;
ROM[16327] <= 32'b11110110010000111000001110010011;
ROM[16328] <= 32'b00000000111000111000001110110011;
ROM[16329] <= 32'b00000000011100010010000000100011;
ROM[16330] <= 32'b00000000010000010000000100010011;
ROM[16331] <= 32'b00000000001100010010000000100011;
ROM[16332] <= 32'b00000000010000010000000100010011;
ROM[16333] <= 32'b00000000010000010010000000100011;
ROM[16334] <= 32'b00000000010000010000000100010011;
ROM[16335] <= 32'b00000000010100010010000000100011;
ROM[16336] <= 32'b00000000010000010000000100010011;
ROM[16337] <= 32'b00000000011000010010000000100011;
ROM[16338] <= 32'b00000000010000010000000100010011;
ROM[16339] <= 32'b00000001010000000000001110010011;
ROM[16340] <= 32'b00000000010000111000001110010011;
ROM[16341] <= 32'b01000000011100010000001110110011;
ROM[16342] <= 32'b00000000011100000000001000110011;
ROM[16343] <= 32'b00000000001000000000000110110011;
ROM[16344] <= 32'b11101001110011111001000011101111;
ROM[16345] <= 32'b00000001000000000000001110010011;
ROM[16346] <= 32'b00000000011100010010000000100011;
ROM[16347] <= 32'b00000000010000010000000100010011;
ROM[16348] <= 32'b00000000000000010000001110110111;
ROM[16349] <= 32'b11111011110000111000001110010011;
ROM[16350] <= 32'b00000000111000111000001110110011;
ROM[16351] <= 32'b00000000011100010010000000100011;
ROM[16352] <= 32'b00000000010000010000000100010011;
ROM[16353] <= 32'b00000000001100010010000000100011;
ROM[16354] <= 32'b00000000010000010000000100010011;
ROM[16355] <= 32'b00000000010000010010000000100011;
ROM[16356] <= 32'b00000000010000010000000100010011;
ROM[16357] <= 32'b00000000010100010010000000100011;
ROM[16358] <= 32'b00000000010000010000000100010011;
ROM[16359] <= 32'b00000000011000010010000000100011;
ROM[16360] <= 32'b00000000010000010000000100010011;
ROM[16361] <= 32'b00000001010000000000001110010011;
ROM[16362] <= 32'b00000000010000111000001110010011;
ROM[16363] <= 32'b01000000011100010000001110110011;
ROM[16364] <= 32'b00000000011100000000001000110011;
ROM[16365] <= 32'b00000000001000000000000110110011;
ROM[16366] <= 32'b11100100010011111001000011101111;
ROM[16367] <= 32'b11111111110000010000000100010011;
ROM[16368] <= 32'b00000000000000010010001110000011;
ROM[16369] <= 32'b11111111110000010000000100010011;
ROM[16370] <= 32'b00000000000000010010010000000011;
ROM[16371] <= 32'b01000000011101000000001110110011;
ROM[16372] <= 32'b00000000011100011010111000100011;
ROM[16373] <= 32'b00000000000000000000001110010011;
ROM[16374] <= 32'b00000000011100010010000000100011;
ROM[16375] <= 32'b00000000010000010000000100010011;
ROM[16376] <= 32'b00000001110000011010001110000011;
ROM[16377] <= 32'b11111111110000010000000100010011;
ROM[16378] <= 32'b00000000000000010010010000000011;
ROM[16379] <= 32'b01000000011101000000001110110011;
ROM[16380] <= 32'b00000010011100011010001000100011;
ROM[16381] <= 32'b00000010010000011010001110000011;
ROM[16382] <= 32'b00000000011100010010000000100011;
ROM[16383] <= 32'b00000000010000010000000100010011;
ROM[16384] <= 32'b00000000000100000000001110010011;
ROM[16385] <= 32'b11111111110000010000000100010011;
ROM[16386] <= 32'b00000000000000010010010000000011;
ROM[16387] <= 32'b01000000011101000000001110110011;
ROM[16388] <= 32'b00000010011100011010001000100011;
ROM[16389] <= 32'b00000000110000011010001110000011;
ROM[16390] <= 32'b00000000011100010010000000100011;
ROM[16391] <= 32'b00000000010000010000000100010011;
ROM[16392] <= 32'b00000001000000000000001110010011;
ROM[16393] <= 32'b00000000011100010010000000100011;
ROM[16394] <= 32'b00000000010000010000000100010011;
ROM[16395] <= 32'b00000000000000010000001110110111;
ROM[16396] <= 32'b00000111100000111000001110010011;
ROM[16397] <= 32'b00000000111000111000001110110011;
ROM[16398] <= 32'b00000000011100010010000000100011;
ROM[16399] <= 32'b00000000010000010000000100010011;
ROM[16400] <= 32'b00000000001100010010000000100011;
ROM[16401] <= 32'b00000000010000010000000100010011;
ROM[16402] <= 32'b00000000010000010010000000100011;
ROM[16403] <= 32'b00000000010000010000000100010011;
ROM[16404] <= 32'b00000000010100010010000000100011;
ROM[16405] <= 32'b00000000010000010000000100010011;
ROM[16406] <= 32'b00000000011000010010000000100011;
ROM[16407] <= 32'b00000000010000010000000100010011;
ROM[16408] <= 32'b00000001010000000000001110010011;
ROM[16409] <= 32'b00000000010000111000001110010011;
ROM[16410] <= 32'b01000000011100010000001110110011;
ROM[16411] <= 32'b00000000011100000000001000110011;
ROM[16412] <= 32'b00000000001000000000000110110011;
ROM[16413] <= 32'b11011000100011111001000011101111;
ROM[16414] <= 32'b00000000000000010000001110110111;
ROM[16415] <= 32'b00001100010000111000001110010011;
ROM[16416] <= 32'b00000000111000111000001110110011;
ROM[16417] <= 32'b00000000011100010010000000100011;
ROM[16418] <= 32'b00000000010000010000000100010011;
ROM[16419] <= 32'b00000000001100010010000000100011;
ROM[16420] <= 32'b00000000010000010000000100010011;
ROM[16421] <= 32'b00000000010000010010000000100011;
ROM[16422] <= 32'b00000000010000010000000100010011;
ROM[16423] <= 32'b00000000010100010010000000100011;
ROM[16424] <= 32'b00000000010000010000000100010011;
ROM[16425] <= 32'b00000000011000010010000000100011;
ROM[16426] <= 32'b00000000010000010000000100010011;
ROM[16427] <= 32'b00000001010000000000001110010011;
ROM[16428] <= 32'b00000000100000111000001110010011;
ROM[16429] <= 32'b01000000011100010000001110110011;
ROM[16430] <= 32'b00000000011100000000001000110011;
ROM[16431] <= 32'b00000000001000000000000110110011;
ROM[16432] <= 32'b10000001010011111001000011101111;
ROM[16433] <= 32'b11111111110000010000000100010011;
ROM[16434] <= 32'b00000000000000010010001110000011;
ROM[16435] <= 32'b00000000011100011010011000100011;
ROM[16436] <= 32'b00000000110000011010001110000011;
ROM[16437] <= 32'b00000000011100010010000000100011;
ROM[16438] <= 32'b00000000010000010000000100010011;
ROM[16439] <= 32'b00000001110000011010001110000011;
ROM[16440] <= 32'b11111111110000010000000100010011;
ROM[16441] <= 32'b00000000000000010010010000000011;
ROM[16442] <= 32'b00000000011101000111001110110011;
ROM[16443] <= 32'b00000000011100011010011000100011;
ROM[16444] <= 32'b00000001100000011010001110000011;
ROM[16445] <= 32'b00000000011100010010000000100011;
ROM[16446] <= 32'b00000000010000010000000100010011;
ROM[16447] <= 32'b00000111110001101010001110000011;
ROM[16448] <= 32'b11111111110000010000000100010011;
ROM[16449] <= 32'b00000000000000010010010000000011;
ROM[16450] <= 32'b00000000011101000000001110110011;
ROM[16451] <= 32'b00000000000000111000001100010011;
ROM[16452] <= 32'b00000000110100110000010000110011;
ROM[16453] <= 32'b00000000000001000010001110000011;
ROM[16454] <= 32'b00000000011100010010000000100011;
ROM[16455] <= 32'b00000000010000010000000100010011;
ROM[16456] <= 32'b00000010010000011010001110000011;
ROM[16457] <= 32'b11111111110000010000000100010011;
ROM[16458] <= 32'b00000000000000010010010000000011;
ROM[16459] <= 32'b00000000011101000111001110110011;
ROM[16460] <= 32'b00000000011100010010000000100011;
ROM[16461] <= 32'b00000000010000010000000100010011;
ROM[16462] <= 32'b00000000110000011010001110000011;
ROM[16463] <= 32'b11111111110000010000000100010011;
ROM[16464] <= 32'b00000000000000010010010000000011;
ROM[16465] <= 32'b00000000011101000110001110110011;
ROM[16466] <= 32'b00000010011100011010010000100011;
ROM[16467] <= 32'b00000001100000011010001110000011;
ROM[16468] <= 32'b00000000011100010010000000100011;
ROM[16469] <= 32'b00000000010000010000000100010011;
ROM[16470] <= 32'b00000111110001101010001110000011;
ROM[16471] <= 32'b11111111110000010000000100010011;
ROM[16472] <= 32'b00000000000000010010010000000011;
ROM[16473] <= 32'b00000000011101000000001110110011;
ROM[16474] <= 32'b00000000011100010010000000100011;
ROM[16475] <= 32'b00000000010000010000000100010011;
ROM[16476] <= 32'b00000010100000011010001110000011;
ROM[16477] <= 32'b00000000011101100010000000100011;
ROM[16478] <= 32'b11111111110000010000000100010011;
ROM[16479] <= 32'b00000000000000010010001110000011;
ROM[16480] <= 32'b00000000000000111000001100010011;
ROM[16481] <= 32'b00000000000001100010001110000011;
ROM[16482] <= 32'b00000000110100110000010000110011;
ROM[16483] <= 32'b00000000011101000010000000100011;
ROM[16484] <= 32'b00110111010000000000000011101111;
ROM[16485] <= 32'b00000000100000011010001110000011;
ROM[16486] <= 32'b00000000011100010010000000100011;
ROM[16487] <= 32'b00000000010000010000000100010011;
ROM[16488] <= 32'b00000000001000000000001110010011;
ROM[16489] <= 32'b11111111110000010000000100010011;
ROM[16490] <= 32'b00000000000000010010010000000011;
ROM[16491] <= 32'b00000000011101000010010010110011;
ROM[16492] <= 32'b00000000100000111010010100110011;
ROM[16493] <= 32'b00000000101001001000001110110011;
ROM[16494] <= 32'b00000000000100111000001110010011;
ROM[16495] <= 32'b00000000000100111111001110010011;
ROM[16496] <= 32'b00000000000000111000101001100011;
ROM[16497] <= 32'b00000000000000010000001110110111;
ROM[16498] <= 32'b00011101100000111000001110010011;
ROM[16499] <= 32'b00000000111000111000001110110011;
ROM[16500] <= 32'b00000000000000111000000011100111;
ROM[16501] <= 32'b00101000110000000000000011101111;
ROM[16502] <= 32'b00000001000000000000001110010011;
ROM[16503] <= 32'b00000000011100010010000000100011;
ROM[16504] <= 32'b00000000010000010000000100010011;
ROM[16505] <= 32'b00000000000000010000001110110111;
ROM[16506] <= 32'b00100011000000111000001110010011;
ROM[16507] <= 32'b00000000111000111000001110110011;
ROM[16508] <= 32'b00000000011100010010000000100011;
ROM[16509] <= 32'b00000000010000010000000100010011;
ROM[16510] <= 32'b00000000001100010010000000100011;
ROM[16511] <= 32'b00000000010000010000000100010011;
ROM[16512] <= 32'b00000000010000010010000000100011;
ROM[16513] <= 32'b00000000010000010000000100010011;
ROM[16514] <= 32'b00000000010100010010000000100011;
ROM[16515] <= 32'b00000000010000010000000100010011;
ROM[16516] <= 32'b00000000011000010010000000100011;
ROM[16517] <= 32'b00000000010000010000000100010011;
ROM[16518] <= 32'b00000001010000000000001110010011;
ROM[16519] <= 32'b00000000010000111000001110010011;
ROM[16520] <= 32'b01000000011100010000001110110011;
ROM[16521] <= 32'b00000000011100000000001000110011;
ROM[16522] <= 32'b00000000001000000000000110110011;
ROM[16523] <= 32'b10111101000011111001000011101111;
ROM[16524] <= 32'b00000000100000000000001110010011;
ROM[16525] <= 32'b00000000011100010010000000100011;
ROM[16526] <= 32'b00000000010000010000000100010011;
ROM[16527] <= 32'b00000000000000010000001110110111;
ROM[16528] <= 32'b00101000100000111000001110010011;
ROM[16529] <= 32'b00000000111000111000001110110011;
ROM[16530] <= 32'b00000000011100010010000000100011;
ROM[16531] <= 32'b00000000010000010000000100010011;
ROM[16532] <= 32'b00000000001100010010000000100011;
ROM[16533] <= 32'b00000000010000010000000100010011;
ROM[16534] <= 32'b00000000010000010010000000100011;
ROM[16535] <= 32'b00000000010000010000000100010011;
ROM[16536] <= 32'b00000000010100010010000000100011;
ROM[16537] <= 32'b00000000010000010000000100010011;
ROM[16538] <= 32'b00000000011000010010000000100011;
ROM[16539] <= 32'b00000000010000010000000100010011;
ROM[16540] <= 32'b00000001010000000000001110010011;
ROM[16541] <= 32'b00000000010000111000001110010011;
ROM[16542] <= 32'b01000000011100010000001110110011;
ROM[16543] <= 32'b00000000011100000000001000110011;
ROM[16544] <= 32'b00000000001000000000000110110011;
ROM[16545] <= 32'b10110111100011111001000011101111;
ROM[16546] <= 32'b11111111110000010000000100010011;
ROM[16547] <= 32'b00000000000000010010001110000011;
ROM[16548] <= 32'b11111111110000010000000100010011;
ROM[16549] <= 32'b00000000000000010010010000000011;
ROM[16550] <= 32'b01000000011101000000001110110011;
ROM[16551] <= 32'b00000010011100011010000000100011;
ROM[16552] <= 32'b00000000000000000000001110010011;
ROM[16553] <= 32'b00000000011100010010000000100011;
ROM[16554] <= 32'b00000000010000010000000100010011;
ROM[16555] <= 32'b00000010000000011010001110000011;
ROM[16556] <= 32'b11111111110000010000000100010011;
ROM[16557] <= 32'b00000000000000010010010000000011;
ROM[16558] <= 32'b01000000011101000000001110110011;
ROM[16559] <= 32'b00000010011100011010001000100011;
ROM[16560] <= 32'b00000010010000011010001110000011;
ROM[16561] <= 32'b00000000011100010010000000100011;
ROM[16562] <= 32'b00000000010000010000000100010011;
ROM[16563] <= 32'b00000000000100000000001110010011;
ROM[16564] <= 32'b11111111110000010000000100010011;
ROM[16565] <= 32'b00000000000000010010010000000011;
ROM[16566] <= 32'b01000000011101000000001110110011;
ROM[16567] <= 32'b00000010011100011010001000100011;
ROM[16568] <= 32'b00000000110000011010001110000011;
ROM[16569] <= 32'b00000000011100010010000000100011;
ROM[16570] <= 32'b00000000010000010000000100010011;
ROM[16571] <= 32'b00000000100000000000001110010011;
ROM[16572] <= 32'b00000000011100010010000000100011;
ROM[16573] <= 32'b00000000010000010000000100010011;
ROM[16574] <= 32'b00000000000000010000001110110111;
ROM[16575] <= 32'b00110100010000111000001110010011;
ROM[16576] <= 32'b00000000111000111000001110110011;
ROM[16577] <= 32'b00000000011100010010000000100011;
ROM[16578] <= 32'b00000000010000010000000100010011;
ROM[16579] <= 32'b00000000001100010010000000100011;
ROM[16580] <= 32'b00000000010000010000000100010011;
ROM[16581] <= 32'b00000000010000010010000000100011;
ROM[16582] <= 32'b00000000010000010000000100010011;
ROM[16583] <= 32'b00000000010100010010000000100011;
ROM[16584] <= 32'b00000000010000010000000100010011;
ROM[16585] <= 32'b00000000011000010010000000100011;
ROM[16586] <= 32'b00000000010000010000000100010011;
ROM[16587] <= 32'b00000001010000000000001110010011;
ROM[16588] <= 32'b00000000010000111000001110010011;
ROM[16589] <= 32'b01000000011100010000001110110011;
ROM[16590] <= 32'b00000000011100000000001000110011;
ROM[16591] <= 32'b00000000001000000000000110110011;
ROM[16592] <= 32'b10101011110011111001000011101111;
ROM[16593] <= 32'b00000000000000010000001110110111;
ROM[16594] <= 32'b00111001000000111000001110010011;
ROM[16595] <= 32'b00000000111000111000001110110011;
ROM[16596] <= 32'b00000000011100010010000000100011;
ROM[16597] <= 32'b00000000010000010000000100010011;
ROM[16598] <= 32'b00000000001100010010000000100011;
ROM[16599] <= 32'b00000000010000010000000100010011;
ROM[16600] <= 32'b00000000010000010010000000100011;
ROM[16601] <= 32'b00000000010000010000000100010011;
ROM[16602] <= 32'b00000000010100010010000000100011;
ROM[16603] <= 32'b00000000010000010000000100010011;
ROM[16604] <= 32'b00000000011000010010000000100011;
ROM[16605] <= 32'b00000000010000010000000100010011;
ROM[16606] <= 32'b00000001010000000000001110010011;
ROM[16607] <= 32'b00000000100000111000001110010011;
ROM[16608] <= 32'b01000000011100010000001110110011;
ROM[16609] <= 32'b00000000011100000000001000110011;
ROM[16610] <= 32'b00000000001000000000000110110011;
ROM[16611] <= 32'b11010100100111111000000011101111;
ROM[16612] <= 32'b11111111110000010000000100010011;
ROM[16613] <= 32'b00000000000000010010001110000011;
ROM[16614] <= 32'b00000000011100011010011000100011;
ROM[16615] <= 32'b00000000110000011010001110000011;
ROM[16616] <= 32'b00000000011100010010000000100011;
ROM[16617] <= 32'b00000000010000010000000100010011;
ROM[16618] <= 32'b00000010000000011010001110000011;
ROM[16619] <= 32'b11111111110000010000000100010011;
ROM[16620] <= 32'b00000000000000010010010000000011;
ROM[16621] <= 32'b00000000011101000111001110110011;
ROM[16622] <= 32'b00000000011100011010011000100011;
ROM[16623] <= 32'b00000001100000011010001110000011;
ROM[16624] <= 32'b00000000011100010010000000100011;
ROM[16625] <= 32'b00000000010000010000000100010011;
ROM[16626] <= 32'b00000111110001101010001110000011;
ROM[16627] <= 32'b11111111110000010000000100010011;
ROM[16628] <= 32'b00000000000000010010010000000011;
ROM[16629] <= 32'b00000000011101000000001110110011;
ROM[16630] <= 32'b00000000000000111000001100010011;
ROM[16631] <= 32'b00000000110100110000010000110011;
ROM[16632] <= 32'b00000000000001000010001110000011;
ROM[16633] <= 32'b00000000011100010010000000100011;
ROM[16634] <= 32'b00000000010000010000000100010011;
ROM[16635] <= 32'b00000010010000011010001110000011;
ROM[16636] <= 32'b11111111110000010000000100010011;
ROM[16637] <= 32'b00000000000000010010010000000011;
ROM[16638] <= 32'b00000000011101000111001110110011;
ROM[16639] <= 32'b00000000011100010010000000100011;
ROM[16640] <= 32'b00000000010000010000000100010011;
ROM[16641] <= 32'b00000000110000011010001110000011;
ROM[16642] <= 32'b11111111110000010000000100010011;
ROM[16643] <= 32'b00000000000000010010010000000011;
ROM[16644] <= 32'b00000000011101000110001110110011;
ROM[16645] <= 32'b00000010011100011010010000100011;
ROM[16646] <= 32'b00000001100000011010001110000011;
ROM[16647] <= 32'b00000000011100010010000000100011;
ROM[16648] <= 32'b00000000010000010000000100010011;
ROM[16649] <= 32'b00000111110001101010001110000011;
ROM[16650] <= 32'b11111111110000010000000100010011;
ROM[16651] <= 32'b00000000000000010010010000000011;
ROM[16652] <= 32'b00000000011101000000001110110011;
ROM[16653] <= 32'b00000000011100010010000000100011;
ROM[16654] <= 32'b00000000010000010000000100010011;
ROM[16655] <= 32'b00000010100000011010001110000011;
ROM[16656] <= 32'b00000000011101100010000000100011;
ROM[16657] <= 32'b11111111110000010000000100010011;
ROM[16658] <= 32'b00000000000000010010001110000011;
ROM[16659] <= 32'b00000000000000111000001100010011;
ROM[16660] <= 32'b00000000000001100010001110000011;
ROM[16661] <= 32'b00000000110100110000010000110011;
ROM[16662] <= 32'b00000000011101000010000000100011;
ROM[16663] <= 32'b00001010100000000000000011101111;
ROM[16664] <= 32'b00000001100000011010001110000011;
ROM[16665] <= 32'b00000000011100010010000000100011;
ROM[16666] <= 32'b00000000010000010000000100010011;
ROM[16667] <= 32'b00000111110001101010001110000011;
ROM[16668] <= 32'b11111111110000010000000100010011;
ROM[16669] <= 32'b00000000000000010010010000000011;
ROM[16670] <= 32'b00000000011101000000001110110011;
ROM[16671] <= 32'b00000000000000111000001100010011;
ROM[16672] <= 32'b00000000110100110000010000110011;
ROM[16673] <= 32'b00000000000001000010001110000011;
ROM[16674] <= 32'b00000000011100010010000000100011;
ROM[16675] <= 32'b00000000010000010000000100010011;
ROM[16676] <= 32'b00010000000000000000001110010011;
ROM[16677] <= 32'b01000000011100000000001110110011;
ROM[16678] <= 32'b11111111110000010000000100010011;
ROM[16679] <= 32'b00000000000000010010010000000011;
ROM[16680] <= 32'b00000000011101000111001110110011;
ROM[16681] <= 32'b00000000011100010010000000100011;
ROM[16682] <= 32'b00000000010000010000000100010011;
ROM[16683] <= 32'b00000000110000011010001110000011;
ROM[16684] <= 32'b11111111110000010000000100010011;
ROM[16685] <= 32'b00000000000000010010010000000011;
ROM[16686] <= 32'b00000000011101000110001110110011;
ROM[16687] <= 32'b00000010011100011010010000100011;
ROM[16688] <= 32'b00000001100000011010001110000011;
ROM[16689] <= 32'b00000000011100010010000000100011;
ROM[16690] <= 32'b00000000010000010000000100010011;
ROM[16691] <= 32'b00000111110001101010001110000011;
ROM[16692] <= 32'b11111111110000010000000100010011;
ROM[16693] <= 32'b00000000000000010010010000000011;
ROM[16694] <= 32'b00000000011101000000001110110011;
ROM[16695] <= 32'b00000000011100010010000000100011;
ROM[16696] <= 32'b00000000010000010000000100010011;
ROM[16697] <= 32'b00000010100000011010001110000011;
ROM[16698] <= 32'b00000000011101100010000000100011;
ROM[16699] <= 32'b11111111110000010000000100010011;
ROM[16700] <= 32'b00000000000000010010001110000011;
ROM[16701] <= 32'b00000000000000111000001100010011;
ROM[16702] <= 32'b00000000000001100010001110000011;
ROM[16703] <= 32'b00000000110100110000010000110011;
ROM[16704] <= 32'b00000000011101000010000000100011;
ROM[16705] <= 32'b00000000010000011010001110000011;
ROM[16706] <= 32'b00000000011100010010000000100011;
ROM[16707] <= 32'b00000000010000010000000100010011;
ROM[16708] <= 32'b00000000101000000000001110010011;
ROM[16709] <= 32'b11111111110000010000000100010011;
ROM[16710] <= 32'b00000000000000010010010000000011;
ROM[16711] <= 32'b00000000011101000000001110110011;
ROM[16712] <= 32'b00000000011100011010001000100011;
ROM[16713] <= 32'b00000001000000011010001110000011;
ROM[16714] <= 32'b00000000011100010010000000100011;
ROM[16715] <= 32'b00000000010000010000000100010011;
ROM[16716] <= 32'b00000000000100000000001110010011;
ROM[16717] <= 32'b11111111110000010000000100010011;
ROM[16718] <= 32'b00000000000000010010010000000011;
ROM[16719] <= 32'b00000000011101000000001110110011;
ROM[16720] <= 32'b00000000011100011010100000100011;
ROM[16721] <= 32'b11100001100011111111000011101111;
ROM[16722] <= 32'b00001000000001101010001110000011;
ROM[16723] <= 32'b00000000011100010010000000100011;
ROM[16724] <= 32'b00000000010000010000000100010011;
ROM[16725] <= 32'b00000010011100000000001110010011;
ROM[16726] <= 32'b11111111110000010000000100010011;
ROM[16727] <= 32'b00000000000000010010010000000011;
ROM[16728] <= 32'b00000000011101000010010010110011;
ROM[16729] <= 32'b00000000100000111010010100110011;
ROM[16730] <= 32'b00000000101001001000001110110011;
ROM[16731] <= 32'b00000000000100111000001110010011;
ROM[16732] <= 32'b00000000000100111111001110010011;
ROM[16733] <= 32'b00000000000000111000101001100011;
ROM[16734] <= 32'b00000000000000010000001110110111;
ROM[16735] <= 32'b01011000110000111000001110010011;
ROM[16736] <= 32'b00000000111000111000001110110011;
ROM[16737] <= 32'b00000000000000111000000011100111;
ROM[16738] <= 32'b00000110000000000000000011101111;
ROM[16739] <= 32'b00000000000000010000001110110111;
ROM[16740] <= 32'b01011101100000111000001110010011;
ROM[16741] <= 32'b00000000111000111000001110110011;
ROM[16742] <= 32'b00000000011100010010000000100011;
ROM[16743] <= 32'b00000000010000010000000100010011;
ROM[16744] <= 32'b00000000001100010010000000100011;
ROM[16745] <= 32'b00000000010000010000000100010011;
ROM[16746] <= 32'b00000000010000010010000000100011;
ROM[16747] <= 32'b00000000010000010000000100010011;
ROM[16748] <= 32'b00000000010100010010000000100011;
ROM[16749] <= 32'b00000000010000010000000100010011;
ROM[16750] <= 32'b00000000011000010010000000100011;
ROM[16751] <= 32'b00000000010000010000000100010011;
ROM[16752] <= 32'b00000001010000000000001110010011;
ROM[16753] <= 32'b00000000000000111000001110010011;
ROM[16754] <= 32'b01000000011100010000001110110011;
ROM[16755] <= 32'b00000000011100000000001000110011;
ROM[16756] <= 32'b00000000001000000000000110110011;
ROM[16757] <= 32'b01001001000000000000000011101111;
ROM[16758] <= 32'b11111111110000010000000100010011;
ROM[16759] <= 32'b00000000000000010010001110000011;
ROM[16760] <= 32'b00000000011101100010000000100011;
ROM[16761] <= 32'b00001000110000000000000011101111;
ROM[16762] <= 32'b00001000010001101010001110000011;
ROM[16763] <= 32'b00000000011100010010000000100011;
ROM[16764] <= 32'b00000000010000010000000100010011;
ROM[16765] <= 32'b00001000000001101010001110000011;
ROM[16766] <= 32'b00000000011100010010000000100011;
ROM[16767] <= 32'b00000000010000010000000100010011;
ROM[16768] <= 32'b00000000000100000000001110010011;
ROM[16769] <= 32'b11111111110000010000000100010011;
ROM[16770] <= 32'b00000000000000010010010000000011;
ROM[16771] <= 32'b00000000011101000000001110110011;
ROM[16772] <= 32'b00000000011100010010000000100011;
ROM[16773] <= 32'b00000000010000010000000100010011;
ROM[16774] <= 32'b00000000000000010000001110110111;
ROM[16775] <= 32'b01100110010000111000001110010011;
ROM[16776] <= 32'b00000000111000111000001110110011;
ROM[16777] <= 32'b00000000011100010010000000100011;
ROM[16778] <= 32'b00000000010000010000000100010011;
ROM[16779] <= 32'b00000000001100010010000000100011;
ROM[16780] <= 32'b00000000010000010000000100010011;
ROM[16781] <= 32'b00000000010000010010000000100011;
ROM[16782] <= 32'b00000000010000010000000100010011;
ROM[16783] <= 32'b00000000010100010010000000100011;
ROM[16784] <= 32'b00000000010000010000000100010011;
ROM[16785] <= 32'b00000000011000010010000000100011;
ROM[16786] <= 32'b00000000010000010000000100010011;
ROM[16787] <= 32'b00000001010000000000001110010011;
ROM[16788] <= 32'b00000000100000111000001110010011;
ROM[16789] <= 32'b01000000011100010000001110110011;
ROM[16790] <= 32'b00000000011100000000001000110011;
ROM[16791] <= 32'b00000000001000000000000110110011;
ROM[16792] <= 32'b10101000110011111111000011101111;
ROM[16793] <= 32'b11111111110000010000000100010011;
ROM[16794] <= 32'b00000000000000010010001110000011;
ROM[16795] <= 32'b00000000011101100010000000100011;
ROM[16796] <= 32'b00000000000000000000001110010011;
ROM[16797] <= 32'b00000000011100010010000000100011;
ROM[16798] <= 32'b00000000010000010000000100010011;
ROM[16799] <= 32'b00000001010000000000001110010011;
ROM[16800] <= 32'b01000000011100011000001110110011;
ROM[16801] <= 32'b00000000000000111010000010000011;
ROM[16802] <= 32'b11111111110000010000000100010011;
ROM[16803] <= 32'b00000000000000010010001110000011;
ROM[16804] <= 32'b00000000011100100010000000100011;
ROM[16805] <= 32'b00000000010000100000000100010011;
ROM[16806] <= 32'b00000001010000000000001110010011;
ROM[16807] <= 32'b01000000011100011000001110110011;
ROM[16808] <= 32'b00000000010000111010000110000011;
ROM[16809] <= 32'b00000000100000111010001000000011;
ROM[16810] <= 32'b00000000110000111010001010000011;
ROM[16811] <= 32'b00000001000000111010001100000011;
ROM[16812] <= 32'b00000000000000001000000011100111;
ROM[16813] <= 32'b00000000000000010010000000100011;
ROM[16814] <= 32'b00000000010000010000000100010011;
ROM[16815] <= 32'b00000000000000000000001110010011;
ROM[16816] <= 32'b00000000011100011010000000100011;
ROM[16817] <= 32'b00000000000000011010001110000011;
ROM[16818] <= 32'b00000000011100010010000000100011;
ROM[16819] <= 32'b00000000010000010000000100010011;
ROM[16820] <= 32'b00000000000000100010001110000011;
ROM[16821] <= 32'b00000000011100010010000000100011;
ROM[16822] <= 32'b00000000010000010000000100010011;
ROM[16823] <= 32'b00000000000000010000001110110111;
ROM[16824] <= 32'b01110010100000111000001110010011;
ROM[16825] <= 32'b00000000111000111000001110110011;
ROM[16826] <= 32'b00000000011100010010000000100011;
ROM[16827] <= 32'b00000000010000010000000100010011;
ROM[16828] <= 32'b00000000001100010010000000100011;
ROM[16829] <= 32'b00000000010000010000000100010011;
ROM[16830] <= 32'b00000000010000010010000000100011;
ROM[16831] <= 32'b00000000010000010000000100010011;
ROM[16832] <= 32'b00000000010100010010000000100011;
ROM[16833] <= 32'b00000000010000010000000100010011;
ROM[16834] <= 32'b00000000011000010010000000100011;
ROM[16835] <= 32'b00000000010000010000000100010011;
ROM[16836] <= 32'b00000001010000000000001110010011;
ROM[16837] <= 32'b00000000010000111000001110010011;
ROM[16838] <= 32'b01000000011100010000001110110011;
ROM[16839] <= 32'b00000000011100000000001000110011;
ROM[16840] <= 32'b00000000001000000000000110110011;
ROM[16841] <= 32'b00110101000000000001000011101111;
ROM[16842] <= 32'b11111111110000010000000100010011;
ROM[16843] <= 32'b00000000000000010010001110000011;
ROM[16844] <= 32'b11111111110000010000000100010011;
ROM[16845] <= 32'b00000000000000010010010000000011;
ROM[16846] <= 32'b00000000011101000010001110110011;
ROM[16847] <= 32'b01000000011100000000001110110011;
ROM[16848] <= 32'b00000000000100111000001110010011;
ROM[16849] <= 32'b00000000000000111000101001100011;
ROM[16850] <= 32'b00000000000000010001001110110111;
ROM[16851] <= 32'b10000011100000111000001110010011;
ROM[16852] <= 32'b00000000111000111000001110110011;
ROM[16853] <= 32'b00000000000000111000000011100111;
ROM[16854] <= 32'b00000000000000100010001110000011;
ROM[16855] <= 32'b00000000011100010010000000100011;
ROM[16856] <= 32'b00000000010000010000000100010011;
ROM[16857] <= 32'b00000000000000011010001110000011;
ROM[16858] <= 32'b00000000011100010010000000100011;
ROM[16859] <= 32'b00000000010000010000000100010011;
ROM[16860] <= 32'b00000000000000010000001110110111;
ROM[16861] <= 32'b01111011110000111000001110010011;
ROM[16862] <= 32'b00000000111000111000001110110011;
ROM[16863] <= 32'b00000000011100010010000000100011;
ROM[16864] <= 32'b00000000010000010000000100010011;
ROM[16865] <= 32'b00000000001100010010000000100011;
ROM[16866] <= 32'b00000000010000010000000100010011;
ROM[16867] <= 32'b00000000010000010010000000100011;
ROM[16868] <= 32'b00000000010000010000000100010011;
ROM[16869] <= 32'b00000000010100010010000000100011;
ROM[16870] <= 32'b00000000010000010000000100010011;
ROM[16871] <= 32'b00000000011000010010000000100011;
ROM[16872] <= 32'b00000000010000010000000100010011;
ROM[16873] <= 32'b00000001010000000000001110010011;
ROM[16874] <= 32'b00000000100000111000001110010011;
ROM[16875] <= 32'b01000000011100010000001110110011;
ROM[16876] <= 32'b00000000011100000000001000110011;
ROM[16877] <= 32'b00000000001000000000000110110011;
ROM[16878] <= 32'b00110000110000000001000011101111;
ROM[16879] <= 32'b00000000000000010001001110110111;
ROM[16880] <= 32'b10000000100000111000001110010011;
ROM[16881] <= 32'b00000000111000111000001110110011;
ROM[16882] <= 32'b00000000011100010010000000100011;
ROM[16883] <= 32'b00000000010000010000000100010011;
ROM[16884] <= 32'b00000000001100010010000000100011;
ROM[16885] <= 32'b00000000010000010000000100010011;
ROM[16886] <= 32'b00000000010000010010000000100011;
ROM[16887] <= 32'b00000000010000010000000100010011;
ROM[16888] <= 32'b00000000010100010010000000100011;
ROM[16889] <= 32'b00000000010000010000000100010011;
ROM[16890] <= 32'b00000000011000010010000000100011;
ROM[16891] <= 32'b00000000010000010000000100010011;
ROM[16892] <= 32'b00000001010000000000001110010011;
ROM[16893] <= 32'b00000000010000111000001110010011;
ROM[16894] <= 32'b01000000011100010000001110110011;
ROM[16895] <= 32'b00000000011100000000001000110011;
ROM[16896] <= 32'b00000000001000000000000110110011;
ROM[16897] <= 32'b10010011110011111111000011101111;
ROM[16898] <= 32'b11111111110000010000000100010011;
ROM[16899] <= 32'b00000000000000010010001110000011;
ROM[16900] <= 32'b00000000011101100010000000100011;
ROM[16901] <= 32'b00000000000000011010001110000011;
ROM[16902] <= 32'b00000000011100010010000000100011;
ROM[16903] <= 32'b00000000010000010000000100010011;
ROM[16904] <= 32'b00000000000100000000001110010011;
ROM[16905] <= 32'b11111111110000010000000100010011;
ROM[16906] <= 32'b00000000000000010010010000000011;
ROM[16907] <= 32'b00000000011101000000001110110011;
ROM[16908] <= 32'b00000000011100011010000000100011;
ROM[16909] <= 32'b11101001000111111111000011101111;
ROM[16910] <= 32'b00000000000000000000001110010011;
ROM[16911] <= 32'b00000000011100010010000000100011;
ROM[16912] <= 32'b00000000010000010000000100010011;
ROM[16913] <= 32'b00000001010000000000001110010011;
ROM[16914] <= 32'b01000000011100011000001110110011;
ROM[16915] <= 32'b00000000000000111010000010000011;
ROM[16916] <= 32'b11111111110000010000000100010011;
ROM[16917] <= 32'b00000000000000010010001110000011;
ROM[16918] <= 32'b00000000011100100010000000100011;
ROM[16919] <= 32'b00000000010000100000000100010011;
ROM[16920] <= 32'b00000001010000000000001110010011;
ROM[16921] <= 32'b01000000011100011000001110110011;
ROM[16922] <= 32'b00000000010000111010000110000011;
ROM[16923] <= 32'b00000000100000111010001000000011;
ROM[16924] <= 32'b00000000110000111010001010000011;
ROM[16925] <= 32'b00000001000000111010001100000011;
ROM[16926] <= 32'b00000000000000001000000011100111;
ROM[16927] <= 32'b00000000000000010010000000100011;
ROM[16928] <= 32'b00000000010000010000000100010011;
ROM[16929] <= 32'b00000000101000000000001110010011;
ROM[16930] <= 32'b00000000011100010010000000100011;
ROM[16931] <= 32'b00000000010000010000000100010011;
ROM[16932] <= 32'b00000000000000010001001110110111;
ROM[16933] <= 32'b10001101110000111000001110010011;
ROM[16934] <= 32'b00000000111000111000001110110011;
ROM[16935] <= 32'b00000000011100010010000000100011;
ROM[16936] <= 32'b00000000010000010000000100010011;
ROM[16937] <= 32'b00000000001100010010000000100011;
ROM[16938] <= 32'b00000000010000010000000100010011;
ROM[16939] <= 32'b00000000010000010010000000100011;
ROM[16940] <= 32'b00000000010000010000000100010011;
ROM[16941] <= 32'b00000000010100010010000000100011;
ROM[16942] <= 32'b00000000010000010000000100010011;
ROM[16943] <= 32'b00000000011000010010000000100011;
ROM[16944] <= 32'b00000000010000010000000100010011;
ROM[16945] <= 32'b00000001010000000000001110010011;
ROM[16946] <= 32'b00000000010000111000001110010011;
ROM[16947] <= 32'b01000000011100010000001110110011;
ROM[16948] <= 32'b00000000011100000000001000110011;
ROM[16949] <= 32'b00000000001000000000000110110011;
ROM[16950] <= 32'b00000010100000000001000011101111;
ROM[16951] <= 32'b11111111110000010000000100010011;
ROM[16952] <= 32'b00000000000000010010001110000011;
ROM[16953] <= 32'b00000000011100011010000000100011;
ROM[16954] <= 32'b00000000000000011010001110000011;
ROM[16955] <= 32'b00000000011100010010000000100011;
ROM[16956] <= 32'b00000000010000010000000100010011;
ROM[16957] <= 32'b00000000000000100010001110000011;
ROM[16958] <= 32'b00000000011100010010000000100011;
ROM[16959] <= 32'b00000000010000010000000100010011;
ROM[16960] <= 32'b00000000000000010001001110110111;
ROM[16961] <= 32'b10010100110000111000001110010011;
ROM[16962] <= 32'b00000000111000111000001110110011;
ROM[16963] <= 32'b00000000011100010010000000100011;
ROM[16964] <= 32'b00000000010000010000000100010011;
ROM[16965] <= 32'b00000000001100010010000000100011;
ROM[16966] <= 32'b00000000010000010000000100010011;
ROM[16967] <= 32'b00000000010000010010000000100011;
ROM[16968] <= 32'b00000000010000010000000100010011;
ROM[16969] <= 32'b00000000010100010010000000100011;
ROM[16970] <= 32'b00000000010000010000000100010011;
ROM[16971] <= 32'b00000000011000010010000000100011;
ROM[16972] <= 32'b00000000010000010000000100010011;
ROM[16973] <= 32'b00000001010000000000001110010011;
ROM[16974] <= 32'b00000000100000111000001110010011;
ROM[16975] <= 32'b01000000011100010000001110110011;
ROM[16976] <= 32'b00000000011100000000001000110011;
ROM[16977] <= 32'b00000000001000000000000110110011;
ROM[16978] <= 32'b00111001010100000001000011101111;
ROM[16979] <= 32'b11111111110000010000000100010011;
ROM[16980] <= 32'b00000000000000010010001110000011;
ROM[16981] <= 32'b00000000011101100010000000100011;
ROM[16982] <= 32'b00000000000000011010001110000011;
ROM[16983] <= 32'b00000000011100010010000000100011;
ROM[16984] <= 32'b00000000010000010000000100010011;
ROM[16985] <= 32'b00000000000000010001001110110111;
ROM[16986] <= 32'b10011011000000111000001110010011;
ROM[16987] <= 32'b00000000111000111000001110110011;
ROM[16988] <= 32'b00000000011100010010000000100011;
ROM[16989] <= 32'b00000000010000010000000100010011;
ROM[16990] <= 32'b00000000001100010010000000100011;
ROM[16991] <= 32'b00000000010000010000000100010011;
ROM[16992] <= 32'b00000000010000010010000000100011;
ROM[16993] <= 32'b00000000010000010000000100010011;
ROM[16994] <= 32'b00000000010100010010000000100011;
ROM[16995] <= 32'b00000000010000010000000100010011;
ROM[16996] <= 32'b00000000011000010010000000100011;
ROM[16997] <= 32'b00000000010000010000000100010011;
ROM[16998] <= 32'b00000001010000000000001110010011;
ROM[16999] <= 32'b00000000010000111000001110010011;
ROM[17000] <= 32'b01000000011100010000001110110011;
ROM[17001] <= 32'b00000000011100000000001000110011;
ROM[17002] <= 32'b00000000001000000000000110110011;
ROM[17003] <= 32'b11010000100111111111000011101111;
ROM[17004] <= 32'b11111111110000010000000100010011;
ROM[17005] <= 32'b00000000000000010010001110000011;
ROM[17006] <= 32'b00000000011101100010000000100011;
ROM[17007] <= 32'b00000000000000011010001110000011;
ROM[17008] <= 32'b00000000011100010010000000100011;
ROM[17009] <= 32'b00000000010000010000000100010011;
ROM[17010] <= 32'b00000000000000010001001110110111;
ROM[17011] <= 32'b10100001010000111000001110010011;
ROM[17012] <= 32'b00000000111000111000001110110011;
ROM[17013] <= 32'b00000000011100010010000000100011;
ROM[17014] <= 32'b00000000010000010000000100010011;
ROM[17015] <= 32'b00000000001100010010000000100011;
ROM[17016] <= 32'b00000000010000010000000100010011;
ROM[17017] <= 32'b00000000010000010010000000100011;
ROM[17018] <= 32'b00000000010000010000000100010011;
ROM[17019] <= 32'b00000000010100010010000000100011;
ROM[17020] <= 32'b00000000010000010000000100010011;
ROM[17021] <= 32'b00000000011000010010000000100011;
ROM[17022] <= 32'b00000000010000010000000100010011;
ROM[17023] <= 32'b00000001010000000000001110010011;
ROM[17024] <= 32'b00000000010000111000001110010011;
ROM[17025] <= 32'b01000000011100010000001110110011;
ROM[17026] <= 32'b00000000011100000000001000110011;
ROM[17027] <= 32'b00000000001000000000000110110011;
ROM[17028] <= 32'b00001100010000000010000011101111;
ROM[17029] <= 32'b11111111110000010000000100010011;
ROM[17030] <= 32'b00000000000000010010001110000011;
ROM[17031] <= 32'b00000000011101100010000000100011;
ROM[17032] <= 32'b00000000000000000000001110010011;
ROM[17033] <= 32'b00000000011100010010000000100011;
ROM[17034] <= 32'b00000000010000010000000100010011;
ROM[17035] <= 32'b00000001010000000000001110010011;
ROM[17036] <= 32'b01000000011100011000001110110011;
ROM[17037] <= 32'b00000000000000111010000010000011;
ROM[17038] <= 32'b11111111110000010000000100010011;
ROM[17039] <= 32'b00000000000000010010001110000011;
ROM[17040] <= 32'b00000000011100100010000000100011;
ROM[17041] <= 32'b00000000010000100000000100010011;
ROM[17042] <= 32'b00000001010000000000001110010011;
ROM[17043] <= 32'b01000000011100011000001110110011;
ROM[17044] <= 32'b00000000010000111010000110000011;
ROM[17045] <= 32'b00000000100000111010001000000011;
ROM[17046] <= 32'b00000000110000111010001010000011;
ROM[17047] <= 32'b00000001000000111010001100000011;
ROM[17048] <= 32'b00000000000000001000000011100111;
ROM[17049] <= 32'b00001000010001101010001110000011;
ROM[17050] <= 32'b00000000011100010010000000100011;
ROM[17051] <= 32'b00000000010000010000000100010011;
ROM[17052] <= 32'b00000001110100000000001110010011;
ROM[17053] <= 32'b11111111110000010000000100010011;
ROM[17054] <= 32'b00000000000000010010010000000011;
ROM[17055] <= 32'b00000000011101000010001110110011;
ROM[17056] <= 32'b00000000000000111000101001100011;
ROM[17057] <= 32'b00000000000000010001001110110111;
ROM[17058] <= 32'b10101001100000111000001110010011;
ROM[17059] <= 32'b00000000111000111000001110110011;
ROM[17060] <= 32'b00000000000000111000000011100111;
ROM[17061] <= 32'b00001001000000000000000011101111;
ROM[17062] <= 32'b00001000010001101010001110000011;
ROM[17063] <= 32'b00000000011100010010000000100011;
ROM[17064] <= 32'b00000000010000010000000100010011;
ROM[17065] <= 32'b00000000000100000000001110010011;
ROM[17066] <= 32'b11111111110000010000000100010011;
ROM[17067] <= 32'b00000000000000010010010000000011;
ROM[17068] <= 32'b00000000011101000000001110110011;
ROM[17069] <= 32'b00000000011100010010000000100011;
ROM[17070] <= 32'b00000000010000010000000100010011;
ROM[17071] <= 32'b00000000000000000000001110010011;
ROM[17072] <= 32'b00000000011100010010000000100011;
ROM[17073] <= 32'b00000000010000010000000100010011;
ROM[17074] <= 32'b00000000000000010001001110110111;
ROM[17075] <= 32'b10110001010000111000001110010011;
ROM[17076] <= 32'b00000000111000111000001110110011;
ROM[17077] <= 32'b00000000011100010010000000100011;
ROM[17078] <= 32'b00000000010000010000000100010011;
ROM[17079] <= 32'b00000000001100010010000000100011;
ROM[17080] <= 32'b00000000010000010000000100010011;
ROM[17081] <= 32'b00000000010000010010000000100011;
ROM[17082] <= 32'b00000000010000010000000100010011;
ROM[17083] <= 32'b00000000010100010010000000100011;
ROM[17084] <= 32'b00000000010000010000000100010011;
ROM[17085] <= 32'b00000000011000010010000000100011;
ROM[17086] <= 32'b00000000010000010000000100010011;
ROM[17087] <= 32'b00000001010000000000001110010011;
ROM[17088] <= 32'b00000000100000111000001110010011;
ROM[17089] <= 32'b01000000011100010000001110110011;
ROM[17090] <= 32'b00000000011100000000001000110011;
ROM[17091] <= 32'b00000000001000000000000110110011;
ROM[17092] <= 32'b11011101110111111110000011101111;
ROM[17093] <= 32'b11111111110000010000000100010011;
ROM[17094] <= 32'b00000000000000010010001110000011;
ROM[17095] <= 32'b00000000011101100010000000100011;
ROM[17096] <= 32'b00000111010000000000000011101111;
ROM[17097] <= 32'b00000000000000000000001110010011;
ROM[17098] <= 32'b00000000011100010010000000100011;
ROM[17099] <= 32'b00000000010000010000000100010011;
ROM[17100] <= 32'b00000000000000000000001110010011;
ROM[17101] <= 32'b00000000011100010010000000100011;
ROM[17102] <= 32'b00000000010000010000000100010011;
ROM[17103] <= 32'b00000000000000010001001110110111;
ROM[17104] <= 32'b10111000100000111000001110010011;
ROM[17105] <= 32'b00000000111000111000001110110011;
ROM[17106] <= 32'b00000000011100010010000000100011;
ROM[17107] <= 32'b00000000010000010000000100010011;
ROM[17108] <= 32'b00000000001100010010000000100011;
ROM[17109] <= 32'b00000000010000010000000100010011;
ROM[17110] <= 32'b00000000010000010010000000100011;
ROM[17111] <= 32'b00000000010000010000000100010011;
ROM[17112] <= 32'b00000000010100010010000000100011;
ROM[17113] <= 32'b00000000010000010000000100010011;
ROM[17114] <= 32'b00000000011000010010000000100011;
ROM[17115] <= 32'b00000000010000010000000100010011;
ROM[17116] <= 32'b00000001010000000000001110010011;
ROM[17117] <= 32'b00000000100000111000001110010011;
ROM[17118] <= 32'b01000000011100010000001110110011;
ROM[17119] <= 32'b00000000011100000000001000110011;
ROM[17120] <= 32'b00000000001000000000000110110011;
ROM[17121] <= 32'b11010110100111111110000011101111;
ROM[17122] <= 32'b11111111110000010000000100010011;
ROM[17123] <= 32'b00000000000000010010001110000011;
ROM[17124] <= 32'b00000000011101100010000000100011;
ROM[17125] <= 32'b00000000000000000000001110010011;
ROM[17126] <= 32'b00000000011100010010000000100011;
ROM[17127] <= 32'b00000000010000010000000100010011;
ROM[17128] <= 32'b00000001010000000000001110010011;
ROM[17129] <= 32'b01000000011100011000001110110011;
ROM[17130] <= 32'b00000000000000111010000010000011;
ROM[17131] <= 32'b11111111110000010000000100010011;
ROM[17132] <= 32'b00000000000000010010001110000011;
ROM[17133] <= 32'b00000000011100100010000000100011;
ROM[17134] <= 32'b00000000010000100000000100010011;
ROM[17135] <= 32'b00000001010000000000001110010011;
ROM[17136] <= 32'b01000000011100011000001110110011;
ROM[17137] <= 32'b00000000010000111010000110000011;
ROM[17138] <= 32'b00000000100000111010001000000011;
ROM[17139] <= 32'b00000000110000111010001010000011;
ROM[17140] <= 32'b00000001000000111010001100000011;
ROM[17141] <= 32'b00000000000000001000000011100111;
ROM[17142] <= 32'b00000000000000010010000000100011;
ROM[17143] <= 32'b00000000010000010000000100010011;
ROM[17144] <= 32'b00000000000000010010000000100011;
ROM[17145] <= 32'b00000000010000010000000100010011;
ROM[17146] <= 32'b00000000000000010010000000100011;
ROM[17147] <= 32'b00000000010000010000000100010011;
ROM[17148] <= 32'b00000000000000010010000000100011;
ROM[17149] <= 32'b00000000010000010000000100010011;
ROM[17150] <= 32'b00000000000000010010000000100011;
ROM[17151] <= 32'b00000000010000010000000100010011;
ROM[17152] <= 32'b00000000000000010010000000100011;
ROM[17153] <= 32'b00000000010000010000000100010011;
ROM[17154] <= 32'b00000000000000010010000000100011;
ROM[17155] <= 32'b00000000010000010000000100010011;
ROM[17156] <= 32'b00000000000000010010000000100011;
ROM[17157] <= 32'b00000000010000010000000100010011;
ROM[17158] <= 32'b00000000000000010010000000100011;
ROM[17159] <= 32'b00000000010000010000000100010011;
ROM[17160] <= 32'b00001000000001101010001110000011;
ROM[17161] <= 32'b00000000011100010010000000100011;
ROM[17162] <= 32'b00000000010000010000000100010011;
ROM[17163] <= 32'b00000000000000000000001110010011;
ROM[17164] <= 32'b11111111110000010000000100010011;
ROM[17165] <= 32'b00000000000000010010010000000011;
ROM[17166] <= 32'b00000000011101000010010010110011;
ROM[17167] <= 32'b00000000100000111010010100110011;
ROM[17168] <= 32'b00000000101001001000001110110011;
ROM[17169] <= 32'b00000000000100111000001110010011;
ROM[17170] <= 32'b00000000000100111111001110010011;
ROM[17171] <= 32'b00000000000000111000101001100011;
ROM[17172] <= 32'b00000000000000010001001110110111;
ROM[17173] <= 32'b11000110010000111000001110010011;
ROM[17174] <= 32'b00000000111000111000001110110011;
ROM[17175] <= 32'b00000000000000111000000011100111;
ROM[17176] <= 32'b00001110000000000000000011101111;
ROM[17177] <= 32'b00001000010001101010001110000011;
ROM[17178] <= 32'b00000000011100010010000000100011;
ROM[17179] <= 32'b00000000010000010000000100010011;
ROM[17180] <= 32'b00000000000000000000001110010011;
ROM[17181] <= 32'b11111111110000010000000100010011;
ROM[17182] <= 32'b00000000000000010010010000000011;
ROM[17183] <= 32'b00000000011101000010010010110011;
ROM[17184] <= 32'b00000000100000111010010100110011;
ROM[17185] <= 32'b00000000101001001000001110110011;
ROM[17186] <= 32'b00000000000100111000001110010011;
ROM[17187] <= 32'b00000000000100111111001110010011;
ROM[17188] <= 32'b01000000011100000000001110110011;
ROM[17189] <= 32'b00000000000100111000001110010011;
ROM[17190] <= 32'b00000000000000111000101001100011;
ROM[17191] <= 32'b00000000000000010001001110110111;
ROM[17192] <= 32'b11001011000000111000001110010011;
ROM[17193] <= 32'b00000000111000111000001110110011;
ROM[17194] <= 32'b00000000000000111000000011100111;
ROM[17195] <= 32'b00001001000000000000000011101111;
ROM[17196] <= 32'b00001000010001101010001110000011;
ROM[17197] <= 32'b00000000011100010010000000100011;
ROM[17198] <= 32'b00000000010000010000000100010011;
ROM[17199] <= 32'b00000000000100000000001110010011;
ROM[17200] <= 32'b11111111110000010000000100010011;
ROM[17201] <= 32'b00000000000000010010010000000011;
ROM[17202] <= 32'b01000000011101000000001110110011;
ROM[17203] <= 32'b00000000011100010010000000100011;
ROM[17204] <= 32'b00000000010000010000000100010011;
ROM[17205] <= 32'b00000010011100000000001110010011;
ROM[17206] <= 32'b00000000011100010010000000100011;
ROM[17207] <= 32'b00000000010000010000000100010011;
ROM[17208] <= 32'b00000000000000010001001110110111;
ROM[17209] <= 32'b11010010110000111000001110010011;
ROM[17210] <= 32'b00000000111000111000001110110011;
ROM[17211] <= 32'b00000000011100010010000000100011;
ROM[17212] <= 32'b00000000010000010000000100010011;
ROM[17213] <= 32'b00000000001100010010000000100011;
ROM[17214] <= 32'b00000000010000010000000100010011;
ROM[17215] <= 32'b00000000010000010010000000100011;
ROM[17216] <= 32'b00000000010000010000000100010011;
ROM[17217] <= 32'b00000000010100010010000000100011;
ROM[17218] <= 32'b00000000010000010000000100010011;
ROM[17219] <= 32'b00000000011000010010000000100011;
ROM[17220] <= 32'b00000000010000010000000100010011;
ROM[17221] <= 32'b00000001010000000000001110010011;
ROM[17222] <= 32'b00000000100000111000001110010011;
ROM[17223] <= 32'b01000000011100010000001110110011;
ROM[17224] <= 32'b00000000011100000000001000110011;
ROM[17225] <= 32'b00000000001000000000000110110011;
ROM[17226] <= 32'b10111100010111111110000011101111;
ROM[17227] <= 32'b11111111110000010000000100010011;
ROM[17228] <= 32'b00000000000000010010001110000011;
ROM[17229] <= 32'b00000000011101100010000000100011;
ROM[17230] <= 32'b00000000010000000000000011101111;
ROM[17231] <= 32'b00001000110000000000000011101111;
ROM[17232] <= 32'b00001000010001101010001110000011;
ROM[17233] <= 32'b00000000011100010010000000100011;
ROM[17234] <= 32'b00000000010000010000000100010011;
ROM[17235] <= 32'b00001000000001101010001110000011;
ROM[17236] <= 32'b00000000011100010010000000100011;
ROM[17237] <= 32'b00000000010000010000000100010011;
ROM[17238] <= 32'b00000000000100000000001110010011;
ROM[17239] <= 32'b11111111110000010000000100010011;
ROM[17240] <= 32'b00000000000000010010010000000011;
ROM[17241] <= 32'b01000000011101000000001110110011;
ROM[17242] <= 32'b00000000011100010010000000100011;
ROM[17243] <= 32'b00000000010000010000000100010011;
ROM[17244] <= 32'b00000000000000010001001110110111;
ROM[17245] <= 32'b11011011110000111000001110010011;
ROM[17246] <= 32'b00000000111000111000001110110011;
ROM[17247] <= 32'b00000000011100010010000000100011;
ROM[17248] <= 32'b00000000010000010000000100010011;
ROM[17249] <= 32'b00000000001100010010000000100011;
ROM[17250] <= 32'b00000000010000010000000100010011;
ROM[17251] <= 32'b00000000010000010010000000100011;
ROM[17252] <= 32'b00000000010000010000000100010011;
ROM[17253] <= 32'b00000000010100010010000000100011;
ROM[17254] <= 32'b00000000010000010000000100010011;
ROM[17255] <= 32'b00000000011000010010000000100011;
ROM[17256] <= 32'b00000000010000010000000100010011;
ROM[17257] <= 32'b00000001010000000000001110010011;
ROM[17258] <= 32'b00000000100000111000001110010011;
ROM[17259] <= 32'b01000000011100010000001110110011;
ROM[17260] <= 32'b00000000011100000000001000110011;
ROM[17261] <= 32'b00000000001000000000000110110011;
ROM[17262] <= 32'b10110011010111111110000011101111;
ROM[17263] <= 32'b11111111110000010000000100010011;
ROM[17264] <= 32'b00000000000000010010001110000011;
ROM[17265] <= 32'b00000000011101100010000000100011;
ROM[17266] <= 32'b00001000010001101010001110000011;
ROM[17267] <= 32'b00000000011100010010000000100011;
ROM[17268] <= 32'b00000000010000010000000100010011;
ROM[17269] <= 32'b00000000101000000000001110010011;
ROM[17270] <= 32'b00000000011100010010000000100011;
ROM[17271] <= 32'b00000000010000010000000100010011;
ROM[17272] <= 32'b00000000000000010001001110110111;
ROM[17273] <= 32'b11100010110000111000001110010011;
ROM[17274] <= 32'b00000000111000111000001110110011;
ROM[17275] <= 32'b00000000011100010010000000100011;
ROM[17276] <= 32'b00000000010000010000000100010011;
ROM[17277] <= 32'b00000000001100010010000000100011;
ROM[17278] <= 32'b00000000010000010000000100010011;
ROM[17279] <= 32'b00000000010000010010000000100011;
ROM[17280] <= 32'b00000000010000010000000100010011;
ROM[17281] <= 32'b00000000010100010010000000100011;
ROM[17282] <= 32'b00000000010000010000000100010011;
ROM[17283] <= 32'b00000000011000010010000000100011;
ROM[17284] <= 32'b00000000010000010000000100010011;
ROM[17285] <= 32'b00000001010000000000001110010011;
ROM[17286] <= 32'b00000000100000111000001110010011;
ROM[17287] <= 32'b01000000011100010000001110110011;
ROM[17288] <= 32'b00000000011100000000001000110011;
ROM[17289] <= 32'b00000000001000000000000110110011;
ROM[17290] <= 32'b10101010110011111000000011101111;
ROM[17291] <= 32'b00000000100000000000001110010011;
ROM[17292] <= 32'b00000000011100010010000000100011;
ROM[17293] <= 32'b00000000010000010000000100010011;
ROM[17294] <= 32'b00000000000000010001001110110111;
ROM[17295] <= 32'b11101000010000111000001110010011;
ROM[17296] <= 32'b00000000111000111000001110110011;
ROM[17297] <= 32'b00000000011100010010000000100011;
ROM[17298] <= 32'b00000000010000010000000100010011;
ROM[17299] <= 32'b00000000001100010010000000100011;
ROM[17300] <= 32'b00000000010000010000000100010011;
ROM[17301] <= 32'b00000000010000010010000000100011;
ROM[17302] <= 32'b00000000010000010000000100010011;
ROM[17303] <= 32'b00000000010100010010000000100011;
ROM[17304] <= 32'b00000000010000010000000100010011;
ROM[17305] <= 32'b00000000011000010010000000100011;
ROM[17306] <= 32'b00000000010000010000000100010011;
ROM[17307] <= 32'b00000001010000000000001110010011;
ROM[17308] <= 32'b00000000100000111000001110010011;
ROM[17309] <= 32'b01000000011100010000001110110011;
ROM[17310] <= 32'b00000000011100000000001000110011;
ROM[17311] <= 32'b00000000001000000000000110110011;
ROM[17312] <= 32'b10100101010011111000000011101111;
ROM[17313] <= 32'b00001000000001101010001110000011;
ROM[17314] <= 32'b00000000011100010010000000100011;
ROM[17315] <= 32'b00000000010000010000000100010011;
ROM[17316] <= 32'b00000000010000000000001110010011;
ROM[17317] <= 32'b00000000011100010010000000100011;
ROM[17318] <= 32'b00000000010000010000000100010011;
ROM[17319] <= 32'b00000000000000010001001110110111;
ROM[17320] <= 32'b11101110100000111000001110010011;
ROM[17321] <= 32'b00000000111000111000001110110011;
ROM[17322] <= 32'b00000000011100010010000000100011;
ROM[17323] <= 32'b00000000010000010000000100010011;
ROM[17324] <= 32'b00000000001100010010000000100011;
ROM[17325] <= 32'b00000000010000010000000100010011;
ROM[17326] <= 32'b00000000010000010010000000100011;
ROM[17327] <= 32'b00000000010000010000000100010011;
ROM[17328] <= 32'b00000000010100010010000000100011;
ROM[17329] <= 32'b00000000010000010000000100010011;
ROM[17330] <= 32'b00000000011000010010000000100011;
ROM[17331] <= 32'b00000000010000010000000100010011;
ROM[17332] <= 32'b00000001010000000000001110010011;
ROM[17333] <= 32'b00000000100000111000001110010011;
ROM[17334] <= 32'b01000000011100010000001110110011;
ROM[17335] <= 32'b00000000011100000000001000110011;
ROM[17336] <= 32'b00000000001000000000000110110011;
ROM[17337] <= 32'b11000001010011111000000011101111;
ROM[17338] <= 32'b11111111110000010000000100010011;
ROM[17339] <= 32'b00000000000000010010001110000011;
ROM[17340] <= 32'b11111111110000010000000100010011;
ROM[17341] <= 32'b00000000000000010010010000000011;
ROM[17342] <= 32'b00000000011101000000001110110011;
ROM[17343] <= 32'b00000000011100011010000000100011;
ROM[17344] <= 32'b00001000000001101010001110000011;
ROM[17345] <= 32'b00000000011100010010000000100011;
ROM[17346] <= 32'b00000000010000010000000100010011;
ROM[17347] <= 32'b00000000001100000000001110010011;
ROM[17348] <= 32'b11111111110000010000000100010011;
ROM[17349] <= 32'b00000000000000010010010000000011;
ROM[17350] <= 32'b00000000011101000111001110110011;
ROM[17351] <= 32'b00000000011100011010010000100011;
ROM[17352] <= 32'b00000000000000000000001110010011;
ROM[17353] <= 32'b00000000011100011010001000100011;
ROM[17354] <= 32'b00000000010000011010001110000011;
ROM[17355] <= 32'b00000000011100010010000000100011;
ROM[17356] <= 32'b00000000010000010000000100010011;
ROM[17357] <= 32'b00000000100000000000001110010011;
ROM[17358] <= 32'b11111111110000010000000100010011;
ROM[17359] <= 32'b00000000000000010010010000000011;
ROM[17360] <= 32'b00000000011101000010001110110011;
ROM[17361] <= 32'b01000000011100000000001110110011;
ROM[17362] <= 32'b00000000000100111000001110010011;
ROM[17363] <= 32'b00000000000000111000101001100011;
ROM[17364] <= 32'b00000000000000010001001110110111;
ROM[17365] <= 32'b01011111110000111000001110010011;
ROM[17366] <= 32'b00000000111000111000001110110011;
ROM[17367] <= 32'b00000000000000111000000011100111;
ROM[17368] <= 32'b00000000010000011010001110000011;
ROM[17369] <= 32'b00000000011100010010000000100011;
ROM[17370] <= 32'b00000000010000010000000100010011;
ROM[17371] <= 32'b00000000010000000000001110010011;
ROM[17372] <= 32'b00000000011100010010000000100011;
ROM[17373] <= 32'b00000000010000010000000100010011;
ROM[17374] <= 32'b00000000000000010001001110110111;
ROM[17375] <= 32'b11111100010000111000001110010011;
ROM[17376] <= 32'b00000000111000111000001110110011;
ROM[17377] <= 32'b00000000011100010010000000100011;
ROM[17378] <= 32'b00000000010000010000000100010011;
ROM[17379] <= 32'b00000000001100010010000000100011;
ROM[17380] <= 32'b00000000010000010000000100010011;
ROM[17381] <= 32'b00000000010000010010000000100011;
ROM[17382] <= 32'b00000000010000010000000100010011;
ROM[17383] <= 32'b00000000010100010010000000100011;
ROM[17384] <= 32'b00000000010000010000000100010011;
ROM[17385] <= 32'b00000000011000010010000000100011;
ROM[17386] <= 32'b00000000010000010000000100010011;
ROM[17387] <= 32'b00000001010000000000001110010011;
ROM[17388] <= 32'b00000000100000111000001110010011;
ROM[17389] <= 32'b01000000011100010000001110110011;
ROM[17390] <= 32'b00000000011100000000001000110011;
ROM[17391] <= 32'b00000000001000000000000110110011;
ROM[17392] <= 32'b10010001010011111000000011101111;
ROM[17393] <= 32'b11111111110000010000000100010011;
ROM[17394] <= 32'b00000000000000010010001110000011;
ROM[17395] <= 32'b00000000011100011010011000100011;
ROM[17396] <= 32'b00000000000000011010001110000011;
ROM[17397] <= 32'b00000000011100010010000000100011;
ROM[17398] <= 32'b00000000010000010000000100010011;
ROM[17399] <= 32'b00000000010000000000001110010011;
ROM[17400] <= 32'b00000000011100010010000000100011;
ROM[17401] <= 32'b00000000010000010000000100010011;
ROM[17402] <= 32'b00000000000000010001001110110111;
ROM[17403] <= 32'b00000011010000111000001110010011;
ROM[17404] <= 32'b00000000111000111000001110110011;
ROM[17405] <= 32'b00000000011100010010000000100011;
ROM[17406] <= 32'b00000000010000010000000100010011;
ROM[17407] <= 32'b00000000001100010010000000100011;
ROM[17408] <= 32'b00000000010000010000000100010011;
ROM[17409] <= 32'b00000000010000010010000000100011;
ROM[17410] <= 32'b00000000010000010000000100010011;
ROM[17411] <= 32'b00000000010100010010000000100011;
ROM[17412] <= 32'b00000000010000010000000100010011;
ROM[17413] <= 32'b00000000011000010010000000100011;
ROM[17414] <= 32'b00000000010000010000000100010011;
ROM[17415] <= 32'b00000001010000000000001110010011;
ROM[17416] <= 32'b00000000100000111000001110010011;
ROM[17417] <= 32'b01000000011100010000001110110011;
ROM[17418] <= 32'b00000000011100000000001000110011;
ROM[17419] <= 32'b00000000001000000000000110110011;
ROM[17420] <= 32'b10001010010011111000000011101111;
ROM[17421] <= 32'b11111111110000010000000100010011;
ROM[17422] <= 32'b00000000000000010010001110000011;
ROM[17423] <= 32'b00000000011100011010100000100011;
ROM[17424] <= 32'b00000000100000011010001110000011;
ROM[17425] <= 32'b00000000011100010010000000100011;
ROM[17426] <= 32'b00000000010000010000000100010011;
ROM[17427] <= 32'b00000000000000000000001110010011;
ROM[17428] <= 32'b11111111110000010000000100010011;
ROM[17429] <= 32'b00000000000000010010010000000011;
ROM[17430] <= 32'b00000000011101000010010010110011;
ROM[17431] <= 32'b00000000100000111010010100110011;
ROM[17432] <= 32'b00000000101001001000001110110011;
ROM[17433] <= 32'b00000000000100111000001110010011;
ROM[17434] <= 32'b00000000000100111111001110010011;
ROM[17435] <= 32'b00000000000000111000101001100011;
ROM[17436] <= 32'b00000000000000010001001110110111;
ROM[17437] <= 32'b00001000010000111000001110010011;
ROM[17438] <= 32'b00000000111000111000001110110011;
ROM[17439] <= 32'b00000000000000111000000011100111;
ROM[17440] <= 32'b00001111110000000000000011101111;
ROM[17441] <= 32'b00000001100000000000001110010011;
ROM[17442] <= 32'b00000000011100010010000000100011;
ROM[17443] <= 32'b00000000010000010000000100010011;
ROM[17444] <= 32'b00000000000000010001001110110111;
ROM[17445] <= 32'b00001101110000111000001110010011;
ROM[17446] <= 32'b00000000111000111000001110110011;
ROM[17447] <= 32'b00000000011100010010000000100011;
ROM[17448] <= 32'b00000000010000010000000100010011;
ROM[17449] <= 32'b00000000001100010010000000100011;
ROM[17450] <= 32'b00000000010000010000000100010011;
ROM[17451] <= 32'b00000000010000010010000000100011;
ROM[17452] <= 32'b00000000010000010000000100010011;
ROM[17453] <= 32'b00000000010100010010000000100011;
ROM[17454] <= 32'b00000000010000010000000100010011;
ROM[17455] <= 32'b00000000011000010010000000100011;
ROM[17456] <= 32'b00000000010000010000000100010011;
ROM[17457] <= 32'b00000001010000000000001110010011;
ROM[17458] <= 32'b00000000010000111000001110010011;
ROM[17459] <= 32'b01000000011100010000001110110011;
ROM[17460] <= 32'b00000000011100000000001000110011;
ROM[17461] <= 32'b00000000001000000000000110110011;
ROM[17462] <= 32'b11010010010011111000000011101111;
ROM[17463] <= 32'b00000000000100000000001110010011;
ROM[17464] <= 32'b11111111110000010000000100010011;
ROM[17465] <= 32'b00000000000000010010010000000011;
ROM[17466] <= 32'b01000000011101000000001110110011;
ROM[17467] <= 32'b00000000011100011010111000100011;
ROM[17468] <= 32'b00000001000000011010001110000011;
ROM[17469] <= 32'b00000000011100010010000000100011;
ROM[17470] <= 32'b00000000010000010000000100010011;
ROM[17471] <= 32'b00000111110001101010001110000011;
ROM[17472] <= 32'b11111111110000010000000100010011;
ROM[17473] <= 32'b00000000000000010010010000000011;
ROM[17474] <= 32'b00000000011101000000001110110011;
ROM[17475] <= 32'b00000000000000111000001100010011;
ROM[17476] <= 32'b00000000110100110000010000110011;
ROM[17477] <= 32'b00000000000001000010001110000011;
ROM[17478] <= 32'b00000000011100010010000000100011;
ROM[17479] <= 32'b00000000010000010000000100010011;
ROM[17480] <= 32'b00000001110000011010001110000011;
ROM[17481] <= 32'b11111111110000010000000100010011;
ROM[17482] <= 32'b00000000000000010010010000000011;
ROM[17483] <= 32'b00000000011101000111001110110011;
ROM[17484] <= 32'b00000010011100011010000000100011;
ROM[17485] <= 32'b00000001000000011010001110000011;
ROM[17486] <= 32'b00000000011100010010000000100011;
ROM[17487] <= 32'b00000000010000010000000100010011;
ROM[17488] <= 32'b00000111110001101010001110000011;
ROM[17489] <= 32'b11111111110000010000000100010011;
ROM[17490] <= 32'b00000000000000010010010000000011;
ROM[17491] <= 32'b00000000011101000000001110110011;
ROM[17492] <= 32'b00000000011100010010000000100011;
ROM[17493] <= 32'b00000000010000010000000100010011;
ROM[17494] <= 32'b00000010000000011010001110000011;
ROM[17495] <= 32'b00000000011101100010000000100011;
ROM[17496] <= 32'b11111111110000010000000100010011;
ROM[17497] <= 32'b00000000000000010010001110000011;
ROM[17498] <= 32'b00000000000000111000001100010011;
ROM[17499] <= 32'b00000000000001100010001110000011;
ROM[17500] <= 32'b00000000110100110000010000110011;
ROM[17501] <= 32'b00000000011101000010000000100011;
ROM[17502] <= 32'b01000100000000000000000011101111;
ROM[17503] <= 32'b00000000100000011010001110000011;
ROM[17504] <= 32'b00000000011100010010000000100011;
ROM[17505] <= 32'b00000000010000010000000100010011;
ROM[17506] <= 32'b00000000000100000000001110010011;
ROM[17507] <= 32'b11111111110000010000000100010011;
ROM[17508] <= 32'b00000000000000010010010000000011;
ROM[17509] <= 32'b00000000011101000010010010110011;
ROM[17510] <= 32'b00000000100000111010010100110011;
ROM[17511] <= 32'b00000000101001001000001110110011;
ROM[17512] <= 32'b00000000000100111000001110010011;
ROM[17513] <= 32'b00000000000100111111001110010011;
ROM[17514] <= 32'b00000000000000111000101001100011;
ROM[17515] <= 32'b00000000000000010001001110110111;
ROM[17516] <= 32'b00011100000000111000001110010011;
ROM[17517] <= 32'b00000000111000111000001110110011;
ROM[17518] <= 32'b00000000000000111000000011100111;
ROM[17519] <= 32'b00011001100000000000000011101111;
ROM[17520] <= 32'b00000001100000000000001110010011;
ROM[17521] <= 32'b00000000011100010010000000100011;
ROM[17522] <= 32'b00000000010000010000000100010011;
ROM[17523] <= 32'b00000000000000010001001110110111;
ROM[17524] <= 32'b00100001100000111000001110010011;
ROM[17525] <= 32'b00000000111000111000001110110011;
ROM[17526] <= 32'b00000000011100010010000000100011;
ROM[17527] <= 32'b00000000010000010000000100010011;
ROM[17528] <= 32'b00000000001100010010000000100011;
ROM[17529] <= 32'b00000000010000010000000100010011;
ROM[17530] <= 32'b00000000010000010010000000100011;
ROM[17531] <= 32'b00000000010000010000000100010011;
ROM[17532] <= 32'b00000000010100010010000000100011;
ROM[17533] <= 32'b00000000010000010000000100010011;
ROM[17534] <= 32'b00000000011000010010000000100011;
ROM[17535] <= 32'b00000000010000010000000100010011;
ROM[17536] <= 32'b00000001010000000000001110010011;
ROM[17537] <= 32'b00000000010000111000001110010011;
ROM[17538] <= 32'b01000000011100010000001110110011;
ROM[17539] <= 32'b00000000011100000000001000110011;
ROM[17540] <= 32'b00000000001000000000000110110011;
ROM[17541] <= 32'b10111110100011111000000011101111;
ROM[17542] <= 32'b00000001000000000000001110010011;
ROM[17543] <= 32'b00000000011100010010000000100011;
ROM[17544] <= 32'b00000000010000010000000100010011;
ROM[17545] <= 32'b00000000000000010001001110110111;
ROM[17546] <= 32'b00100111000000111000001110010011;
ROM[17547] <= 32'b00000000111000111000001110110011;
ROM[17548] <= 32'b00000000011100010010000000100011;
ROM[17549] <= 32'b00000000010000010000000100010011;
ROM[17550] <= 32'b00000000001100010010000000100011;
ROM[17551] <= 32'b00000000010000010000000100010011;
ROM[17552] <= 32'b00000000010000010010000000100011;
ROM[17553] <= 32'b00000000010000010000000100010011;
ROM[17554] <= 32'b00000000010100010010000000100011;
ROM[17555] <= 32'b00000000010000010000000100010011;
ROM[17556] <= 32'b00000000011000010010000000100011;
ROM[17557] <= 32'b00000000010000010000000100010011;
ROM[17558] <= 32'b00000001010000000000001110010011;
ROM[17559] <= 32'b00000000010000111000001110010011;
ROM[17560] <= 32'b01000000011100010000001110110011;
ROM[17561] <= 32'b00000000011100000000001000110011;
ROM[17562] <= 32'b00000000001000000000000110110011;
ROM[17563] <= 32'b10111001000011111000000011101111;
ROM[17564] <= 32'b11111111110000010000000100010011;
ROM[17565] <= 32'b00000000000000010010001110000011;
ROM[17566] <= 32'b11111111110000010000000100010011;
ROM[17567] <= 32'b00000000000000010010010000000011;
ROM[17568] <= 32'b01000000011101000000001110110011;
ROM[17569] <= 32'b00000000011100011010101000100011;
ROM[17570] <= 32'b00000000000000000000001110010011;
ROM[17571] <= 32'b00000000011100010010000000100011;
ROM[17572] <= 32'b00000000010000010000000100010011;
ROM[17573] <= 32'b00000001010000011010001110000011;
ROM[17574] <= 32'b11111111110000010000000100010011;
ROM[17575] <= 32'b00000000000000010010010000000011;
ROM[17576] <= 32'b01000000011101000000001110110011;
ROM[17577] <= 32'b00000000011100011010111000100011;
ROM[17578] <= 32'b00000001110000011010001110000011;
ROM[17579] <= 32'b00000000011100010010000000100011;
ROM[17580] <= 32'b00000000010000010000000100010011;
ROM[17581] <= 32'b00000000000100000000001110010011;
ROM[17582] <= 32'b11111111110000010000000100010011;
ROM[17583] <= 32'b00000000000000010010010000000011;
ROM[17584] <= 32'b01000000011101000000001110110011;
ROM[17585] <= 32'b00000000011100011010111000100011;
ROM[17586] <= 32'b00000001000000011010001110000011;
ROM[17587] <= 32'b00000000011100010010000000100011;
ROM[17588] <= 32'b00000000010000010000000100010011;
ROM[17589] <= 32'b00000111110001101010001110000011;
ROM[17590] <= 32'b11111111110000010000000100010011;
ROM[17591] <= 32'b00000000000000010010010000000011;
ROM[17592] <= 32'b00000000011101000000001110110011;
ROM[17593] <= 32'b00000000000000111000001100010011;
ROM[17594] <= 32'b00000000110100110000010000110011;
ROM[17595] <= 32'b00000000000001000010001110000011;
ROM[17596] <= 32'b00000000011100010010000000100011;
ROM[17597] <= 32'b00000000010000010000000100010011;
ROM[17598] <= 32'b00000001110000011010001110000011;
ROM[17599] <= 32'b11111111110000010000000100010011;
ROM[17600] <= 32'b00000000000000010010010000000011;
ROM[17601] <= 32'b00000000011101000111001110110011;
ROM[17602] <= 32'b00000010011100011010000000100011;
ROM[17603] <= 32'b00000001000000011010001110000011;
ROM[17604] <= 32'b00000000011100010010000000100011;
ROM[17605] <= 32'b00000000010000010000000100010011;
ROM[17606] <= 32'b00000111110001101010001110000011;
ROM[17607] <= 32'b11111111110000010000000100010011;
ROM[17608] <= 32'b00000000000000010010010000000011;
ROM[17609] <= 32'b00000000011101000000001110110011;
ROM[17610] <= 32'b00000000011100010010000000100011;
ROM[17611] <= 32'b00000000010000010000000100010011;
ROM[17612] <= 32'b00000010000000011010001110000011;
ROM[17613] <= 32'b00000000011101100010000000100011;
ROM[17614] <= 32'b11111111110000010000000100010011;
ROM[17615] <= 32'b00000000000000010010001110000011;
ROM[17616] <= 32'b00000000000000111000001100010011;
ROM[17617] <= 32'b00000000000001100010001110000011;
ROM[17618] <= 32'b00000000110100110000010000110011;
ROM[17619] <= 32'b00000000011101000010000000100011;
ROM[17620] <= 32'b00100110100000000000000011101111;
ROM[17621] <= 32'b00000000100000011010001110000011;
ROM[17622] <= 32'b00000000011100010010000000100011;
ROM[17623] <= 32'b00000000010000010000000100010011;
ROM[17624] <= 32'b00000000001000000000001110010011;
ROM[17625] <= 32'b11111111110000010000000100010011;
ROM[17626] <= 32'b00000000000000010010010000000011;
ROM[17627] <= 32'b00000000011101000010010010110011;
ROM[17628] <= 32'b00000000100000111010010100110011;
ROM[17629] <= 32'b00000000101001001000001110110011;
ROM[17630] <= 32'b00000000000100111000001110010011;
ROM[17631] <= 32'b00000000000100111111001110010011;
ROM[17632] <= 32'b00000000000000111000101001100011;
ROM[17633] <= 32'b00000000000000010001001110110111;
ROM[17634] <= 32'b00111001100000111000001110010011;
ROM[17635] <= 32'b00000000111000111000001110110011;
ROM[17636] <= 32'b00000000000000111000000011100111;
ROM[17637] <= 32'b00011001100000000000000011101111;
ROM[17638] <= 32'b00000001000000000000001110010011;
ROM[17639] <= 32'b00000000011100010010000000100011;
ROM[17640] <= 32'b00000000010000010000000100010011;
ROM[17641] <= 32'b00000000000000010001001110110111;
ROM[17642] <= 32'b00111111000000111000001110010011;
ROM[17643] <= 32'b00000000111000111000001110110011;
ROM[17644] <= 32'b00000000011100010010000000100011;
ROM[17645] <= 32'b00000000010000010000000100010011;
ROM[17646] <= 32'b00000000001100010010000000100011;
ROM[17647] <= 32'b00000000010000010000000100010011;
ROM[17648] <= 32'b00000000010000010010000000100011;
ROM[17649] <= 32'b00000000010000010000000100010011;
ROM[17650] <= 32'b00000000010100010010000000100011;
ROM[17651] <= 32'b00000000010000010000000100010011;
ROM[17652] <= 32'b00000000011000010010000000100011;
ROM[17653] <= 32'b00000000010000010000000100010011;
ROM[17654] <= 32'b00000001010000000000001110010011;
ROM[17655] <= 32'b00000000010000111000001110010011;
ROM[17656] <= 32'b01000000011100010000001110110011;
ROM[17657] <= 32'b00000000011100000000001000110011;
ROM[17658] <= 32'b00000000001000000000000110110011;
ROM[17659] <= 32'b10100001000011111000000011101111;
ROM[17660] <= 32'b00000000100000000000001110010011;
ROM[17661] <= 32'b00000000011100010010000000100011;
ROM[17662] <= 32'b00000000010000010000000100010011;
ROM[17663] <= 32'b00000000000000010001001110110111;
ROM[17664] <= 32'b01000100100000111000001110010011;
ROM[17665] <= 32'b00000000111000111000001110110011;
ROM[17666] <= 32'b00000000011100010010000000100011;
ROM[17667] <= 32'b00000000010000010000000100010011;
ROM[17668] <= 32'b00000000001100010010000000100011;
ROM[17669] <= 32'b00000000010000010000000100010011;
ROM[17670] <= 32'b00000000010000010010000000100011;
ROM[17671] <= 32'b00000000010000010000000100010011;
ROM[17672] <= 32'b00000000010100010010000000100011;
ROM[17673] <= 32'b00000000010000010000000100010011;
ROM[17674] <= 32'b00000000011000010010000000100011;
ROM[17675] <= 32'b00000000010000010000000100010011;
ROM[17676] <= 32'b00000001010000000000001110010011;
ROM[17677] <= 32'b00000000010000111000001110010011;
ROM[17678] <= 32'b01000000011100010000001110110011;
ROM[17679] <= 32'b00000000011100000000001000110011;
ROM[17680] <= 32'b00000000001000000000000110110011;
ROM[17681] <= 32'b10011011100011111000000011101111;
ROM[17682] <= 32'b11111111110000010000000100010011;
ROM[17683] <= 32'b00000000000000010010001110000011;
ROM[17684] <= 32'b11111111110000010000000100010011;
ROM[17685] <= 32'b00000000000000010010010000000011;
ROM[17686] <= 32'b01000000011101000000001110110011;
ROM[17687] <= 32'b00000000011100011010110000100011;
ROM[17688] <= 32'b00000000000000000000001110010011;
ROM[17689] <= 32'b00000000011100010010000000100011;
ROM[17690] <= 32'b00000000010000010000000100010011;
ROM[17691] <= 32'b00000001100000011010001110000011;
ROM[17692] <= 32'b11111111110000010000000100010011;
ROM[17693] <= 32'b00000000000000010010010000000011;
ROM[17694] <= 32'b01000000011101000000001110110011;
ROM[17695] <= 32'b00000000011100011010111000100011;
ROM[17696] <= 32'b00000001110000011010001110000011;
ROM[17697] <= 32'b00000000011100010010000000100011;
ROM[17698] <= 32'b00000000010000010000000100010011;
ROM[17699] <= 32'b00000000000100000000001110010011;
ROM[17700] <= 32'b11111111110000010000000100010011;
ROM[17701] <= 32'b00000000000000010010010000000011;
ROM[17702] <= 32'b01000000011101000000001110110011;
ROM[17703] <= 32'b00000000011100011010111000100011;
ROM[17704] <= 32'b00000001000000011010001110000011;
ROM[17705] <= 32'b00000000011100010010000000100011;
ROM[17706] <= 32'b00000000010000010000000100010011;
ROM[17707] <= 32'b00000111110001101010001110000011;
ROM[17708] <= 32'b11111111110000010000000100010011;
ROM[17709] <= 32'b00000000000000010010010000000011;
ROM[17710] <= 32'b00000000011101000000001110110011;
ROM[17711] <= 32'b00000000000000111000001100010011;
ROM[17712] <= 32'b00000000110100110000010000110011;
ROM[17713] <= 32'b00000000000001000010001110000011;
ROM[17714] <= 32'b00000000011100010010000000100011;
ROM[17715] <= 32'b00000000010000010000000100010011;
ROM[17716] <= 32'b00000001110000011010001110000011;
ROM[17717] <= 32'b11111111110000010000000100010011;
ROM[17718] <= 32'b00000000000000010010010000000011;
ROM[17719] <= 32'b00000000011101000111001110110011;
ROM[17720] <= 32'b00000010011100011010000000100011;
ROM[17721] <= 32'b00000001000000011010001110000011;
ROM[17722] <= 32'b00000000011100010010000000100011;
ROM[17723] <= 32'b00000000010000010000000100010011;
ROM[17724] <= 32'b00000111110001101010001110000011;
ROM[17725] <= 32'b11111111110000010000000100010011;
ROM[17726] <= 32'b00000000000000010010010000000011;
ROM[17727] <= 32'b00000000011101000000001110110011;
ROM[17728] <= 32'b00000000011100010010000000100011;
ROM[17729] <= 32'b00000000010000010000000100010011;
ROM[17730] <= 32'b00000010000000011010001110000011;
ROM[17731] <= 32'b00000000011101100010000000100011;
ROM[17732] <= 32'b11111111110000010000000100010011;
ROM[17733] <= 32'b00000000000000010010001110000011;
ROM[17734] <= 32'b00000000000000111000001100010011;
ROM[17735] <= 32'b00000000000001100010001110000011;
ROM[17736] <= 32'b00000000110100110000010000110011;
ROM[17737] <= 32'b00000000011101000010000000100011;
ROM[17738] <= 32'b00001001000000000000000011101111;
ROM[17739] <= 32'b00000001000000011010001110000011;
ROM[17740] <= 32'b00000000011100010010000000100011;
ROM[17741] <= 32'b00000000010000010000000100010011;
ROM[17742] <= 32'b00000111110001101010001110000011;
ROM[17743] <= 32'b11111111110000010000000100010011;
ROM[17744] <= 32'b00000000000000010010010000000011;
ROM[17745] <= 32'b00000000011101000000001110110011;
ROM[17746] <= 32'b00000000000000111000001100010011;
ROM[17747] <= 32'b00000000110100110000010000110011;
ROM[17748] <= 32'b00000000000001000010001110000011;
ROM[17749] <= 32'b00000000011100010010000000100011;
ROM[17750] <= 32'b00000000010000010000000100010011;
ROM[17751] <= 32'b00010000000000000000001110010011;
ROM[17752] <= 32'b01000000011100000000001110110011;
ROM[17753] <= 32'b11111111110000010000000100010011;
ROM[17754] <= 32'b00000000000000010010010000000011;
ROM[17755] <= 32'b00000000011101000111001110110011;
ROM[17756] <= 32'b00000010011100011010000000100011;
ROM[17757] <= 32'b00000001000000011010001110000011;
ROM[17758] <= 32'b00000000011100010010000000100011;
ROM[17759] <= 32'b00000000010000010000000100010011;
ROM[17760] <= 32'b00000111110001101010001110000011;
ROM[17761] <= 32'b11111111110000010000000100010011;
ROM[17762] <= 32'b00000000000000010010010000000011;
ROM[17763] <= 32'b00000000011101000000001110110011;
ROM[17764] <= 32'b00000000011100010010000000100011;
ROM[17765] <= 32'b00000000010000010000000100010011;
ROM[17766] <= 32'b00000010000000011010001110000011;
ROM[17767] <= 32'b00000000011101100010000000100011;
ROM[17768] <= 32'b11111111110000010000000100010011;
ROM[17769] <= 32'b00000000000000010010001110000011;
ROM[17770] <= 32'b00000000000000111000001100010011;
ROM[17771] <= 32'b00000000000001100010001110000011;
ROM[17772] <= 32'b00000000110100110000010000110011;
ROM[17773] <= 32'b00000000011101000010000000100011;
ROM[17774] <= 32'b00000000000000011010001110000011;
ROM[17775] <= 32'b00000000011100010010000000100011;
ROM[17776] <= 32'b00000000010000010000000100010011;
ROM[17777] <= 32'b00000000101000000000001110010011;
ROM[17778] <= 32'b11111111110000010000000100010011;
ROM[17779] <= 32'b00000000000000010010010000000011;
ROM[17780] <= 32'b00000000011101000000001110110011;
ROM[17781] <= 32'b00000000011100011010000000100011;
ROM[17782] <= 32'b00000000010000011010001110000011;
ROM[17783] <= 32'b00000000011100010010000000100011;
ROM[17784] <= 32'b00000000010000010000000100010011;
ROM[17785] <= 32'b00000000000100000000001110010011;
ROM[17786] <= 32'b11111111110000010000000100010011;
ROM[17787] <= 32'b00000000000000010010010000000011;
ROM[17788] <= 32'b00000000011101000000001110110011;
ROM[17789] <= 32'b00000000011100011010001000100011;
ROM[17790] <= 32'b10010011000111111111000011101111;
ROM[17791] <= 32'b00000000000000000000001110010011;
ROM[17792] <= 32'b00000000011100010010000000100011;
ROM[17793] <= 32'b00000000010000010000000100010011;
ROM[17794] <= 32'b00000001010000000000001110010011;
ROM[17795] <= 32'b01000000011100011000001110110011;
ROM[17796] <= 32'b00000000000000111010000010000011;
ROM[17797] <= 32'b11111111110000010000000100010011;
ROM[17798] <= 32'b00000000000000010010001110000011;
ROM[17799] <= 32'b00000000011100100010000000100011;
ROM[17800] <= 32'b00000000010000100000000100010011;
ROM[17801] <= 32'b00000001010000000000001110010011;
ROM[17802] <= 32'b01000000011100011000001110110011;
ROM[17803] <= 32'b00000000010000111010000110000011;
ROM[17804] <= 32'b00000000100000111010001000000011;
ROM[17805] <= 32'b00000000110000111010001010000011;
ROM[17806] <= 32'b00000001000000111010001100000011;
ROM[17807] <= 32'b00000000000000001000000011100111;
ROM[17808] <= 32'b00000000000000010010000000100011;
ROM[17809] <= 32'b00000000010000010000000100010011;
ROM[17810] <= 32'b00000000110000000000001110010011;
ROM[17811] <= 32'b00000000011100010010000000100011;
ROM[17812] <= 32'b00000000010000010000000100010011;
ROM[17813] <= 32'b00000000000000010001001110110111;
ROM[17814] <= 32'b01101010000000111000001110010011;
ROM[17815] <= 32'b00000000111000111000001110110011;
ROM[17816] <= 32'b00000000011100010010000000100011;
ROM[17817] <= 32'b00000000010000010000000100010011;
ROM[17818] <= 32'b00000000001100010010000000100011;
ROM[17819] <= 32'b00000000010000010000000100010011;
ROM[17820] <= 32'b00000000010000010010000000100011;
ROM[17821] <= 32'b00000000010000010000000100010011;
ROM[17822] <= 32'b00000000010100010010000000100011;
ROM[17823] <= 32'b00000000010000010000000100010011;
ROM[17824] <= 32'b00000000011000010010000000100011;
ROM[17825] <= 32'b00000000010000010000000100010011;
ROM[17826] <= 32'b00000001010000000000001110010011;
ROM[17827] <= 32'b00000000010000111000001110010011;
ROM[17828] <= 32'b01000000011100010000001110110011;
ROM[17829] <= 32'b00000000011100000000001000110011;
ROM[17830] <= 32'b00000000001000000000000110110011;
ROM[17831] <= 32'b11110110000111110111000011101111;
ROM[17832] <= 32'b11111111110000010000000100010011;
ROM[17833] <= 32'b00000000000000010010001110000011;
ROM[17834] <= 32'b00000000011100011010000000100011;
ROM[17835] <= 32'b00000010001000000000001110010011;
ROM[17836] <= 32'b00000000011100010010000000100011;
ROM[17837] <= 32'b00000000010000010000000100010011;
ROM[17838] <= 32'b00000000000000011010001110000011;
ROM[17839] <= 32'b00000000011100010010000000100011;
ROM[17840] <= 32'b00000000010000010000000100010011;
ROM[17841] <= 32'b00000000000000010001001110110111;
ROM[17842] <= 32'b01110001000000111000001110010011;
ROM[17843] <= 32'b00000000111000111000001110110011;
ROM[17844] <= 32'b00000000011100010010000000100011;
ROM[17845] <= 32'b00000000010000010000000100010011;
ROM[17846] <= 32'b00000000001100010010000000100011;
ROM[17847] <= 32'b00000000010000010000000100010011;
ROM[17848] <= 32'b00000000010000010010000000100011;
ROM[17849] <= 32'b00000000010000010000000100010011;
ROM[17850] <= 32'b00000000010100010010000000100011;
ROM[17851] <= 32'b00000000010000010000000100010011;
ROM[17852] <= 32'b00000000011000010010000000100011;
ROM[17853] <= 32'b00000000010000010000000100010011;
ROM[17854] <= 32'b00000001010000000000001110010011;
ROM[17855] <= 32'b00000000100000111000001110010011;
ROM[17856] <= 32'b01000000011100010000001110110011;
ROM[17857] <= 32'b00000000011100000000001000110011;
ROM[17858] <= 32'b00000000001000000000000110110011;
ROM[17859] <= 32'b10011100100111110111000011101111;
ROM[17860] <= 32'b11111111110000010000000100010011;
ROM[17861] <= 32'b00000000000000010010001110000011;
ROM[17862] <= 32'b00000000011100011010000000100011;
ROM[17863] <= 32'b00000000000000011010001110000011;
ROM[17864] <= 32'b00000000011100010010000000100011;
ROM[17865] <= 32'b00000000010000010000000100010011;
ROM[17866] <= 32'b01011000000000000000001110010011;
ROM[17867] <= 32'b11111111110000010000000100010011;
ROM[17868] <= 32'b00000000000000010010010000000011;
ROM[17869] <= 32'b00000000011101000000001110110011;
ROM[17870] <= 32'b00000000011100011010000000100011;
ROM[17871] <= 32'b00000000000000000000001110010011;
ROM[17872] <= 32'b00000000011100010010000000100011;
ROM[17873] <= 32'b00000000010000010000000100010011;
ROM[17874] <= 32'b00000000000000011010001110000011;
ROM[17875] <= 32'b11111111110000010000000100010011;
ROM[17876] <= 32'b00000000000000010010010000000011;
ROM[17877] <= 32'b01000000011101000000001110110011;
ROM[17878] <= 32'b00001000011101101010011000100011;
ROM[17879] <= 32'b00000000000000000000001110010011;
ROM[17880] <= 32'b01000000011100000000001110110011;
ROM[17881] <= 32'b00000000000100111000001110010011;
ROM[17882] <= 32'b00001000011101101010100000100011;
ROM[17883] <= 32'b00000000000000000000001110010011;
ROM[17884] <= 32'b00000000011100010010000000100011;
ROM[17885] <= 32'b00000000010000010000000100010011;
ROM[17886] <= 32'b00000001010000000000001110010011;
ROM[17887] <= 32'b01000000011100011000001110110011;
ROM[17888] <= 32'b00000000000000111010000010000011;
ROM[17889] <= 32'b11111111110000010000000100010011;
ROM[17890] <= 32'b00000000000000010010001110000011;
ROM[17891] <= 32'b00000000011100100010000000100011;
ROM[17892] <= 32'b00000000010000100000000100010011;
ROM[17893] <= 32'b00000001010000000000001110010011;
ROM[17894] <= 32'b01000000011100011000001110110011;
ROM[17895] <= 32'b00000000010000111010000110000011;
ROM[17896] <= 32'b00000000100000111010001000000011;
ROM[17897] <= 32'b00000000110000111010001010000011;
ROM[17898] <= 32'b00000001000000111010001100000011;
ROM[17899] <= 32'b00000000000000001000000011100111;
ROM[17900] <= 32'b00000000000000010010000000100011;
ROM[17901] <= 32'b00000000010000010000000100010011;
ROM[17902] <= 32'b00000000000000010010000000100011;
ROM[17903] <= 32'b00000000010000010000000100010011;
ROM[17904] <= 32'b00000000000000000000001110010011;
ROM[17905] <= 32'b00000000011100011010000000100011;
ROM[17906] <= 32'b00000000000000011010001110000011;
ROM[17907] <= 32'b00000000011100010010000000100011;
ROM[17908] <= 32'b00000000010000010000000100010011;
ROM[17909] <= 32'b00000000000000000001001110110111;
ROM[17910] <= 32'b10010110000000111000001110010011;
ROM[17911] <= 32'b11111111110000010000000100010011;
ROM[17912] <= 32'b00000000000000010010010000000011;
ROM[17913] <= 32'b00000000011101000010001110110011;
ROM[17914] <= 32'b01000000011100000000001110110011;
ROM[17915] <= 32'b00000000000100111000001110010011;
ROM[17916] <= 32'b00000000000000111000101001100011;
ROM[17917] <= 32'b00000000000000010010001110110111;
ROM[17918] <= 32'b10001011110000111000001110010011;
ROM[17919] <= 32'b00000000111000111000001110110011;
ROM[17920] <= 32'b00000000000000111000000011100111;
ROM[17921] <= 32'b00000000000000011010001110000011;
ROM[17922] <= 32'b00000000011100010010000000100011;
ROM[17923] <= 32'b00000000010000010000000100010011;
ROM[17924] <= 32'b00000000000000011010001110000011;
ROM[17925] <= 32'b11111111110000010000000100010011;
ROM[17926] <= 32'b00000000000000010010010000000011;
ROM[17927] <= 32'b00000000011101000000001110110011;
ROM[17928] <= 32'b00000000011100010010000000100011;
ROM[17929] <= 32'b00000000010000010000000100010011;
ROM[17930] <= 32'b00000000000000011010001110000011;
ROM[17931] <= 32'b11111111110000010000000100010011;
ROM[17932] <= 32'b00000000000000010010010000000011;
ROM[17933] <= 32'b00000000011101000000001110110011;
ROM[17934] <= 32'b00000000011100010010000000100011;
ROM[17935] <= 32'b00000000010000010000000100010011;
ROM[17936] <= 32'b00000000000000011010001110000011;
ROM[17937] <= 32'b11111111110000010000000100010011;
ROM[17938] <= 32'b00000000000000010010010000000011;
ROM[17939] <= 32'b00000000011101000000001110110011;
ROM[17940] <= 32'b00000000011100011010001000100011;
ROM[17941] <= 32'b00000000010000011010001110000011;
ROM[17942] <= 32'b00000000011100010010000000100011;
ROM[17943] <= 32'b00000000010000010000000100010011;
ROM[17944] <= 32'b00001000110001101010001110000011;
ROM[17945] <= 32'b11111111110000010000000100010011;
ROM[17946] <= 32'b00000000000000010010010000000011;
ROM[17947] <= 32'b00000000011101000000001110110011;
ROM[17948] <= 32'b00000000011100010010000000100011;
ROM[17949] <= 32'b00000000010000010000000100010011;
ROM[17950] <= 32'b00000000000000000000001110010011;
ROM[17951] <= 32'b00000000011101100010000000100011;
ROM[17952] <= 32'b11111111110000010000000100010011;
ROM[17953] <= 32'b00000000000000010010001110000011;
ROM[17954] <= 32'b00000000000000111000001100010011;
ROM[17955] <= 32'b00000000000001100010001110000011;
ROM[17956] <= 32'b00000000110100110000010000110011;
ROM[17957] <= 32'b00000000011101000010000000100011;
ROM[17958] <= 32'b00000000000000011010001110000011;
ROM[17959] <= 32'b00000000011100010010000000100011;
ROM[17960] <= 32'b00000000010000010000000100010011;
ROM[17961] <= 32'b00000000000100000000001110010011;
ROM[17962] <= 32'b11111111110000010000000100010011;
ROM[17963] <= 32'b00000000000000010010010000000011;
ROM[17964] <= 32'b00000000011101000000001110110011;
ROM[17965] <= 32'b00000000011100011010000000100011;
ROM[17966] <= 32'b11110001000111111111000011101111;
ROM[17967] <= 32'b00000000000000000000001110010011;
ROM[17968] <= 32'b00000000011100010010000000100011;
ROM[17969] <= 32'b00000000010000010000000100010011;
ROM[17970] <= 32'b00000001010000000000001110010011;
ROM[17971] <= 32'b01000000011100011000001110110011;
ROM[17972] <= 32'b00000000000000111010000010000011;
ROM[17973] <= 32'b11111111110000010000000100010011;
ROM[17974] <= 32'b00000000000000010010001110000011;
ROM[17975] <= 32'b00000000011100100010000000100011;
ROM[17976] <= 32'b00000000010000100000000100010011;
ROM[17977] <= 32'b00000001010000000000001110010011;
ROM[17978] <= 32'b01000000011100011000001110110011;
ROM[17979] <= 32'b00000000010000111010000110000011;
ROM[17980] <= 32'b00000000100000111010001000000011;
ROM[17981] <= 32'b00000000110000111010001010000011;
ROM[17982] <= 32'b00000001000000111010001100000011;
ROM[17983] <= 32'b00000000000000001000000011100111;
ROM[17984] <= 32'b00000000001100000000001110010011;
ROM[17985] <= 32'b00000000011100010010000000100011;
ROM[17986] <= 32'b00000000010000010000000100010011;
ROM[17987] <= 32'b00000000000000010010001110110111;
ROM[17988] <= 32'b10010101100000111000001110010011;
ROM[17989] <= 32'b00000000111000111000001110110011;
ROM[17990] <= 32'b00000000011100010010000000100011;
ROM[17991] <= 32'b00000000010000010000000100010011;
ROM[17992] <= 32'b00000000001100010010000000100011;
ROM[17993] <= 32'b00000000010000010000000100010011;
ROM[17994] <= 32'b00000000010000010010000000100011;
ROM[17995] <= 32'b00000000010000010000000100010011;
ROM[17996] <= 32'b00000000010100010010000000100011;
ROM[17997] <= 32'b00000000010000010000000100010011;
ROM[17998] <= 32'b00000000011000010010000000100011;
ROM[17999] <= 32'b00000000010000010000000100010011;
ROM[18000] <= 32'b00000001010000000000001110010011;
ROM[18001] <= 32'b00000000010000111000001110010011;
ROM[18002] <= 32'b01000000011100010000001110110011;
ROM[18003] <= 32'b00000000011100000000001000110011;
ROM[18004] <= 32'b00000000001000000000000110110011;
ROM[18005] <= 32'b10101011000111111000000011101111;
ROM[18006] <= 32'b11111111110000010000000100010011;
ROM[18007] <= 32'b00000000000000010010001110000011;
ROM[18008] <= 32'b00000000000000111000001010010011;
ROM[18009] <= 32'b00000000000000100010001110000011;
ROM[18010] <= 32'b00000000011100010010000000100011;
ROM[18011] <= 32'b00000000010000010000000100010011;
ROM[18012] <= 32'b00000000000000000000001110010011;
ROM[18013] <= 32'b11111111110000010000000100010011;
ROM[18014] <= 32'b00000000000000010010010000000011;
ROM[18015] <= 32'b00000000011101000010010010110011;
ROM[18016] <= 32'b00000000100000111010010100110011;
ROM[18017] <= 32'b00000000101001001000001110110011;
ROM[18018] <= 32'b00000000000100111000001110010011;
ROM[18019] <= 32'b00000000000100111111001110010011;
ROM[18020] <= 32'b00000000000000111000101001100011;
ROM[18021] <= 32'b00000000000000010010001110110111;
ROM[18022] <= 32'b10011010100000111000001110010011;
ROM[18023] <= 32'b00000000111000111000001110110011;
ROM[18024] <= 32'b00000000000000111000000011100111;
ROM[18025] <= 32'b00000001000000000000000011101111;
ROM[18026] <= 32'b00000000000100000000001110010011;
ROM[18027] <= 32'b00000000011100100010000000100011;
ROM[18028] <= 32'b00000000010000000000000011101111;
ROM[18029] <= 32'b00000000000000000000001110010011;
ROM[18030] <= 32'b00000000110100101000010000110011;
ROM[18031] <= 32'b00000000011101000010001000100011;
ROM[18032] <= 32'b00000000000000100010001110000011;
ROM[18033] <= 32'b00000000110100101000010000110011;
ROM[18034] <= 32'b00000000011101000010000000100011;
ROM[18035] <= 32'b00000000000000100010001110000011;
ROM[18036] <= 32'b00000000011100010010000000100011;
ROM[18037] <= 32'b00000000010000010000000100010011;
ROM[18038] <= 32'b00000000000000010010001110110111;
ROM[18039] <= 32'b10100010010000111000001110010011;
ROM[18040] <= 32'b00000000111000111000001110110011;
ROM[18041] <= 32'b00000000011100010010000000100011;
ROM[18042] <= 32'b00000000010000010000000100010011;
ROM[18043] <= 32'b00000000001100010010000000100011;
ROM[18044] <= 32'b00000000010000010000000100010011;
ROM[18045] <= 32'b00000000010000010010000000100011;
ROM[18046] <= 32'b00000000010000010000000100010011;
ROM[18047] <= 32'b00000000010100010010000000100011;
ROM[18048] <= 32'b00000000010000010000000100010011;
ROM[18049] <= 32'b00000000011000010010000000100011;
ROM[18050] <= 32'b00000000010000010000000100010011;
ROM[18051] <= 32'b00000001010000000000001110010011;
ROM[18052] <= 32'b00000000010000111000001110010011;
ROM[18053] <= 32'b01000000011100010000001110110011;
ROM[18054] <= 32'b00000000011100000000001000110011;
ROM[18055] <= 32'b00000000001000000000000110110011;
ROM[18056] <= 32'b10100010000111101110000011101111;
ROM[18057] <= 32'b11111111110000010000000100010011;
ROM[18058] <= 32'b00000000000000010010001110000011;
ROM[18059] <= 32'b00000000110100101000010000110011;
ROM[18060] <= 32'b00000000011101000010010000100011;
ROM[18061] <= 32'b00000000010100010010000000100011;
ROM[18062] <= 32'b00000000010000010000000100010011;
ROM[18063] <= 32'b00000001010000000000001110010011;
ROM[18064] <= 32'b01000000011100011000001110110011;
ROM[18065] <= 32'b00000000000000111010000010000011;
ROM[18066] <= 32'b11111111110000010000000100010011;
ROM[18067] <= 32'b00000000000000010010001110000011;
ROM[18068] <= 32'b00000000011100100010000000100011;
ROM[18069] <= 32'b00000000010000100000000100010011;
ROM[18070] <= 32'b00000001010000000000001110010011;
ROM[18071] <= 32'b01000000011100011000001110110011;
ROM[18072] <= 32'b00000000010000111010000110000011;
ROM[18073] <= 32'b00000000100000111010001000000011;
ROM[18074] <= 32'b00000000110000111010001010000011;
ROM[18075] <= 32'b00000001000000111010001100000011;
ROM[18076] <= 32'b00000000000000001000000011100111;
ROM[18077] <= 32'b00000000000000100010001110000011;
ROM[18078] <= 32'b00000000000000111000001010010011;
ROM[18079] <= 32'b00000000110100101000010000110011;
ROM[18080] <= 32'b00000000010001000010001110000011;
ROM[18081] <= 32'b00000000011100010010000000100011;
ROM[18082] <= 32'b00000000010000010000000100010011;
ROM[18083] <= 32'b00000001010000000000001110010011;
ROM[18084] <= 32'b01000000011100011000001110110011;
ROM[18085] <= 32'b00000000000000111010000010000011;
ROM[18086] <= 32'b11111111110000010000000100010011;
ROM[18087] <= 32'b00000000000000010010001110000011;
ROM[18088] <= 32'b00000000011100100010000000100011;
ROM[18089] <= 32'b00000000010000100000000100010011;
ROM[18090] <= 32'b00000001010000000000001110010011;
ROM[18091] <= 32'b01000000011100011000001110110011;
ROM[18092] <= 32'b00000000010000111010000110000011;
ROM[18093] <= 32'b00000000100000111010001000000011;
ROM[18094] <= 32'b00000000110000111010001010000011;
ROM[18095] <= 32'b00000001000000111010001100000011;
ROM[18096] <= 32'b00000000000000001000000011100111;
ROM[18097] <= 32'b00000000000000010010000000100011;
ROM[18098] <= 32'b00000000010000010000000100010011;
ROM[18099] <= 32'b00000000000000100010001110000011;
ROM[18100] <= 32'b00000000000000111000001010010011;
ROM[18101] <= 32'b00000000010000100010001110000011;
ROM[18102] <= 32'b00000000011100010010000000100011;
ROM[18103] <= 32'b00000000010000010000000100010011;
ROM[18104] <= 32'b00000000010000000000001110010011;
ROM[18105] <= 32'b00000000011100010010000000100011;
ROM[18106] <= 32'b00000000010000010000000100010011;
ROM[18107] <= 32'b00000000000000010010001110110111;
ROM[18108] <= 32'b10110011100000111000001110010011;
ROM[18109] <= 32'b00000000111000111000001110110011;
ROM[18110] <= 32'b00000000011100010010000000100011;
ROM[18111] <= 32'b00000000010000010000000100010011;
ROM[18112] <= 32'b00000000001100010010000000100011;
ROM[18113] <= 32'b00000000010000010000000100010011;
ROM[18114] <= 32'b00000000010000010010000000100011;
ROM[18115] <= 32'b00000000010000010000000100010011;
ROM[18116] <= 32'b00000000010100010010000000100011;
ROM[18117] <= 32'b00000000010000010000000100010011;
ROM[18118] <= 32'b00000000011000010010000000100011;
ROM[18119] <= 32'b00000000010000010000000100010011;
ROM[18120] <= 32'b00000001010000000000001110010011;
ROM[18121] <= 32'b00000000100000111000001110010011;
ROM[18122] <= 32'b01000000011100010000001110110011;
ROM[18123] <= 32'b00000000011100000000001000110011;
ROM[18124] <= 32'b00000000001000000000000110110011;
ROM[18125] <= 32'b11011010000011110111000011101111;
ROM[18126] <= 32'b11111111110000010000000100010011;
ROM[18127] <= 32'b00000000000000010010001110000011;
ROM[18128] <= 32'b00000000011100011010000000100011;
ROM[18129] <= 32'b00000000000000011010001110000011;
ROM[18130] <= 32'b00000000011100010010000000100011;
ROM[18131] <= 32'b00000000010000010000000100010011;
ROM[18132] <= 32'b00000000110100101000010000110011;
ROM[18133] <= 32'b00000000100001000010001110000011;
ROM[18134] <= 32'b11111111110000010000000100010011;
ROM[18135] <= 32'b00000000000000010010010000000011;
ROM[18136] <= 32'b00000000011101000000001110110011;
ROM[18137] <= 32'b00000000000000111000001100010011;
ROM[18138] <= 32'b00000000110100110000010000110011;
ROM[18139] <= 32'b00000000000001000010001110000011;
ROM[18140] <= 32'b00000000011100010010000000100011;
ROM[18141] <= 32'b00000000010000010000000100010011;
ROM[18142] <= 32'b00000001010000000000001110010011;
ROM[18143] <= 32'b01000000011100011000001110110011;
ROM[18144] <= 32'b00000000000000111010000010000011;
ROM[18145] <= 32'b11111111110000010000000100010011;
ROM[18146] <= 32'b00000000000000010010001110000011;
ROM[18147] <= 32'b00000000011100100010000000100011;
ROM[18148] <= 32'b00000000010000100000000100010011;
ROM[18149] <= 32'b00000001010000000000001110010011;
ROM[18150] <= 32'b01000000011100011000001110110011;
ROM[18151] <= 32'b00000000010000111010000110000011;
ROM[18152] <= 32'b00000000100000111010001000000011;
ROM[18153] <= 32'b00000000110000111010001010000011;
ROM[18154] <= 32'b00000001000000111010001100000011;
ROM[18155] <= 32'b00000000000000001000000011100111;
ROM[18156] <= 32'b00000000000000010010000000100011;
ROM[18157] <= 32'b00000000010000010000000100010011;
ROM[18158] <= 32'b00000000000000100010001110000011;
ROM[18159] <= 32'b00000000000000111000001010010011;
ROM[18160] <= 32'b00000000010000100010001110000011;
ROM[18161] <= 32'b00000000011100010010000000100011;
ROM[18162] <= 32'b00000000010000010000000100010011;
ROM[18163] <= 32'b00000000010000000000001110010011;
ROM[18164] <= 32'b00000000011100010010000000100011;
ROM[18165] <= 32'b00000000010000010000000100010011;
ROM[18166] <= 32'b00000000000000010010001110110111;
ROM[18167] <= 32'b11000010010000111000001110010011;
ROM[18168] <= 32'b00000000111000111000001110110011;
ROM[18169] <= 32'b00000000011100010010000000100011;
ROM[18170] <= 32'b00000000010000010000000100010011;
ROM[18171] <= 32'b00000000001100010010000000100011;
ROM[18172] <= 32'b00000000010000010000000100010011;
ROM[18173] <= 32'b00000000010000010010000000100011;
ROM[18174] <= 32'b00000000010000010000000100010011;
ROM[18175] <= 32'b00000000010100010010000000100011;
ROM[18176] <= 32'b00000000010000010000000100010011;
ROM[18177] <= 32'b00000000011000010010000000100011;
ROM[18178] <= 32'b00000000010000010000000100010011;
ROM[18179] <= 32'b00000001010000000000001110010011;
ROM[18180] <= 32'b00000000100000111000001110010011;
ROM[18181] <= 32'b01000000011100010000001110110011;
ROM[18182] <= 32'b00000000011100000000001000110011;
ROM[18183] <= 32'b00000000001000000000000110110011;
ROM[18184] <= 32'b11001011010011110111000011101111;
ROM[18185] <= 32'b11111111110000010000000100010011;
ROM[18186] <= 32'b00000000000000010010001110000011;
ROM[18187] <= 32'b00000000011100011010000000100011;
ROM[18188] <= 32'b00000000000000011010001110000011;
ROM[18189] <= 32'b00000000011100010010000000100011;
ROM[18190] <= 32'b00000000010000010000000100010011;
ROM[18191] <= 32'b00000000110100101000010000110011;
ROM[18192] <= 32'b00000000100001000010001110000011;
ROM[18193] <= 32'b11111111110000010000000100010011;
ROM[18194] <= 32'b00000000000000010010010000000011;
ROM[18195] <= 32'b00000000011101000000001110110011;
ROM[18196] <= 32'b00000000011100010010000000100011;
ROM[18197] <= 32'b00000000010000010000000100010011;
ROM[18198] <= 32'b00000000100000100010001110000011;
ROM[18199] <= 32'b00000000011101100010000000100011;
ROM[18200] <= 32'b11111111110000010000000100010011;
ROM[18201] <= 32'b00000000000000010010001110000011;
ROM[18202] <= 32'b00000000000000111000001100010011;
ROM[18203] <= 32'b00000000000001100010001110000011;
ROM[18204] <= 32'b00000000110100110000010000110011;
ROM[18205] <= 32'b00000000011101000010000000100011;
ROM[18206] <= 32'b00000000000000000000001110010011;
ROM[18207] <= 32'b00000000011100010010000000100011;
ROM[18208] <= 32'b00000000010000010000000100010011;
ROM[18209] <= 32'b00000001010000000000001110010011;
ROM[18210] <= 32'b01000000011100011000001110110011;
ROM[18211] <= 32'b00000000000000111010000010000011;
ROM[18212] <= 32'b11111111110000010000000100010011;
ROM[18213] <= 32'b00000000000000010010001110000011;
ROM[18214] <= 32'b00000000011100100010000000100011;
ROM[18215] <= 32'b00000000010000100000000100010011;
ROM[18216] <= 32'b00000001010000000000001110010011;
ROM[18217] <= 32'b01000000011100011000001110110011;
ROM[18218] <= 32'b00000000010000111010000110000011;
ROM[18219] <= 32'b00000000100000111010001000000011;
ROM[18220] <= 32'b00000000110000111010001010000011;
ROM[18221] <= 32'b00000001000000111010001100000011;
ROM[18222] <= 32'b00000000000000001000000011100111;
ROM[18223] <= 32'b00000000000000010010000000100011;
ROM[18224] <= 32'b00000000010000010000000100010011;
ROM[18225] <= 32'b00000000000000100010001110000011;
ROM[18226] <= 32'b00000000000000111000001010010011;
ROM[18227] <= 32'b00000000110100101000010000110011;
ROM[18228] <= 32'b00000000010001000010001110000011;
ROM[18229] <= 32'b00000000011100010010000000100011;
ROM[18230] <= 32'b00000000010000010000000100010011;
ROM[18231] <= 32'b00000000010000000000001110010011;
ROM[18232] <= 32'b00000000011100010010000000100011;
ROM[18233] <= 32'b00000000010000010000000100010011;
ROM[18234] <= 32'b00000000000000010010001110110111;
ROM[18235] <= 32'b11010011010000111000001110010011;
ROM[18236] <= 32'b00000000111000111000001110110011;
ROM[18237] <= 32'b00000000011100010010000000100011;
ROM[18238] <= 32'b00000000010000010000000100010011;
ROM[18239] <= 32'b00000000001100010010000000100011;
ROM[18240] <= 32'b00000000010000010000000100010011;
ROM[18241] <= 32'b00000000010000010010000000100011;
ROM[18242] <= 32'b00000000010000010000000100010011;
ROM[18243] <= 32'b00000000010100010010000000100011;
ROM[18244] <= 32'b00000000010000010000000100010011;
ROM[18245] <= 32'b00000000011000010010000000100011;
ROM[18246] <= 32'b00000000010000010000000100010011;
ROM[18247] <= 32'b00000001010000000000001110010011;
ROM[18248] <= 32'b00000000100000111000001110010011;
ROM[18249] <= 32'b01000000011100010000001110110011;
ROM[18250] <= 32'b00000000011100000000001000110011;
ROM[18251] <= 32'b00000000001000000000000110110011;
ROM[18252] <= 32'b10111010010011110111000011101111;
ROM[18253] <= 32'b11111111110000010000000100010011;
ROM[18254] <= 32'b00000000000000010010001110000011;
ROM[18255] <= 32'b00000000011100011010000000100011;
ROM[18256] <= 32'b00000000110100101000010000110011;
ROM[18257] <= 32'b00000000010001000010001110000011;
ROM[18258] <= 32'b00000000011100010010000000100011;
ROM[18259] <= 32'b00000000010000010000000100010011;
ROM[18260] <= 32'b00000000110100101000010000110011;
ROM[18261] <= 32'b00000000000001000010001110000011;
ROM[18262] <= 32'b11111111110000010000000100010011;
ROM[18263] <= 32'b00000000000000010010010000000011;
ROM[18264] <= 32'b00000000011101000010001110110011;
ROM[18265] <= 32'b00000000000000111000101001100011;
ROM[18266] <= 32'b00000000000000010010001110110111;
ROM[18267] <= 32'b11010111110000111000001110010011;
ROM[18268] <= 32'b00000000111000111000001110110011;
ROM[18269] <= 32'b00000000000000111000000011100111;
ROM[18270] <= 32'b00000111100000000000000011101111;
ROM[18271] <= 32'b00000000000000011010001110000011;
ROM[18272] <= 32'b00000000011100010010000000100011;
ROM[18273] <= 32'b00000000010000010000000100010011;
ROM[18274] <= 32'b00000000110100101000010000110011;
ROM[18275] <= 32'b00000000100001000010001110000011;
ROM[18276] <= 32'b11111111110000010000000100010011;
ROM[18277] <= 32'b00000000000000010010010000000011;
ROM[18278] <= 32'b00000000011101000000001110110011;
ROM[18279] <= 32'b00000000011100010010000000100011;
ROM[18280] <= 32'b00000000010000010000000100010011;
ROM[18281] <= 32'b00000000010000100010001110000011;
ROM[18282] <= 32'b00000000011101100010000000100011;
ROM[18283] <= 32'b11111111110000010000000100010011;
ROM[18284] <= 32'b00000000000000010010001110000011;
ROM[18285] <= 32'b00000000000000111000001100010011;
ROM[18286] <= 32'b00000000000001100010001110000011;
ROM[18287] <= 32'b00000000110100110000010000110011;
ROM[18288] <= 32'b00000000011101000010000000100011;
ROM[18289] <= 32'b00000000110100101000010000110011;
ROM[18290] <= 32'b00000000010001000010001110000011;
ROM[18291] <= 32'b00000000011100010010000000100011;
ROM[18292] <= 32'b00000000010000010000000100010011;
ROM[18293] <= 32'b00000000000100000000001110010011;
ROM[18294] <= 32'b11111111110000010000000100010011;
ROM[18295] <= 32'b00000000000000010010010000000011;
ROM[18296] <= 32'b00000000011101000000001110110011;
ROM[18297] <= 32'b00000000110100101000010000110011;
ROM[18298] <= 32'b00000000011101000010001000100011;
ROM[18299] <= 32'b00000000010000000000000011101111;
ROM[18300] <= 32'b00000000110100101000010000110011;
ROM[18301] <= 32'b00000000100001000010001110000011;
ROM[18302] <= 32'b00000000011100010010000000100011;
ROM[18303] <= 32'b00000000010000010000000100010011;
ROM[18304] <= 32'b00000001010000000000001110010011;
ROM[18305] <= 32'b01000000011100011000001110110011;
ROM[18306] <= 32'b00000000000000111010000010000011;
ROM[18307] <= 32'b11111111110000010000000100010011;
ROM[18308] <= 32'b00000000000000010010001110000011;
ROM[18309] <= 32'b00000000011100100010000000100011;
ROM[18310] <= 32'b00000000010000100000000100010011;
ROM[18311] <= 32'b00000001010000000000001110010011;
ROM[18312] <= 32'b01000000011100011000001110110011;
ROM[18313] <= 32'b00000000010000111010000110000011;
ROM[18314] <= 32'b00000000100000111010001000000011;
ROM[18315] <= 32'b00000000110000111010001010000011;
ROM[18316] <= 32'b00000001000000111010001100000011;
ROM[18317] <= 32'b00000000000000001000000011100111;
ROM[18318] <= 32'b00000000000000100010001110000011;
ROM[18319] <= 32'b00000000000000111000001010010011;
ROM[18320] <= 32'b00000000110100101000010000110011;
ROM[18321] <= 32'b00000000010001000010001110000011;
ROM[18322] <= 32'b00000000011100010010000000100011;
ROM[18323] <= 32'b00000000010000010000000100010011;
ROM[18324] <= 32'b00000000000000000000001110010011;
ROM[18325] <= 32'b11111111110000010000000100010011;
ROM[18326] <= 32'b00000000000000010010010000000011;
ROM[18327] <= 32'b00000000100000111010001110110011;
ROM[18328] <= 32'b00000000000000111000101001100011;
ROM[18329] <= 32'b00000000000000010010001110110111;
ROM[18330] <= 32'b11100111100000111000001110010011;
ROM[18331] <= 32'b00000000111000111000001110110011;
ROM[18332] <= 32'b00000000000000111000000011100111;
ROM[18333] <= 32'b00000011000000000000000011101111;
ROM[18334] <= 32'b00000000110100101000010000110011;
ROM[18335] <= 32'b00000000010001000010001110000011;
ROM[18336] <= 32'b00000000011100010010000000100011;
ROM[18337] <= 32'b00000000010000010000000100010011;
ROM[18338] <= 32'b00000000000100000000001110010011;
ROM[18339] <= 32'b11111111110000010000000100010011;
ROM[18340] <= 32'b00000000000000010010010000000011;
ROM[18341] <= 32'b01000000011101000000001110110011;
ROM[18342] <= 32'b00000000110100101000010000110011;
ROM[18343] <= 32'b00000000011101000010001000100011;
ROM[18344] <= 32'b00000000010000000000000011101111;
ROM[18345] <= 32'b00000000000000000000001110010011;
ROM[18346] <= 32'b00000000011100010010000000100011;
ROM[18347] <= 32'b00000000010000010000000100010011;
ROM[18348] <= 32'b00000001010000000000001110010011;
ROM[18349] <= 32'b01000000011100011000001110110011;
ROM[18350] <= 32'b00000000000000111010000010000011;
ROM[18351] <= 32'b11111111110000010000000100010011;
ROM[18352] <= 32'b00000000000000010010001110000011;
ROM[18353] <= 32'b00000000011100100010000000100011;
ROM[18354] <= 32'b00000000010000100000000100010011;
ROM[18355] <= 32'b00000001010000000000001110010011;
ROM[18356] <= 32'b01000000011100011000001110110011;
ROM[18357] <= 32'b00000000010000111010000110000011;
ROM[18358] <= 32'b00000000100000111010001000000011;
ROM[18359] <= 32'b00000000110000111010001010000011;
ROM[18360] <= 32'b00000001000000111010001100000011;
ROM[18361] <= 32'b00000000000000001000000011100111;
ROM[18362] <= 32'b00000000000000010010000000100011;
ROM[18363] <= 32'b00000000010000010000000100010011;
ROM[18364] <= 32'b00000000000000010010000000100011;
ROM[18365] <= 32'b00000000010000010000000100010011;
ROM[18366] <= 32'b00000000000000010010000000100011;
ROM[18367] <= 32'b00000000010000010000000100010011;
ROM[18368] <= 32'b00000000000000100010001110000011;
ROM[18369] <= 32'b00000000000000111000001010010011;
ROM[18370] <= 32'b00000000000000000000001110010011;
ROM[18371] <= 32'b00000000011100011010000000100011;
ROM[18372] <= 32'b00000000110100101000010000110011;
ROM[18373] <= 32'b00000000010001000010001110000011;
ROM[18374] <= 32'b00000000011100010010000000100011;
ROM[18375] <= 32'b00000000010000010000000100010011;
ROM[18376] <= 32'b00000000000000000000001110010011;
ROM[18377] <= 32'b11111111110000010000000100010011;
ROM[18378] <= 32'b00000000000000010010010000000011;
ROM[18379] <= 32'b00000000100000111010001110110011;
ROM[18380] <= 32'b00000000011100010010000000100011;
ROM[18381] <= 32'b00000000010000010000000100010011;
ROM[18382] <= 32'b00000000000000000000001110010011;
ROM[18383] <= 32'b00000000011100010010000000100011;
ROM[18384] <= 32'b00000000010000010000000100010011;
ROM[18385] <= 32'b00000000110100101000010000110011;
ROM[18386] <= 32'b00000000100001000010001110000011;
ROM[18387] <= 32'b11111111110000010000000100010011;
ROM[18388] <= 32'b00000000000000010010010000000011;
ROM[18389] <= 32'b00000000011101000000001110110011;
ROM[18390] <= 32'b00000000000000111000001100010011;
ROM[18391] <= 32'b00000000110100110000010000110011;
ROM[18392] <= 32'b00000000000001000010001110000011;
ROM[18393] <= 32'b00000000011100010010000000100011;
ROM[18394] <= 32'b00000000010000010000000100010011;
ROM[18395] <= 32'b00000010110100000000001110010011;
ROM[18396] <= 32'b11111111110000010000000100010011;
ROM[18397] <= 32'b00000000000000010010010000000011;
ROM[18398] <= 32'b00000000011101000010010010110011;
ROM[18399] <= 32'b00000000100000111010010100110011;
ROM[18400] <= 32'b00000000101001001000001110110011;
ROM[18401] <= 32'b00000000000100111000001110010011;
ROM[18402] <= 32'b00000000000100111111001110010011;
ROM[18403] <= 32'b11111111110000010000000100010011;
ROM[18404] <= 32'b00000000000000010010010000000011;
ROM[18405] <= 32'b00000000011101000111001110110011;
ROM[18406] <= 32'b00000000000000111000101001100011;
ROM[18407] <= 32'b00000000000000010010001110110111;
ROM[18408] <= 32'b11111011000000111000001110010011;
ROM[18409] <= 32'b00000000111000111000001110110011;
ROM[18410] <= 32'b00000000000000111000000011100111;
ROM[18411] <= 32'b00000010000000000000000011101111;
ROM[18412] <= 32'b00000000000000000000001110010011;
ROM[18413] <= 32'b01000000011100000000001110110011;
ROM[18414] <= 32'b00000000000100111000001110010011;
ROM[18415] <= 32'b00000000011100011010010000100011;
ROM[18416] <= 32'b00000000000100000000001110010011;
ROM[18417] <= 32'b00000000011100011010001000100011;
ROM[18418] <= 32'b00000001010000000000000011101111;
ROM[18419] <= 32'b00000000000000000000001110010011;
ROM[18420] <= 32'b00000000011100011010010000100011;
ROM[18421] <= 32'b00000000000000000000001110010011;
ROM[18422] <= 32'b00000000011100011010001000100011;
ROM[18423] <= 32'b00000000010000011010001110000011;
ROM[18424] <= 32'b00000000011100010010000000100011;
ROM[18425] <= 32'b00000000010000010000000100010011;
ROM[18426] <= 32'b00000000110100101000010000110011;
ROM[18427] <= 32'b00000000010001000010001110000011;
ROM[18428] <= 32'b11111111110000010000000100010011;
ROM[18429] <= 32'b00000000000000010010010000000011;
ROM[18430] <= 32'b00000000011101000010001110110011;
ROM[18431] <= 32'b00000000011100010010000000100011;
ROM[18432] <= 32'b00000000010000010000000100010011;
ROM[18433] <= 32'b00000000010000000000001110010011;
ROM[18434] <= 32'b00000000011100010010000000100011;
ROM[18435] <= 32'b00000000010000010000000100010011;
ROM[18436] <= 32'b00000000010000011010001110000011;
ROM[18437] <= 32'b00000000011100010010000000100011;
ROM[18438] <= 32'b00000000010000010000000100010011;
ROM[18439] <= 32'b00000000000000010010001110110111;
ROM[18440] <= 32'b00000110100000111000001110010011;
ROM[18441] <= 32'b00000000111000111000001110110011;
ROM[18442] <= 32'b00000000011100010010000000100011;
ROM[18443] <= 32'b00000000010000010000000100010011;
ROM[18444] <= 32'b00000000001100010010000000100011;
ROM[18445] <= 32'b00000000010000010000000100010011;
ROM[18446] <= 32'b00000000010000010010000000100011;
ROM[18447] <= 32'b00000000010000010000000100010011;
ROM[18448] <= 32'b00000000010100010010000000100011;
ROM[18449] <= 32'b00000000010000010000000100010011;
ROM[18450] <= 32'b00000000011000010010000000100011;
ROM[18451] <= 32'b00000000010000010000000100010011;
ROM[18452] <= 32'b00000001010000000000001110010011;
ROM[18453] <= 32'b00000000100000111000001110010011;
ROM[18454] <= 32'b01000000011100010000001110110011;
ROM[18455] <= 32'b00000000011100000000001000110011;
ROM[18456] <= 32'b00000000001000000000000110110011;
ROM[18457] <= 32'b10000111000011110111000011101111;
ROM[18458] <= 32'b00000000110100101000010000110011;
ROM[18459] <= 32'b00000000100001000010001110000011;
ROM[18460] <= 32'b11111111110000010000000100010011;
ROM[18461] <= 32'b00000000000000010010010000000011;
ROM[18462] <= 32'b00000000011101000000001110110011;
ROM[18463] <= 32'b00000000000000111000001100010011;
ROM[18464] <= 32'b00000000110100110000010000110011;
ROM[18465] <= 32'b00000000000001000010001110000011;
ROM[18466] <= 32'b00000000011100010010000000100011;
ROM[18467] <= 32'b00000000010000010000000100010011;
ROM[18468] <= 32'b00000000000000010010001110110111;
ROM[18469] <= 32'b00001101110000111000001110010011;
ROM[18470] <= 32'b00000000111000111000001110110011;
ROM[18471] <= 32'b00000000011100010010000000100011;
ROM[18472] <= 32'b00000000010000010000000100010011;
ROM[18473] <= 32'b00000000001100010010000000100011;
ROM[18474] <= 32'b00000000010000010000000100010011;
ROM[18475] <= 32'b00000000010000010010000000100011;
ROM[18476] <= 32'b00000000010000010000000100010011;
ROM[18477] <= 32'b00000000010100010010000000100011;
ROM[18478] <= 32'b00000000010000010000000100010011;
ROM[18479] <= 32'b00000000011000010010000000100011;
ROM[18480] <= 32'b00000000010000010000000100010011;
ROM[18481] <= 32'b00000001010000000000001110010011;
ROM[18482] <= 32'b00000000010000111000001110010011;
ROM[18483] <= 32'b01000000011100010000001110110011;
ROM[18484] <= 32'b00000000011100000000001000110011;
ROM[18485] <= 32'b00000000001000000000000110110011;
ROM[18486] <= 32'b00100101100000000000000011101111;
ROM[18487] <= 32'b11111111110000010000000100010011;
ROM[18488] <= 32'b00000000000000010010001110000011;
ROM[18489] <= 32'b11111111110000010000000100010011;
ROM[18490] <= 32'b00000000000000010010010000000011;
ROM[18491] <= 32'b00000000011101000111001110110011;
ROM[18492] <= 32'b01000000011100000000001110110011;
ROM[18493] <= 32'b00000000000100111000001110010011;
ROM[18494] <= 32'b00000000000000111000101001100011;
ROM[18495] <= 32'b00000000000000010010001110110111;
ROM[18496] <= 32'b00101000010000111000001110010011;
ROM[18497] <= 32'b00000000111000111000001110110011;
ROM[18498] <= 32'b00000000000000111000000011100111;
ROM[18499] <= 32'b00000000000000011010001110000011;
ROM[18500] <= 32'b00000000011100010010000000100011;
ROM[18501] <= 32'b00000000010000010000000100010011;
ROM[18502] <= 32'b00000000101000000000001110010011;
ROM[18503] <= 32'b00000000011100010010000000100011;
ROM[18504] <= 32'b00000000010000010000000100010011;
ROM[18505] <= 32'b00000000000000010010001110110111;
ROM[18506] <= 32'b00010111000000111000001110010011;
ROM[18507] <= 32'b00000000111000111000001110110011;
ROM[18508] <= 32'b00000000011100010010000000100011;
ROM[18509] <= 32'b00000000010000010000000100010011;
ROM[18510] <= 32'b00000000001100010010000000100011;
ROM[18511] <= 32'b00000000010000010000000100010011;
ROM[18512] <= 32'b00000000010000010010000000100011;
ROM[18513] <= 32'b00000000010000010000000100010011;
ROM[18514] <= 32'b00000000010100010010000000100011;
ROM[18515] <= 32'b00000000010000010000000100010011;
ROM[18516] <= 32'b00000000011000010010000000100011;
ROM[18517] <= 32'b00000000010000010000000100010011;
ROM[18518] <= 32'b00000001010000000000001110010011;
ROM[18519] <= 32'b00000000100000111000001110010011;
ROM[18520] <= 32'b01000000011100010000001110110011;
ROM[18521] <= 32'b00000000011100000000001000110011;
ROM[18522] <= 32'b00000000001000000000000110110011;
ROM[18523] <= 32'b11110110100111110110000011101111;
ROM[18524] <= 32'b00000000010000000000001110010011;
ROM[18525] <= 32'b00000000011100010010000000100011;
ROM[18526] <= 32'b00000000010000010000000100010011;
ROM[18527] <= 32'b00000000010000011010001110000011;
ROM[18528] <= 32'b00000000011100010010000000100011;
ROM[18529] <= 32'b00000000010000010000000100010011;
ROM[18530] <= 32'b00000000000000010010001110110111;
ROM[18531] <= 32'b00011101010000111000001110010011;
ROM[18532] <= 32'b00000000111000111000001110110011;
ROM[18533] <= 32'b00000000011100010010000000100011;
ROM[18534] <= 32'b00000000010000010000000100010011;
ROM[18535] <= 32'b00000000001100010010000000100011;
ROM[18536] <= 32'b00000000010000010000000100010011;
ROM[18537] <= 32'b00000000010000010010000000100011;
ROM[18538] <= 32'b00000000010000010000000100010011;
ROM[18539] <= 32'b00000000010100010010000000100011;
ROM[18540] <= 32'b00000000010000010000000100010011;
ROM[18541] <= 32'b00000000011000010010000000100011;
ROM[18542] <= 32'b00000000010000010000000100010011;
ROM[18543] <= 32'b00000001010000000000001110010011;
ROM[18544] <= 32'b00000000100000111000001110010011;
ROM[18545] <= 32'b01000000011100010000001110110011;
ROM[18546] <= 32'b00000000011100000000001000110011;
ROM[18547] <= 32'b00000000001000000000000110110011;
ROM[18548] <= 32'b11110000010111110110000011101111;
ROM[18549] <= 32'b00000000110100101000010000110011;
ROM[18550] <= 32'b00000000100001000010001110000011;
ROM[18551] <= 32'b11111111110000010000000100010011;
ROM[18552] <= 32'b00000000000000010010010000000011;
ROM[18553] <= 32'b00000000011101000000001110110011;
ROM[18554] <= 32'b00000000000000111000001100010011;
ROM[18555] <= 32'b00000000110100110000010000110011;
ROM[18556] <= 32'b00000000000001000010001110000011;
ROM[18557] <= 32'b00000000011100010010000000100011;
ROM[18558] <= 32'b00000000010000010000000100010011;
ROM[18559] <= 32'b00000000000000010010001110110111;
ROM[18560] <= 32'b00100100100000111000001110010011;
ROM[18561] <= 32'b00000000111000111000001110110011;
ROM[18562] <= 32'b00000000011100010010000000100011;
ROM[18563] <= 32'b00000000010000010000000100010011;
ROM[18564] <= 32'b00000000001100010010000000100011;
ROM[18565] <= 32'b00000000010000010000000100010011;
ROM[18566] <= 32'b00000000010000010010000000100011;
ROM[18567] <= 32'b00000000010000010000000100010011;
ROM[18568] <= 32'b00000000010100010010000000100011;
ROM[18569] <= 32'b00000000010000010000000100010011;
ROM[18570] <= 32'b00000000011000010010000000100011;
ROM[18571] <= 32'b00000000010000010000000100010011;
ROM[18572] <= 32'b00000001010000000000001110010011;
ROM[18573] <= 32'b00000000010000111000001110010011;
ROM[18574] <= 32'b01000000011100010000001110110011;
ROM[18575] <= 32'b00000000011100000000001000110011;
ROM[18576] <= 32'b00000000001000000000000110110011;
ROM[18577] <= 32'b00011000100000000000000011101111;
ROM[18578] <= 32'b11111111110000010000000100010011;
ROM[18579] <= 32'b00000000000000010010001110000011;
ROM[18580] <= 32'b11111111110000010000000100010011;
ROM[18581] <= 32'b00000000000000010010010000000011;
ROM[18582] <= 32'b00000000011101000000001110110011;
ROM[18583] <= 32'b00000000011100011010000000100011;
ROM[18584] <= 32'b00000000010000011010001110000011;
ROM[18585] <= 32'b00000000011100010010000000100011;
ROM[18586] <= 32'b00000000010000010000000100010011;
ROM[18587] <= 32'b00000000000100000000001110010011;
ROM[18588] <= 32'b11111111110000010000000100010011;
ROM[18589] <= 32'b00000000000000010010010000000011;
ROM[18590] <= 32'b00000000011101000000001110110011;
ROM[18591] <= 32'b00000000011100011010001000100011;
ROM[18592] <= 32'b11010101110111111111000011101111;
ROM[18593] <= 32'b00000000100000011010001110000011;
ROM[18594] <= 32'b00000000000000111000101001100011;
ROM[18595] <= 32'b00000000000000010010001110110111;
ROM[18596] <= 32'b00101010000000111000001110010011;
ROM[18597] <= 32'b00000000111000111000001110110011;
ROM[18598] <= 32'b00000000000000111000000011100111;
ROM[18599] <= 32'b00000101000000000000000011101111;
ROM[18600] <= 32'b00000000000000011010001110000011;
ROM[18601] <= 32'b01000000011100000000001110110011;
ROM[18602] <= 32'b00000000011100010010000000100011;
ROM[18603] <= 32'b00000000010000010000000100010011;
ROM[18604] <= 32'b00000001010000000000001110010011;
ROM[18605] <= 32'b01000000011100011000001110110011;
ROM[18606] <= 32'b00000000000000111010000010000011;
ROM[18607] <= 32'b11111111110000010000000100010011;
ROM[18608] <= 32'b00000000000000010010001110000011;
ROM[18609] <= 32'b00000000011100100010000000100011;
ROM[18610] <= 32'b00000000010000100000000100010011;
ROM[18611] <= 32'b00000001010000000000001110010011;
ROM[18612] <= 32'b01000000011100011000001110110011;
ROM[18613] <= 32'b00000000010000111010000110000011;
ROM[18614] <= 32'b00000000100000111010001000000011;
ROM[18615] <= 32'b00000000110000111010001010000011;
ROM[18616] <= 32'b00000001000000111010001100000011;
ROM[18617] <= 32'b00000000000000001000000011100111;
ROM[18618] <= 32'b00000100100000000000000011101111;
ROM[18619] <= 32'b00000000000000011010001110000011;
ROM[18620] <= 32'b00000000011100010010000000100011;
ROM[18621] <= 32'b00000000010000010000000100010011;
ROM[18622] <= 32'b00000001010000000000001110010011;
ROM[18623] <= 32'b01000000011100011000001110110011;
ROM[18624] <= 32'b00000000000000111010000010000011;
ROM[18625] <= 32'b11111111110000010000000100010011;
ROM[18626] <= 32'b00000000000000010010001110000011;
ROM[18627] <= 32'b00000000011100100010000000100011;
ROM[18628] <= 32'b00000000010000100000000100010011;
ROM[18629] <= 32'b00000001010000000000001110010011;
ROM[18630] <= 32'b01000000011100011000001110110011;
ROM[18631] <= 32'b00000000010000111010000110000011;
ROM[18632] <= 32'b00000000100000111010001000000011;
ROM[18633] <= 32'b00000000110000111010001010000011;
ROM[18634] <= 32'b00000001000000111010001100000011;
ROM[18635] <= 32'b00000000000000001000000011100111;
ROM[18636] <= 32'b00000000000000100010001110000011;
ROM[18637] <= 32'b00000000011100010010000000100011;
ROM[18638] <= 32'b00000000010000010000000100010011;
ROM[18639] <= 32'b00000011000000000000001110010011;
ROM[18640] <= 32'b11111111110000010000000100010011;
ROM[18641] <= 32'b00000000000000010010010000000011;
ROM[18642] <= 32'b00000000011101000010001110110011;
ROM[18643] <= 32'b01000000011100000000001110110011;
ROM[18644] <= 32'b00000000000100111000001110010011;
ROM[18645] <= 32'b00000000011100010010000000100011;
ROM[18646] <= 32'b00000000010000010000000100010011;
ROM[18647] <= 32'b00000000000000100010001110000011;
ROM[18648] <= 32'b00000000011100010010000000100011;
ROM[18649] <= 32'b00000000010000010000000100010011;
ROM[18650] <= 32'b00000011100100000000001110010011;
ROM[18651] <= 32'b11111111110000010000000100010011;
ROM[18652] <= 32'b00000000000000010010010000000011;
ROM[18653] <= 32'b00000000100000111010001110110011;
ROM[18654] <= 32'b01000000011100000000001110110011;
ROM[18655] <= 32'b00000000000100111000001110010011;
ROM[18656] <= 32'b11111111110000010000000100010011;
ROM[18657] <= 32'b00000000000000010010010000000011;
ROM[18658] <= 32'b00000000011101000111001110110011;
ROM[18659] <= 32'b00000000011100010010000000100011;
ROM[18660] <= 32'b00000000010000010000000100010011;
ROM[18661] <= 32'b00000001010000000000001110010011;
ROM[18662] <= 32'b01000000011100011000001110110011;
ROM[18663] <= 32'b00000000000000111010000010000011;
ROM[18664] <= 32'b11111111110000010000000100010011;
ROM[18665] <= 32'b00000000000000010010001110000011;
ROM[18666] <= 32'b00000000011100100010000000100011;
ROM[18667] <= 32'b00000000010000100000000100010011;
ROM[18668] <= 32'b00000001010000000000001110010011;
ROM[18669] <= 32'b01000000011100011000001110110011;
ROM[18670] <= 32'b00000000010000111010000110000011;
ROM[18671] <= 32'b00000000100000111010001000000011;
ROM[18672] <= 32'b00000000110000111010001010000011;
ROM[18673] <= 32'b00000001000000111010001100000011;
ROM[18674] <= 32'b00000000000000001000000011100111;
ROM[18675] <= 32'b00000000000000100010001110000011;
ROM[18676] <= 32'b00000000011100010010000000100011;
ROM[18677] <= 32'b00000000010000010000000100010011;
ROM[18678] <= 32'b00000011000000000000001110010011;
ROM[18679] <= 32'b11111111110000010000000100010011;
ROM[18680] <= 32'b00000000000000010010010000000011;
ROM[18681] <= 32'b01000000011101000000001110110011;
ROM[18682] <= 32'b00000000011100010010000000100011;
ROM[18683] <= 32'b00000000010000010000000100010011;
ROM[18684] <= 32'b00000001010000000000001110010011;
ROM[18685] <= 32'b01000000011100011000001110110011;
ROM[18686] <= 32'b00000000000000111010000010000011;
ROM[18687] <= 32'b11111111110000010000000100010011;
ROM[18688] <= 32'b00000000000000010010001110000011;
ROM[18689] <= 32'b00000000011100100010000000100011;
ROM[18690] <= 32'b00000000010000100000000100010011;
ROM[18691] <= 32'b00000001010000000000001110010011;
ROM[18692] <= 32'b01000000011100011000001110110011;
ROM[18693] <= 32'b00000000010000111010000110000011;
ROM[18694] <= 32'b00000000100000111010001000000011;
ROM[18695] <= 32'b00000000110000111010001010000011;
ROM[18696] <= 32'b00000001000000111010001100000011;
ROM[18697] <= 32'b00000000000000001000000011100111;
ROM[18698] <= 32'b00000000000000100010001110000011;
ROM[18699] <= 32'b00000000011100010010000000100011;
ROM[18700] <= 32'b00000000010000010000000100010011;
ROM[18701] <= 32'b00000011000000000000001110010011;
ROM[18702] <= 32'b11111111110000010000000100010011;
ROM[18703] <= 32'b00000000000000010010010000000011;
ROM[18704] <= 32'b00000000011101000000001110110011;
ROM[18705] <= 32'b00000000011100010010000000100011;
ROM[18706] <= 32'b00000000010000010000000100010011;
ROM[18707] <= 32'b00000001010000000000001110010011;
ROM[18708] <= 32'b01000000011100011000001110110011;
ROM[18709] <= 32'b00000000000000111010000010000011;
ROM[18710] <= 32'b11111111110000010000000100010011;
ROM[18711] <= 32'b00000000000000010010001110000011;
ROM[18712] <= 32'b00000000011100100010000000100011;
ROM[18713] <= 32'b00000000010000100000000100010011;
ROM[18714] <= 32'b00000001010000000000001110010011;
ROM[18715] <= 32'b01000000011100011000001110110011;
ROM[18716] <= 32'b00000000010000111010000110000011;
ROM[18717] <= 32'b00000000100000111010001000000011;
ROM[18718] <= 32'b00000000110000111010001010000011;
ROM[18719] <= 32'b00000001000000111010001100000011;
ROM[18720] <= 32'b00000000000000001000000011100111;
ROM[18721] <= 32'b00000000000000100010001110000011;
ROM[18722] <= 32'b00000000000000111000001010010011;
ROM[18723] <= 32'b00000000000000000000001110010011;
ROM[18724] <= 32'b00000000110100101000010000110011;
ROM[18725] <= 32'b00000000011101000010001000100011;
ROM[18726] <= 32'b00000000000000000000001110010011;
ROM[18727] <= 32'b00000000011100010010000000100011;
ROM[18728] <= 32'b00000000010000010000000100010011;
ROM[18729] <= 32'b00000001010000000000001110010011;
ROM[18730] <= 32'b01000000011100011000001110110011;
ROM[18731] <= 32'b00000000000000111010000010000011;
ROM[18732] <= 32'b11111111110000010000000100010011;
ROM[18733] <= 32'b00000000000000010010001110000011;
ROM[18734] <= 32'b00000000011100100010000000100011;
ROM[18735] <= 32'b00000000010000100000000100010011;
ROM[18736] <= 32'b00000001010000000000001110010011;
ROM[18737] <= 32'b01000000011100011000001110110011;
ROM[18738] <= 32'b00000000010000111010000110000011;
ROM[18739] <= 32'b00000000100000111010001000000011;
ROM[18740] <= 32'b00000000110000111010001010000011;
ROM[18741] <= 32'b00000001000000111010001100000011;
ROM[18742] <= 32'b00000000000000001000000011100111;
ROM[18743] <= 32'b00000000000000100010001110000011;
ROM[18744] <= 32'b00000000000000111000001010010011;
ROM[18745] <= 32'b00000000010100010010000000100011;
ROM[18746] <= 32'b00000000010000010000000100010011;
ROM[18747] <= 32'b00000000000000010010001110110111;
ROM[18748] <= 32'b01010011100000111000001110010011;
ROM[18749] <= 32'b00000000111000111000001110110011;
ROM[18750] <= 32'b00000000011100010010000000100011;
ROM[18751] <= 32'b00000000010000010000000100010011;
ROM[18752] <= 32'b00000000001100010010000000100011;
ROM[18753] <= 32'b00000000010000010000000100010011;
ROM[18754] <= 32'b00000000010000010010000000100011;
ROM[18755] <= 32'b00000000010000010000000100010011;
ROM[18756] <= 32'b00000000010100010010000000100011;
ROM[18757] <= 32'b00000000010000010000000100010011;
ROM[18758] <= 32'b00000000011000010010000000100011;
ROM[18759] <= 32'b00000000010000010000000100010011;
ROM[18760] <= 32'b00000001010000000000001110010011;
ROM[18761] <= 32'b00000000010000111000001110010011;
ROM[18762] <= 32'b01000000011100010000001110110011;
ROM[18763] <= 32'b00000000011100000000001000110011;
ROM[18764] <= 32'b00000000001000000000000110110011;
ROM[18765] <= 32'b11110101000111111111000011101111;
ROM[18766] <= 32'b11111111110000010000000100010011;
ROM[18767] <= 32'b00000000000000010010001110000011;
ROM[18768] <= 32'b00000000011101100010000000100011;
ROM[18769] <= 32'b00000000000000000000001110010011;
ROM[18770] <= 32'b00000000110100101000010000110011;
ROM[18771] <= 32'b00000000011101000010001000100011;
ROM[18772] <= 32'b00000000010000100010001110000011;
ROM[18773] <= 32'b00000000011100010010000000100011;
ROM[18774] <= 32'b00000000010000010000000100010011;
ROM[18775] <= 32'b00000000000000000000001110010011;
ROM[18776] <= 32'b11111111110000010000000100010011;
ROM[18777] <= 32'b00000000000000010010010000000011;
ROM[18778] <= 32'b00000000011101000010001110110011;
ROM[18779] <= 32'b00000000000000111000101001100011;
ROM[18780] <= 32'b00000000000000010010001110110111;
ROM[18781] <= 32'b01011000010000111000001110010011;
ROM[18782] <= 32'b00000000111000111000001110110011;
ROM[18783] <= 32'b00000000000000111000000011100111;
ROM[18784] <= 32'b00001000000000000000000011101111;
ROM[18785] <= 32'b00000000010000100010001110000011;
ROM[18786] <= 32'b01000000011100000000001110110011;
ROM[18787] <= 32'b00000000011100100010001000100011;
ROM[18788] <= 32'b00000000010100010010000000100011;
ROM[18789] <= 32'b00000000010000010000000100010011;
ROM[18790] <= 32'b00000010110100000000001110010011;
ROM[18791] <= 32'b00000000011100010010000000100011;
ROM[18792] <= 32'b00000000010000010000000100010011;
ROM[18793] <= 32'b00000000000000010010001110110111;
ROM[18794] <= 32'b01011111000000111000001110010011;
ROM[18795] <= 32'b00000000111000111000001110110011;
ROM[18796] <= 32'b00000000011100010010000000100011;
ROM[18797] <= 32'b00000000010000010000000100010011;
ROM[18798] <= 32'b00000000001100010010000000100011;
ROM[18799] <= 32'b00000000010000010000000100010011;
ROM[18800] <= 32'b00000000010000010010000000100011;
ROM[18801] <= 32'b00000000010000010000000100010011;
ROM[18802] <= 32'b00000000010100010010000000100011;
ROM[18803] <= 32'b00000000010000010000000100010011;
ROM[18804] <= 32'b00000000011000010010000000100011;
ROM[18805] <= 32'b00000000010000010000000100010011;
ROM[18806] <= 32'b00000001010000000000001110010011;
ROM[18807] <= 32'b00000000100000111000001110010011;
ROM[18808] <= 32'b01000000011100010000001110110011;
ROM[18809] <= 32'b00000000011100000000001000110011;
ROM[18810] <= 32'b00000000001000000000000110110011;
ROM[18811] <= 32'b11101101000011111111000011101111;
ROM[18812] <= 32'b11111111110000010000000100010011;
ROM[18813] <= 32'b00000000000000010010001110000011;
ROM[18814] <= 32'b00000000011101100010000000100011;
ROM[18815] <= 32'b00000000010000000000000011101111;
ROM[18816] <= 32'b00000000010100010010000000100011;
ROM[18817] <= 32'b00000000010000010000000100010011;
ROM[18818] <= 32'b00000000010000100010001110000011;
ROM[18819] <= 32'b00000000011100010010000000100011;
ROM[18820] <= 32'b00000000010000010000000100010011;
ROM[18821] <= 32'b00000000000000010010001110110111;
ROM[18822] <= 32'b01100110000000111000001110010011;
ROM[18823] <= 32'b00000000111000111000001110110011;
ROM[18824] <= 32'b00000000011100010010000000100011;
ROM[18825] <= 32'b00000000010000010000000100010011;
ROM[18826] <= 32'b00000000001100010010000000100011;
ROM[18827] <= 32'b00000000010000010000000100010011;
ROM[18828] <= 32'b00000000010000010010000000100011;
ROM[18829] <= 32'b00000000010000010000000100010011;
ROM[18830] <= 32'b00000000010100010010000000100011;
ROM[18831] <= 32'b00000000010000010000000100010011;
ROM[18832] <= 32'b00000000011000010010000000100011;
ROM[18833] <= 32'b00000000010000010000000100010011;
ROM[18834] <= 32'b00000001010000000000001110010011;
ROM[18835] <= 32'b00000000100000111000001110010011;
ROM[18836] <= 32'b01000000011100010000001110110011;
ROM[18837] <= 32'b00000000011100000000001000110011;
ROM[18838] <= 32'b00000000001000000000000110110011;
ROM[18839] <= 32'b00000101010000000000000011101111;
ROM[18840] <= 32'b11111111110000010000000100010011;
ROM[18841] <= 32'b00000000000000010010001110000011;
ROM[18842] <= 32'b00000000011101100010000000100011;
ROM[18843] <= 32'b00000000000000000000001110010011;
ROM[18844] <= 32'b00000000011100010010000000100011;
ROM[18845] <= 32'b00000000010000010000000100010011;
ROM[18846] <= 32'b00000001010000000000001110010011;
ROM[18847] <= 32'b01000000011100011000001110110011;
ROM[18848] <= 32'b00000000000000111010000010000011;
ROM[18849] <= 32'b11111111110000010000000100010011;
ROM[18850] <= 32'b00000000000000010010001110000011;
ROM[18851] <= 32'b00000000011100100010000000100011;
ROM[18852] <= 32'b00000000010000100000000100010011;
ROM[18853] <= 32'b00000001010000000000001110010011;
ROM[18854] <= 32'b01000000011100011000001110110011;
ROM[18855] <= 32'b00000000010000111010000110000011;
ROM[18856] <= 32'b00000000100000111010001000000011;
ROM[18857] <= 32'b00000000110000111010001010000011;
ROM[18858] <= 32'b00000001000000111010001100000011;
ROM[18859] <= 32'b00000000000000001000000011100111;
ROM[18860] <= 32'b00000000000000010010000000100011;
ROM[18861] <= 32'b00000000010000010000000100010011;
ROM[18862] <= 32'b00000000000000100010001110000011;
ROM[18863] <= 32'b00000000000000111000001010010011;
ROM[18864] <= 32'b00000000010000100010001110000011;
ROM[18865] <= 32'b00000000011100010010000000100011;
ROM[18866] <= 32'b00000000010000010000000100010011;
ROM[18867] <= 32'b00000000101000000000001110010011;
ROM[18868] <= 32'b11111111110000010000000100010011;
ROM[18869] <= 32'b00000000000000010010010000000011;
ROM[18870] <= 32'b00000000011101000010001110110011;
ROM[18871] <= 32'b00000000000000111000101001100011;
ROM[18872] <= 32'b00000000000000010010001110110111;
ROM[18873] <= 32'b01101111010000111000001110010011;
ROM[18874] <= 32'b00000000111000111000001110110011;
ROM[18875] <= 32'b00000000000000111000000011100111;
ROM[18876] <= 32'b00001100000000000000000011101111;
ROM[18877] <= 32'b00000000010100010010000000100011;
ROM[18878] <= 32'b00000000010000010000000100010011;
ROM[18879] <= 32'b00000000010000100010001110000011;
ROM[18880] <= 32'b00000000011100010010000000100011;
ROM[18881] <= 32'b00000000010000010000000100010011;
ROM[18882] <= 32'b00000000000000010010001110110111;
ROM[18883] <= 32'b01110101010000111000001110010011;
ROM[18884] <= 32'b00000000111000111000001110110011;
ROM[18885] <= 32'b00000000011100010010000000100011;
ROM[18886] <= 32'b00000000010000010000000100010011;
ROM[18887] <= 32'b00000000001100010010000000100011;
ROM[18888] <= 32'b00000000010000010000000100010011;
ROM[18889] <= 32'b00000000010000010010000000100011;
ROM[18890] <= 32'b00000000010000010000000100010011;
ROM[18891] <= 32'b00000000010100010010000000100011;
ROM[18892] <= 32'b00000000010000010000000100010011;
ROM[18893] <= 32'b00000000011000010010000000100011;
ROM[18894] <= 32'b00000000010000010000000100010011;
ROM[18895] <= 32'b00000001010000000000001110010011;
ROM[18896] <= 32'b00000000010000111000001110010011;
ROM[18897] <= 32'b01000000011100010000001110110011;
ROM[18898] <= 32'b00000000011100000000001000110011;
ROM[18899] <= 32'b00000000001000000000000110110011;
ROM[18900] <= 32'b11001101100111111111000011101111;
ROM[18901] <= 32'b00000000000000010010001110110111;
ROM[18902] <= 32'b01111010000000111000001110010011;
ROM[18903] <= 32'b00000000111000111000001110110011;
ROM[18904] <= 32'b00000000011100010010000000100011;
ROM[18905] <= 32'b00000000010000010000000100010011;
ROM[18906] <= 32'b00000000001100010010000000100011;
ROM[18907] <= 32'b00000000010000010000000100010011;
ROM[18908] <= 32'b00000000010000010010000000100011;
ROM[18909] <= 32'b00000000010000010000000100010011;
ROM[18910] <= 32'b00000000010100010010000000100011;
ROM[18911] <= 32'b00000000010000010000000100010011;
ROM[18912] <= 32'b00000000011000010010000000100011;
ROM[18913] <= 32'b00000000010000010000000100010011;
ROM[18914] <= 32'b00000001010000000000001110010011;
ROM[18915] <= 32'b00000000100000111000001110010011;
ROM[18916] <= 32'b01000000011100010000001110110011;
ROM[18917] <= 32'b00000000011100000000001000110011;
ROM[18918] <= 32'b00000000001000000000000110110011;
ROM[18919] <= 32'b11010010000011111111000011101111;
ROM[18920] <= 32'b11111111110000010000000100010011;
ROM[18921] <= 32'b00000000000000010010001110000011;
ROM[18922] <= 32'b00000000011101100010000000100011;
ROM[18923] <= 32'b00100001100000000000000011101111;
ROM[18924] <= 32'b00000000010000100010001110000011;
ROM[18925] <= 32'b00000000011100010010000000100011;
ROM[18926] <= 32'b00000000010000010000000100010011;
ROM[18927] <= 32'b00000000101000000000001110010011;
ROM[18928] <= 32'b00000000011100010010000000100011;
ROM[18929] <= 32'b00000000010000010000000100010011;
ROM[18930] <= 32'b00000000000000010011001110110111;
ROM[18931] <= 32'b10000001010000111000001110010011;
ROM[18932] <= 32'b00000000111000111000001110110011;
ROM[18933] <= 32'b00000000011100010010000000100011;
ROM[18934] <= 32'b00000000010000010000000100010011;
ROM[18935] <= 32'b00000000001100010010000000100011;
ROM[18936] <= 32'b00000000010000010000000100010011;
ROM[18937] <= 32'b00000000010000010010000000100011;
ROM[18938] <= 32'b00000000010000010000000100010011;
ROM[18939] <= 32'b00000000010100010010000000100011;
ROM[18940] <= 32'b00000000010000010000000100010011;
ROM[18941] <= 32'b00000000011000010010000000100011;
ROM[18942] <= 32'b00000000010000010000000100010011;
ROM[18943] <= 32'b00000001010000000000001110010011;
ROM[18944] <= 32'b00000000100000111000001110010011;
ROM[18945] <= 32'b01000000011100010000001110110011;
ROM[18946] <= 32'b00000000011100000000001000110011;
ROM[18947] <= 32'b00000000001000000000000110110011;
ROM[18948] <= 32'b10101110100111110110000011101111;
ROM[18949] <= 32'b11111111110000010000000100010011;
ROM[18950] <= 32'b00000000000000010010001110000011;
ROM[18951] <= 32'b00000000011100011010000000100011;
ROM[18952] <= 32'b00000000010100010010000000100011;
ROM[18953] <= 32'b00000000010000010000000100010011;
ROM[18954] <= 32'b00000000000000011010001110000011;
ROM[18955] <= 32'b00000000011100010010000000100011;
ROM[18956] <= 32'b00000000010000010000000100010011;
ROM[18957] <= 32'b00000000000000010011001110110111;
ROM[18958] <= 32'b10001000000000111000001110010011;
ROM[18959] <= 32'b00000000111000111000001110110011;
ROM[18960] <= 32'b00000000011100010010000000100011;
ROM[18961] <= 32'b00000000010000010000000100010011;
ROM[18962] <= 32'b00000000001100010010000000100011;
ROM[18963] <= 32'b00000000010000010000000100010011;
ROM[18964] <= 32'b00000000010000010010000000100011;
ROM[18965] <= 32'b00000000010000010000000100010011;
ROM[18966] <= 32'b00000000010100010010000000100011;
ROM[18967] <= 32'b00000000010000010000000100010011;
ROM[18968] <= 32'b00000000011000010010000000100011;
ROM[18969] <= 32'b00000000010000010000000100010011;
ROM[18970] <= 32'b00000001010000000000001110010011;
ROM[18971] <= 32'b00000000100000111000001110010011;
ROM[18972] <= 32'b01000000011100010000001110110011;
ROM[18973] <= 32'b00000000011100000000001000110011;
ROM[18974] <= 32'b00000000001000000000000110110011;
ROM[18975] <= 32'b11100011010111111111000011101111;
ROM[18976] <= 32'b11111111110000010000000100010011;
ROM[18977] <= 32'b00000000000000010010001110000011;
ROM[18978] <= 32'b00000000011101100010000000100011;
ROM[18979] <= 32'b00000000010100010010000000100011;
ROM[18980] <= 32'b00000000010000010000000100010011;
ROM[18981] <= 32'b00000000010000100010001110000011;
ROM[18982] <= 32'b00000000011100010010000000100011;
ROM[18983] <= 32'b00000000010000010000000100010011;
ROM[18984] <= 32'b00000000000000011010001110000011;
ROM[18985] <= 32'b00000000011100010010000000100011;
ROM[18986] <= 32'b00000000010000010000000100010011;
ROM[18987] <= 32'b00000000101000000000001110010011;
ROM[18988] <= 32'b00000000011100010010000000100011;
ROM[18989] <= 32'b00000000010000010000000100010011;
ROM[18990] <= 32'b00000000000000010011001110110111;
ROM[18991] <= 32'b10010000010000111000001110010011;
ROM[18992] <= 32'b00000000111000111000001110110011;
ROM[18993] <= 32'b00000000011100010010000000100011;
ROM[18994] <= 32'b00000000010000010000000100010011;
ROM[18995] <= 32'b00000000001100010010000000100011;
ROM[18996] <= 32'b00000000010000010000000100010011;
ROM[18997] <= 32'b00000000010000010010000000100011;
ROM[18998] <= 32'b00000000010000010000000100010011;
ROM[18999] <= 32'b00000000010100010010000000100011;
ROM[19000] <= 32'b00000000010000010000000100010011;
ROM[19001] <= 32'b00000000011000010010000000100011;
ROM[19002] <= 32'b00000000010000010000000100010011;
ROM[19003] <= 32'b00000001010000000000001110010011;
ROM[19004] <= 32'b00000000100000111000001110010011;
ROM[19005] <= 32'b01000000011100010000001110110011;
ROM[19006] <= 32'b00000000011100000000001000110011;
ROM[19007] <= 32'b00000000001000000000000110110011;
ROM[19008] <= 32'b11111101010011110110000011101111;
ROM[19009] <= 32'b11111111110000010000000100010011;
ROM[19010] <= 32'b00000000000000010010001110000011;
ROM[19011] <= 32'b11111111110000010000000100010011;
ROM[19012] <= 32'b00000000000000010010010000000011;
ROM[19013] <= 32'b01000000011101000000001110110011;
ROM[19014] <= 32'b00000000011100010010000000100011;
ROM[19015] <= 32'b00000000010000010000000100010011;
ROM[19016] <= 32'b00000000000000010011001110110111;
ROM[19017] <= 32'b10010110110000111000001110010011;
ROM[19018] <= 32'b00000000111000111000001110110011;
ROM[19019] <= 32'b00000000011100010010000000100011;
ROM[19020] <= 32'b00000000010000010000000100010011;
ROM[19021] <= 32'b00000000001100010010000000100011;
ROM[19022] <= 32'b00000000010000010000000100010011;
ROM[19023] <= 32'b00000000010000010010000000100011;
ROM[19024] <= 32'b00000000010000010000000100010011;
ROM[19025] <= 32'b00000000010100010010000000100011;
ROM[19026] <= 32'b00000000010000010000000100010011;
ROM[19027] <= 32'b00000000011000010010000000100011;
ROM[19028] <= 32'b00000000010000010000000100010011;
ROM[19029] <= 32'b00000001010000000000001110010011;
ROM[19030] <= 32'b00000000010000111000001110010011;
ROM[19031] <= 32'b01000000011100010000001110110011;
ROM[19032] <= 32'b00000000011100000000001000110011;
ROM[19033] <= 32'b00000000001000000000000110110011;
ROM[19034] <= 32'b10101100000111111111000011101111;
ROM[19035] <= 32'b00000000000000010011001110110111;
ROM[19036] <= 32'b10011011100000111000001110010011;
ROM[19037] <= 32'b00000000111000111000001110110011;
ROM[19038] <= 32'b00000000011100010010000000100011;
ROM[19039] <= 32'b00000000010000010000000100010011;
ROM[19040] <= 32'b00000000001100010010000000100011;
ROM[19041] <= 32'b00000000010000010000000100010011;
ROM[19042] <= 32'b00000000010000010010000000100011;
ROM[19043] <= 32'b00000000010000010000000100010011;
ROM[19044] <= 32'b00000000010100010010000000100011;
ROM[19045] <= 32'b00000000010000010000000100010011;
ROM[19046] <= 32'b00000000011000010010000000100011;
ROM[19047] <= 32'b00000000010000010000000100010011;
ROM[19048] <= 32'b00000001010000000000001110010011;
ROM[19049] <= 32'b00000000100000111000001110010011;
ROM[19050] <= 32'b01000000011100010000001110110011;
ROM[19051] <= 32'b00000000011100000000001000110011;
ROM[19052] <= 32'b00000000001000000000000110110011;
ROM[19053] <= 32'b10110000100011111111000011101111;
ROM[19054] <= 32'b11111111110000010000000100010011;
ROM[19055] <= 32'b00000000000000010010001110000011;
ROM[19056] <= 32'b00000000011101100010000000100011;
ROM[19057] <= 32'b00000000000000000000001110010011;
ROM[19058] <= 32'b00000000011100010010000000100011;
ROM[19059] <= 32'b00000000010000010000000100010011;
ROM[19060] <= 32'b00000001010000000000001110010011;
ROM[19061] <= 32'b01000000011100011000001110110011;
ROM[19062] <= 32'b00000000000000111010000010000011;
ROM[19063] <= 32'b11111111110000010000000100010011;
ROM[19064] <= 32'b00000000000000010010001110000011;
ROM[19065] <= 32'b00000000011100100010000000100011;
ROM[19066] <= 32'b00000000010000100000000100010011;
ROM[19067] <= 32'b00000001010000000000001110010011;
ROM[19068] <= 32'b01000000011100011000001110110011;
ROM[19069] <= 32'b00000000010000111010000110000011;
ROM[19070] <= 32'b00000000100000111010001000000011;
ROM[19071] <= 32'b00000000110000111010001010000011;
ROM[19072] <= 32'b00000001000000111010001100000011;
ROM[19073] <= 32'b00000000000000001000000011100111;
ROM[19074] <= 32'b00000000110100000000001110010011;
ROM[19075] <= 32'b00000000011100010010000000100011;
ROM[19076] <= 32'b00000000010000010000000100010011;
ROM[19077] <= 32'b00000001010000000000001110010011;
ROM[19078] <= 32'b01000000011100011000001110110011;
ROM[19079] <= 32'b00000000000000111010000010000011;
ROM[19080] <= 32'b11111111110000010000000100010011;
ROM[19081] <= 32'b00000000000000010010001110000011;
ROM[19082] <= 32'b00000000011100100010000000100011;
ROM[19083] <= 32'b00000000010000100000000100010011;
ROM[19084] <= 32'b00000001010000000000001110010011;
ROM[19085] <= 32'b01000000011100011000001110110011;
ROM[19086] <= 32'b00000000010000111010000110000011;
ROM[19087] <= 32'b00000000100000111010001000000011;
ROM[19088] <= 32'b00000000110000111010001010000011;
ROM[19089] <= 32'b00000001000000111010001100000011;
ROM[19090] <= 32'b00000000000000001000000011100111;
ROM[19091] <= 32'b00000000100000000000001110010011;
ROM[19092] <= 32'b00000000011100010010000000100011;
ROM[19093] <= 32'b00000000010000010000000100010011;
ROM[19094] <= 32'b00000001010000000000001110010011;
ROM[19095] <= 32'b01000000011100011000001110110011;
ROM[19096] <= 32'b00000000000000111010000010000011;
ROM[19097] <= 32'b11111111110000010000000100010011;
ROM[19098] <= 32'b00000000000000010010001110000011;
ROM[19099] <= 32'b00000000011100100010000000100011;
ROM[19100] <= 32'b00000000010000100000000100010011;
ROM[19101] <= 32'b00000001010000000000001110010011;
ROM[19102] <= 32'b01000000011100011000001110110011;
ROM[19103] <= 32'b00000000010000111010000110000011;
ROM[19104] <= 32'b00000000100000111010001000000011;
ROM[19105] <= 32'b00000000110000111010001010000011;
ROM[19106] <= 32'b00000001000000111010001100000011;
ROM[19107] <= 32'b00000000000000001000000011100111;
ROM[19108] <= 32'b00000010001000000000001110010011;
ROM[19109] <= 32'b00000000011100010010000000100011;
ROM[19110] <= 32'b00000000010000010000000100010011;
ROM[19111] <= 32'b00000001010000000000001110010011;
ROM[19112] <= 32'b01000000011100011000001110110011;
ROM[19113] <= 32'b00000000000000111010000010000011;
ROM[19114] <= 32'b11111111110000010000000100010011;
ROM[19115] <= 32'b00000000000000010010001110000011;
ROM[19116] <= 32'b00000000011100100010000000100011;
ROM[19117] <= 32'b00000000010000100000000100010011;
ROM[19118] <= 32'b00000001010000000000001110010011;
ROM[19119] <= 32'b01000000011100011000001110110011;
ROM[19120] <= 32'b00000000010000111010000110000011;
ROM[19121] <= 32'b00000000100000111010001000000011;
ROM[19122] <= 32'b00000000110000111010001010000011;
ROM[19123] <= 32'b00000001000000111010001100000011;
ROM[19124] <= 32'b00000000000000001000000011100111;
ROM[19125] <= 32'b00000000000000100010001110000011;
ROM[19126] <= 32'b00000000000000111000001010010011;
ROM[19127] <= 32'b00000000110100101000010000110011;
ROM[19128] <= 32'b00000000100001000010001110000011;
ROM[19129] <= 32'b00000000011100010010000000100011;
ROM[19130] <= 32'b00000000010000010000000100010011;
ROM[19131] <= 32'b00000000000000010011001110110111;
ROM[19132] <= 32'b10110011100000111000001110010011;
ROM[19133] <= 32'b00000000111000111000001110110011;
ROM[19134] <= 32'b00000000011100010010000000100011;
ROM[19135] <= 32'b00000000010000010000000100010011;
ROM[19136] <= 32'b00000000001100010010000000100011;
ROM[19137] <= 32'b00000000010000010000000100010011;
ROM[19138] <= 32'b00000000010000010010000000100011;
ROM[19139] <= 32'b00000000010000010000000100010011;
ROM[19140] <= 32'b00000000010100010010000000100011;
ROM[19141] <= 32'b00000000010000010000000100010011;
ROM[19142] <= 32'b00000000011000010010000000100011;
ROM[19143] <= 32'b00000000010000010000000100010011;
ROM[19144] <= 32'b00000001010000000000001110010011;
ROM[19145] <= 32'b00000000010000111000001110010011;
ROM[19146] <= 32'b01000000011100010000001110110011;
ROM[19147] <= 32'b00000000011100000000001000110011;
ROM[19148] <= 32'b00000000001000000000000110110011;
ROM[19149] <= 32'b10011001110111101101000011101111;
ROM[19150] <= 32'b11111111110000010000000100010011;
ROM[19151] <= 32'b00000000000000010010001110000011;
ROM[19152] <= 32'b00000000011101100010000000100011;
ROM[19153] <= 32'b00000000000000000000001110010011;
ROM[19154] <= 32'b00000000011100010010000000100011;
ROM[19155] <= 32'b00000000010000010000000100010011;
ROM[19156] <= 32'b00000001010000000000001110010011;
ROM[19157] <= 32'b01000000011100011000001110110011;
ROM[19158] <= 32'b00000000000000111010000010000011;
ROM[19159] <= 32'b11111111110000010000000100010011;
ROM[19160] <= 32'b00000000000000010010001110000011;
ROM[19161] <= 32'b00000000011100100010000000100011;
ROM[19162] <= 32'b00000000010000100000000100010011;
ROM[19163] <= 32'b00000001010000000000001110010011;
ROM[19164] <= 32'b01000000011100011000001110110011;
ROM[19165] <= 32'b00000000010000111010000110000011;
ROM[19166] <= 32'b00000000100000111010001000000011;
ROM[19167] <= 32'b00000000110000111010001010000011;
ROM[19168] <= 32'b00000001000000111010001100000011;
ROM[19169] <= 32'b00000000000000001000000011100111;
ROM[19170] <= 32'b00000000000000010011001110110111;
ROM[19171] <= 32'b10111101010000111000001110010011;
ROM[19172] <= 32'b00000000111000111000001110110011;
ROM[19173] <= 32'b00000000011100010010000000100011;
ROM[19174] <= 32'b00000000010000010000000100010011;
ROM[19175] <= 32'b00000000001100010010000000100011;
ROM[19176] <= 32'b00000000010000010000000100010011;
ROM[19177] <= 32'b00000000010000010010000000100011;
ROM[19178] <= 32'b00000000010000010000000100010011;
ROM[19179] <= 32'b00000000010100010010000000100011;
ROM[19180] <= 32'b00000000010000010000000100010011;
ROM[19181] <= 32'b00000000011000010010000000100011;
ROM[19182] <= 32'b00000000010000010000000100010011;
ROM[19183] <= 32'b00000001010000000000001110010011;
ROM[19184] <= 32'b00000000000000111000001110010011;
ROM[19185] <= 32'b01000000011100010000001110110011;
ROM[19186] <= 32'b00000000011100000000001000110011;
ROM[19187] <= 32'b00000000001000000000000110110011;
ROM[19188] <= 32'b10110000010111110110000011101111;
ROM[19189] <= 32'b11111111110000010000000100010011;
ROM[19190] <= 32'b00000000000000010010001110000011;
ROM[19191] <= 32'b00000000011101100010000000100011;
ROM[19192] <= 32'b00000000000000010011001110110111;
ROM[19193] <= 32'b11000010110000111000001110010011;
ROM[19194] <= 32'b00000000111000111000001110110011;
ROM[19195] <= 32'b00000000011100010010000000100011;
ROM[19196] <= 32'b00000000010000010000000100010011;
ROM[19197] <= 32'b00000000001100010010000000100011;
ROM[19198] <= 32'b00000000010000010000000100010011;
ROM[19199] <= 32'b00000000010000010010000000100011;
ROM[19200] <= 32'b00000000010000010000000100010011;
ROM[19201] <= 32'b00000000010100010010000000100011;
ROM[19202] <= 32'b00000000010000010000000100010011;
ROM[19203] <= 32'b00000000011000010010000000100011;
ROM[19204] <= 32'b00000000010000010000000100010011;
ROM[19205] <= 32'b00000001010000000000001110010011;
ROM[19206] <= 32'b00000000000000111000001110010011;
ROM[19207] <= 32'b01000000011100010000001110110011;
ROM[19208] <= 32'b00000000011100000000001000110011;
ROM[19209] <= 32'b00000000001000000000000110110011;
ROM[19210] <= 32'b11010101010011110101000011101111;
ROM[19211] <= 32'b11111111110000010000000100010011;
ROM[19212] <= 32'b00000000000000010010001110000011;
ROM[19213] <= 32'b00000000011101100010000000100011;
ROM[19214] <= 32'b00000000000000010011001110110111;
ROM[19215] <= 32'b11001000010000111000001110010011;
ROM[19216] <= 32'b00000000111000111000001110110011;
ROM[19217] <= 32'b00000000011100010010000000100011;
ROM[19218] <= 32'b00000000010000010000000100010011;
ROM[19219] <= 32'b00000000001100010010000000100011;
ROM[19220] <= 32'b00000000010000010000000100010011;
ROM[19221] <= 32'b00000000010000010010000000100011;
ROM[19222] <= 32'b00000000010000010000000100010011;
ROM[19223] <= 32'b00000000010100010010000000100011;
ROM[19224] <= 32'b00000000010000010000000100010011;
ROM[19225] <= 32'b00000000011000010010000000100011;
ROM[19226] <= 32'b00000000010000010000000100010011;
ROM[19227] <= 32'b00000001010000000000001110010011;
ROM[19228] <= 32'b00000000000000111000001110010011;
ROM[19229] <= 32'b01000000011100010000001110110011;
ROM[19230] <= 32'b00000000011100000000001000110011;
ROM[19231] <= 32'b00000000001000000000000110110011;
ROM[19232] <= 32'b10111100000111110111000011101111;
ROM[19233] <= 32'b11111111110000010000000100010011;
ROM[19234] <= 32'b00000000000000010010001110000011;
ROM[19235] <= 32'b00000000011101100010000000100011;
ROM[19236] <= 32'b00000000000000010011001110110111;
ROM[19237] <= 32'b11001101110000111000001110010011;
ROM[19238] <= 32'b00000000111000111000001110110011;
ROM[19239] <= 32'b00000000011100010010000000100011;
ROM[19240] <= 32'b00000000010000010000000100010011;
ROM[19241] <= 32'b00000000001100010010000000100011;
ROM[19242] <= 32'b00000000010000010000000100010011;
ROM[19243] <= 32'b00000000010000010010000000100011;
ROM[19244] <= 32'b00000000010000010000000100010011;
ROM[19245] <= 32'b00000000010100010010000000100011;
ROM[19246] <= 32'b00000000010000010000000100010011;
ROM[19247] <= 32'b00000000011000010010000000100011;
ROM[19248] <= 32'b00000000010000010000000100010011;
ROM[19249] <= 32'b00000001010000000000001110010011;
ROM[19250] <= 32'b00000000000000111000001110010011;
ROM[19251] <= 32'b01000000011100010000001110110011;
ROM[19252] <= 32'b00000000011100000000001000110011;
ROM[19253] <= 32'b00000000001000000000000110110011;
ROM[19254] <= 32'b11011111110011110010000011101111;
ROM[19255] <= 32'b11111111110000010000000100010011;
ROM[19256] <= 32'b00000000000000010010001110000011;
ROM[19257] <= 32'b00000000011101100010000000100011;
ROM[19258] <= 32'b00000000000000010011001110110111;
ROM[19259] <= 32'b11010011010000111000001110010011;
ROM[19260] <= 32'b00000000111000111000001110110011;
ROM[19261] <= 32'b00000000011100010010000000100011;
ROM[19262] <= 32'b00000000010000010000000100010011;
ROM[19263] <= 32'b00000000001100010010000000100011;
ROM[19264] <= 32'b00000000010000010000000100010011;
ROM[19265] <= 32'b00000000010000010010000000100011;
ROM[19266] <= 32'b00000000010000010000000100010011;
ROM[19267] <= 32'b00000000010100010010000000100011;
ROM[19268] <= 32'b00000000010000010000000100010011;
ROM[19269] <= 32'b00000000011000010010000000100011;
ROM[19270] <= 32'b00000000010000010000000100010011;
ROM[19271] <= 32'b00000001010000000000001110010011;
ROM[19272] <= 32'b00000000000000111000001110010011;
ROM[19273] <= 32'b01000000011100010000001110110011;
ROM[19274] <= 32'b00000000011100000000001000110011;
ROM[19275] <= 32'b00000000001000000000000110110011;
ROM[19276] <= 32'b11111011110111110010000011101111;
ROM[19277] <= 32'b11111111110000010000000100010011;
ROM[19278] <= 32'b00000000000000010010001110000011;
ROM[19279] <= 32'b00000000011101100010000000100011;
ROM[19280] <= 32'b00000000000000010011001110110111;
ROM[19281] <= 32'b11011000110000111000001110010011;
ROM[19282] <= 32'b00000000111000111000001110110011;
ROM[19283] <= 32'b00000000011100010010000000100011;
ROM[19284] <= 32'b00000000010000010000000100010011;
ROM[19285] <= 32'b00000000001100010010000000100011;
ROM[19286] <= 32'b00000000010000010000000100010011;
ROM[19287] <= 32'b00000000010000010010000000100011;
ROM[19288] <= 32'b00000000010000010000000100010011;
ROM[19289] <= 32'b00000000010100010010000000100011;
ROM[19290] <= 32'b00000000010000010000000100010011;
ROM[19291] <= 32'b00000000011000010010000000100011;
ROM[19292] <= 32'b00000000010000010000000100010011;
ROM[19293] <= 32'b00000001010000000000001110010011;
ROM[19294] <= 32'b00000000000000111000001110010011;
ROM[19295] <= 32'b01000000011100010000001110110011;
ROM[19296] <= 32'b00000000011100000000001000110011;
ROM[19297] <= 32'b00000000001000000000000110110011;
ROM[19298] <= 32'b00000101010000000000000011101111;
ROM[19299] <= 32'b11111111110000010000000100010011;
ROM[19300] <= 32'b00000000000000010010001110000011;
ROM[19301] <= 32'b00000000011101100010000000100011;
ROM[19302] <= 32'b00000000000000000000001110010011;
ROM[19303] <= 32'b00000000011100010010000000100011;
ROM[19304] <= 32'b00000000010000010000000100010011;
ROM[19305] <= 32'b00000001010000000000001110010011;
ROM[19306] <= 32'b01000000011100011000001110110011;
ROM[19307] <= 32'b00000000000000111010000010000011;
ROM[19308] <= 32'b11111111110000010000000100010011;
ROM[19309] <= 32'b00000000000000010010001110000011;
ROM[19310] <= 32'b00000000011100100010000000100011;
ROM[19311] <= 32'b00000000010000100000000100010011;
ROM[19312] <= 32'b00000001010000000000001110010011;
ROM[19313] <= 32'b01000000011100011000001110110011;
ROM[19314] <= 32'b00000000010000111010000110000011;
ROM[19315] <= 32'b00000000100000111010001000000011;
ROM[19316] <= 32'b00000000110000111010001010000011;
ROM[19317] <= 32'b00000001000000111010001100000011;
ROM[19318] <= 32'b00000000000000001000000011100111;
ROM[19319] <= 32'b00000000000000000000001110010011;
ROM[19320] <= 32'b01000000011100000000001110110011;
ROM[19321] <= 32'b00000000000100111000001110010011;
ROM[19322] <= 32'b01000000011100000000001110110011;
ROM[19323] <= 32'b00000000000100111000001110010011;
ROM[19324] <= 32'b00000000000000111000101001100011;
ROM[19325] <= 32'b00000000000000010011001110110111;
ROM[19326] <= 32'b11100000100000111000001110010011;
ROM[19327] <= 32'b00000000111000111000001110110011;
ROM[19328] <= 32'b00000000000000111000000011100111;
ROM[19329] <= 32'b11111101100111111111000011101111;
ROM[19330] <= 32'b00000000000000000000001110010011;
ROM[19331] <= 32'b00000000011100010010000000100011;
ROM[19332] <= 32'b00000000010000010000000100010011;
ROM[19333] <= 32'b00000001010000000000001110010011;
ROM[19334] <= 32'b01000000011100011000001110110011;
ROM[19335] <= 32'b00000000000000111010000010000011;
ROM[19336] <= 32'b11111111110000010000000100010011;
ROM[19337] <= 32'b00000000000000010010001110000011;
ROM[19338] <= 32'b00000000011100100010000000100011;
ROM[19339] <= 32'b00000000010000100000000100010011;
ROM[19340] <= 32'b00000001010000000000001110010011;
ROM[19341] <= 32'b01000000011100011000001110110011;
ROM[19342] <= 32'b00000000010000111010000110000011;
ROM[19343] <= 32'b00000000100000111010001000000011;
ROM[19344] <= 32'b00000000110000111010001010000011;
ROM[19345] <= 32'b00000001000000111010001100000011;
ROM[19346] <= 32'b00000000000000001000000011100111;
ROM[19347] <= 32'b00000000000000010010000000100011;
ROM[19348] <= 32'b00000000010000010000000100010011;
ROM[19349] <= 32'b00000000000000010010000000100011;
ROM[19350] <= 32'b00000000010000010000000100010011;
ROM[19351] <= 32'b00000000000000000000001110010011;
ROM[19352] <= 32'b00000000011100011010000000100011;
ROM[19353] <= 32'b00000000000000011010001110000011;
ROM[19354] <= 32'b00000000011100010010000000100011;
ROM[19355] <= 32'b00000000010000010000000100010011;
ROM[19356] <= 32'b00000000000000100010001110000011;
ROM[19357] <= 32'b11111111110000010000000100010011;
ROM[19358] <= 32'b00000000000000010010010000000011;
ROM[19359] <= 32'b00000000011101000010001110110011;
ROM[19360] <= 32'b01000000011100000000001110110011;
ROM[19361] <= 32'b00000000000100111000001110010011;
ROM[19362] <= 32'b00000000000000111000101001100011;
ROM[19363] <= 32'b00000000000000010011001110110111;
ROM[19364] <= 32'b11110010010000111000001110010011;
ROM[19365] <= 32'b00000000111000111000001110110011;
ROM[19366] <= 32'b00000000000000111000000011100111;
ROM[19367] <= 32'b00000000000000000000001110010011;
ROM[19368] <= 32'b00000000011100011010001000100011;
ROM[19369] <= 32'b00000000010000011010001110000011;
ROM[19370] <= 32'b00000000011100010010000000100011;
ROM[19371] <= 32'b00000000010000010000000100010011;
ROM[19372] <= 32'b00000110010000000000001110010011;
ROM[19373] <= 32'b11111111110000010000000100010011;
ROM[19374] <= 32'b00000000000000010010010000000011;
ROM[19375] <= 32'b00000000011101000010001110110011;
ROM[19376] <= 32'b01000000011100000000001110110011;
ROM[19377] <= 32'b00000000000100111000001110010011;
ROM[19378] <= 32'b00000000000000111000101001100011;
ROM[19379] <= 32'b00000000000000010011001110110111;
ROM[19380] <= 32'b11110000000000111000001110010011;
ROM[19381] <= 32'b00000000111000111000001110110011;
ROM[19382] <= 32'b00000000000000111000000011100111;
ROM[19383] <= 32'b00000000010000011010001110000011;
ROM[19384] <= 32'b00000000011100010010000000100011;
ROM[19385] <= 32'b00000000010000010000000100010011;
ROM[19386] <= 32'b00000000000100000000001110010011;
ROM[19387] <= 32'b11111111110000010000000100010011;
ROM[19388] <= 32'b00000000000000010010010000000011;
ROM[19389] <= 32'b00000000011101000000001110110011;
ROM[19390] <= 32'b00000000011100011010001000100011;
ROM[19391] <= 32'b11111010100111111111000011101111;
ROM[19392] <= 32'b00000000000000011010001110000011;
ROM[19393] <= 32'b00000000011100010010000000100011;
ROM[19394] <= 32'b00000000010000010000000100010011;
ROM[19395] <= 32'b00000000000100000000001110010011;
ROM[19396] <= 32'b11111111110000010000000100010011;
ROM[19397] <= 32'b00000000000000010010010000000011;
ROM[19398] <= 32'b00000000011101000000001110110011;
ROM[19399] <= 32'b00000000011100011010000000100011;
ROM[19400] <= 32'b11110100010111111111000011101111;
ROM[19401] <= 32'b00000000000000000000001110010011;
ROM[19402] <= 32'b00000000011100010010000000100011;
ROM[19403] <= 32'b00000000010000010000000100010011;
ROM[19404] <= 32'b00000001010000000000001110010011;
ROM[19405] <= 32'b01000000011100011000001110110011;
ROM[19406] <= 32'b00000000000000111010000010000011;
ROM[19407] <= 32'b11111111110000010000000100010011;
ROM[19408] <= 32'b00000000000000010010001110000011;
ROM[19409] <= 32'b00000000011100100010000000100011;
ROM[19410] <= 32'b00000000010000100000000100010011;
ROM[19411] <= 32'b00000001010000000000001110010011;
ROM[19412] <= 32'b01000000011100011000001110110011;
ROM[19413] <= 32'b00000000010000111010000110000011;
ROM[19414] <= 32'b00000000100000111010001000000011;
ROM[19415] <= 32'b00000000110000111010001010000011;
ROM[19416] <= 32'b00000001000000111010001100000011;
ROM[19417] <= 32'b00000000000000001000000011100111;
ROM[19418] <= 32'b00000000000000111000000010010011;
        end
    assign address = addr[16:2];
    assign Inst = ROM[address];
        
endmodule