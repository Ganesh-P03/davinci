module ROM (                    //Instruction Memory
    input [16:0] addr,
    input clock,
    output [31:0] Inst
    );
    wire [14:0] address;
    
    (* ram_style="block" *)
    reg [31:0] ROM[32767:0];

    initial
        begin
ROM[0] <= 32'b00000000000000000010011100110111;
ROM[1] <= 32'b01011000000001110000011100010011;
ROM[2] <= 32'b00000000000000100010011010110111;
ROM[3] <= 32'b01011000000001101000011010010011;
ROM[4] <= 32'b00000100000001101010000000100011;
ROM[5] <= 32'b00000100000001101010001000100011;
ROM[6] <= 32'b00000100000001101010010000100011;
ROM[7] <= 32'b00000100000001101010011000100011;
ROM[8] <= 32'b00000100000001101010100000100011;
ROM[9] <= 32'b00000100000001101010101000100011;
ROM[10] <= 32'b00000100000001101010110000100011;
ROM[11] <= 32'b00000100000001101010111000100011;
ROM[12] <= 32'b00000110000001101010000000100011;
ROM[13] <= 32'b00000110000001101010001000100011;
ROM[14] <= 32'b00000110000001101010010000100011;
ROM[15] <= 32'b00000110000001101010011000100011;
ROM[16] <= 32'b00000110000001101010100000100011;
ROM[17] <= 32'b00000110000001101010101000100011;
ROM[18] <= 32'b00000110000001101010110000100011;
ROM[19] <= 32'b00000110000001101010111000100011;
ROM[20] <= 32'b00001000000001101010000000100011;
ROM[21] <= 32'b00001000000001101010001000100011;
ROM[22] <= 32'b00001000000001101010010000100011;
ROM[23] <= 32'b00001000000001101010011000100011;
ROM[24] <= 32'b00001000000001101010100000100011;
ROM[25] <= 32'b00001000000001101010101000100011;
ROM[26] <= 32'b00001000000001101010110000100011;
ROM[27] <= 32'b00001000000001101010111000100011;
ROM[28] <= 32'b00001010000001101010000000100011;
ROM[29] <= 32'b00001010000001101010001000100011;
ROM[30] <= 32'b00001010000001101010010000100011;
ROM[31] <= 32'b00001010000001101010011000100011;
ROM[32] <= 32'b00001010000001101010100000100011;
ROM[33] <= 32'b00001010000001101010101000100011;
ROM[34] <= 32'b00001010000001101010110000100011;
ROM[35] <= 32'b00001010000001101010111000100011;
ROM[36] <= 32'b00001100000001101010000000100011;
ROM[37] <= 32'b00001100000001101010001000100011;
ROM[38] <= 32'b00001100000001101010010000100011;
ROM[39] <= 32'b00001100000001101010011000100011;
ROM[40] <= 32'b00001100000001101010100000100011;
ROM[41] <= 32'b00001100000001101010101000100011;
ROM[42] <= 32'b00001100000001101010110000100011;
ROM[43] <= 32'b00001100000001101010111000100011;
ROM[44] <= 32'b00001110000001101010000000100011;
ROM[45] <= 32'b00001110000001101010001000100011;
ROM[46] <= 32'b00001110000001101010010000100011;
ROM[47] <= 32'b00001110000001101010011000100011;
ROM[48] <= 32'b00001110000001101010100000100011;
ROM[49] <= 32'b00001110000001101010101000100011;
ROM[50] <= 32'b00001110000001101010110000100011;
ROM[51] <= 32'b00001110000001101010111000100011;
ROM[52] <= 32'b00010000000001101010000000100011;
ROM[53] <= 32'b00010000000001101010001000100011;
ROM[54] <= 32'b00010000000001101010010000100011;
ROM[55] <= 32'b00010000000001101010011000100011;
ROM[56] <= 32'b00010000000001101010100000100011;
ROM[57] <= 32'b00010000000001101010101000100011;
ROM[58] <= 32'b00010000000001101010110000100011;
ROM[59] <= 32'b00010000000001101010111000100011;
ROM[60] <= 32'b00010010000001101010000000100011;
ROM[61] <= 32'b00010010000001101010001000100011;
ROM[62] <= 32'b00010010000001101010010000100011;
ROM[63] <= 32'b00010010000001101010011000100011;
ROM[64] <= 32'b00010010000001101010100000100011;
ROM[65] <= 32'b00010010000001101010101000100011;
ROM[66] <= 32'b00010010000001101010110000100011;
ROM[67] <= 32'b00010010000001101010111000100011;
ROM[68] <= 32'b00010100000001101010000000100011;
ROM[69] <= 32'b00010100000001101010001000100011;
ROM[70] <= 32'b00010100000001101010010000100011;
ROM[71] <= 32'b00010100000001101010011000100011;
ROM[72] <= 32'b00010100000001101010100000100011;
ROM[73] <= 32'b00010100000001101010101000100011;
ROM[74] <= 32'b00010100000001101010110000100011;
ROM[75] <= 32'b00010100000001101010111000100011;
ROM[76] <= 32'b00010110000001101010000000100011;
ROM[77] <= 32'b00010110000001101010001000100011;
ROM[78] <= 32'b00010110000001101010010000100011;
ROM[79] <= 32'b00010110000001101010011000100011;
ROM[80] <= 32'b00010110000001101010100000100011;
ROM[81] <= 32'b00010110000001101010101000100011;
ROM[82] <= 32'b00010110000001101010110000100011;
ROM[83] <= 32'b00010110000001101010111000100011;
ROM[84] <= 32'b00011000000001101010000000100011;
ROM[85] <= 32'b00011000000001101010001000100011;
ROM[86] <= 32'b00011000000001101010010000100011;
ROM[87] <= 32'b00011000000001101010011000100011;
ROM[88] <= 32'b00011000000001101010100000100011;
ROM[89] <= 32'b00011000000001101010101000100011;
ROM[90] <= 32'b00011000000001101010110000100011;
ROM[91] <= 32'b00011000000001101010111000100011;
ROM[92] <= 32'b00011010000001101010000000100011;
ROM[93] <= 32'b00011010000001101010001000100011;
ROM[94] <= 32'b00011010000001101010010000100011;
ROM[95] <= 32'b00011010000001101010011000100011;
ROM[96] <= 32'b00011010000001101010100000100011;
ROM[97] <= 32'b00011010000001101010101000100011;
ROM[98] <= 32'b00011010000001101010110000100011;
ROM[99] <= 32'b00011010000001101010111000100011;
ROM[100] <= 32'b00011100000001101010000000100011;
ROM[101] <= 32'b00011100000001101010001000100011;
ROM[102] <= 32'b00011100000001101010010000100011;
ROM[103] <= 32'b00011100000001101010011000100011;
ROM[104] <= 32'b00011100000001101010100000100011;
ROM[105] <= 32'b00011100000001101010101000100011;
ROM[106] <= 32'b00011100000001101010110000100011;
ROM[107] <= 32'b00011100000001101010111000100011;
ROM[108] <= 32'b00011110000001101010000000100011;
ROM[109] <= 32'b00011110000001101010001000100011;
ROM[110] <= 32'b00011110000001101010010000100011;
ROM[111] <= 32'b00011110000001101010011000100011;
ROM[112] <= 32'b00011110000001101010100000100011;
ROM[113] <= 32'b00011110000001101010101000100011;
ROM[114] <= 32'b00011110000001101010110000100011;
ROM[115] <= 32'b00011110000001101010111000100011;
ROM[116] <= 32'b00100000000001101010000000100011;
ROM[117] <= 32'b00100000000001101010001000100011;
ROM[118] <= 32'b00100000000001101010010000100011;
ROM[119] <= 32'b00100000000001101010011000100011;
ROM[120] <= 32'b00100000000001101010100000100011;
ROM[121] <= 32'b00100000000001101010101000100011;
ROM[122] <= 32'b00100000000001101010110000100011;
ROM[123] <= 32'b00100000000001101010111000100011;
ROM[124] <= 32'b00100010000001101010000000100011;
ROM[125] <= 32'b00100010000001101010001000100011;
ROM[126] <= 32'b00100010000001101010010000100011;
ROM[127] <= 32'b00100010000001101010011000100011;
ROM[128] <= 32'b00100010000001101010100000100011;
ROM[129] <= 32'b00100010000001101010101000100011;
ROM[130] <= 32'b00100010000001101010110000100011;
ROM[131] <= 32'b00100010000001101010111000100011;
ROM[132] <= 32'b00100100000001101010000000100011;
ROM[133] <= 32'b00100100000001101010001000100011;
ROM[134] <= 32'b00100100000001101010010000100011;
ROM[135] <= 32'b00100100000001101010011000100011;
ROM[136] <= 32'b00100100000001101010100000100011;
ROM[137] <= 32'b00100100000001101010101000100011;
ROM[138] <= 32'b00100100000001101010110000100011;
ROM[139] <= 32'b00100100000001101010111000100011;
ROM[140] <= 32'b00100110000001101010000000100011;
ROM[141] <= 32'b00100110000001101010001000100011;
ROM[142] <= 32'b00100110000001101010010000100011;
ROM[143] <= 32'b00100110000001101010011000100011;
ROM[144] <= 32'b00100110000001101010100000100011;
ROM[145] <= 32'b00100110000001101010101000100011;
ROM[146] <= 32'b00100110000001101010110000100011;
ROM[147] <= 32'b00100110000001101010111000100011;
ROM[148] <= 32'b00101000000001101010000000100011;
ROM[149] <= 32'b00101000000001101010001000100011;
ROM[150] <= 32'b00101000000001101010010000100011;
ROM[151] <= 32'b00101000000001101010011000100011;
ROM[152] <= 32'b00101000000001101010100000100011;
ROM[153] <= 32'b00101000000001101010101000100011;
ROM[154] <= 32'b00101000000001101010110000100011;
ROM[155] <= 32'b00101000000001101010111000100011;
ROM[156] <= 32'b00101010000001101010000000100011;
ROM[157] <= 32'b00101010000001101010001000100011;
ROM[158] <= 32'b00101010000001101010010000100011;
ROM[159] <= 32'b00101010000001101010011000100011;
ROM[160] <= 32'b00101010000001101010100000100011;
ROM[161] <= 32'b00101010000001101010101000100011;
ROM[162] <= 32'b00101010000001101010110000100011;
ROM[163] <= 32'b00101010000001101010111000100011;
ROM[164] <= 32'b00101100000001101010000000100011;
ROM[165] <= 32'b00101100000001101010001000100011;
ROM[166] <= 32'b00101100000001101010010000100011;
ROM[167] <= 32'b00101100000001101010011000100011;
ROM[168] <= 32'b00101100000001101010100000100011;
ROM[169] <= 32'b00101100000001101010101000100011;
ROM[170] <= 32'b00101100000001101010110000100011;
ROM[171] <= 32'b00101100000001101010111000100011;
ROM[172] <= 32'b00101110000001101010000000100011;
ROM[173] <= 32'b00101110000001101010001000100011;
ROM[174] <= 32'b00101110000001101010010000100011;
ROM[175] <= 32'b00101110000001101010011000100011;
ROM[176] <= 32'b00101110000001101010100000100011;
ROM[177] <= 32'b00101110000001101010101000100011;
ROM[178] <= 32'b00101110000001101010110000100011;
ROM[179] <= 32'b00101110000001101010111000100011;
ROM[180] <= 32'b00110000000001101010000000100011;
ROM[181] <= 32'b00110000000001101010001000100011;
ROM[182] <= 32'b00110000000001101010010000100011;
ROM[183] <= 32'b00110000000001101010011000100011;
ROM[184] <= 32'b00110000000001101010100000100011;
ROM[185] <= 32'b00110000000001101010101000100011;
ROM[186] <= 32'b00110000000001101010110000100011;
ROM[187] <= 32'b00110000000001101010111000100011;
ROM[188] <= 32'b00110010000001101010000000100011;
ROM[189] <= 32'b00110010000001101010001000100011;
ROM[190] <= 32'b00110010000001101010010000100011;
ROM[191] <= 32'b00110010000001101010011000100011;
ROM[192] <= 32'b00110010000001101010100000100011;
ROM[193] <= 32'b00110010000001101010101000100011;
ROM[194] <= 32'b00110010000001101010110000100011;
ROM[195] <= 32'b00110010000001101010111000100011;
ROM[196] <= 32'b00110100000001101010000000100011;
ROM[197] <= 32'b00110100000001101010001000100011;
ROM[198] <= 32'b00110100000001101010010000100011;
ROM[199] <= 32'b00110100000001101010011000100011;
ROM[200] <= 32'b00110100000001101010100000100011;
ROM[201] <= 32'b00110100000001101010101000100011;
ROM[202] <= 32'b00110100000001101010110000100011;
ROM[203] <= 32'b00110100000001101010111000100011;
ROM[204] <= 32'b00110110000001101010000000100011;
ROM[205] <= 32'b00110110000001101010001000100011;
ROM[206] <= 32'b00110110000001101010010000100011;
ROM[207] <= 32'b00110110000001101010011000100011;
ROM[208] <= 32'b00110110000001101010100000100011;
ROM[209] <= 32'b00110110000001101010101000100011;
ROM[210] <= 32'b00110110000001101010110000100011;
ROM[211] <= 32'b00110110000001101010111000100011;
ROM[212] <= 32'b00111000000001101010000000100011;
ROM[213] <= 32'b00111000000001101010001000100011;
ROM[214] <= 32'b00111000000001101010010000100011;
ROM[215] <= 32'b00111000000001101010011000100011;
ROM[216] <= 32'b00111000000001101010100000100011;
ROM[217] <= 32'b00111000000001101010101000100011;
ROM[218] <= 32'b00111000000001101010110000100011;
ROM[219] <= 32'b00111000000001101010111000100011;
ROM[220] <= 32'b00111010000001101010000000100011;
ROM[221] <= 32'b00111010000001101010001000100011;
ROM[222] <= 32'b00111010000001101010010000100011;
ROM[223] <= 32'b00111010000001101010011000100011;
ROM[224] <= 32'b00111010000001101010100000100011;
ROM[225] <= 32'b00111010000001101010101000100011;
ROM[226] <= 32'b00111010000001101010110000100011;
ROM[227] <= 32'b00111010000001101010111000100011;
ROM[228] <= 32'b00111100000001101010000000100011;
ROM[229] <= 32'b00111100000001101010001000100011;
ROM[230] <= 32'b00111100000001101010010000100011;
ROM[231] <= 32'b00111100000001101010011000100011;
ROM[232] <= 32'b00111100000001101010100000100011;
ROM[233] <= 32'b00111100000001101010101000100011;
ROM[234] <= 32'b00111100000001101010110000100011;
ROM[235] <= 32'b00111100000001101010111000100011;
ROM[236] <= 32'b00111110000001101010000000100011;
ROM[237] <= 32'b00111110000001101010001000100011;
ROM[238] <= 32'b00111110000001101010010000100011;
ROM[239] <= 32'b00111110000001101010011000100011;
ROM[240] <= 32'b00111110000001101010100000100011;
ROM[241] <= 32'b00111110000001101010101000100011;
ROM[242] <= 32'b00111110000001101010110000100011;
ROM[243] <= 32'b00111110000001101010111000100011;
ROM[244] <= 32'b00000000000001101000011000010011;
ROM[245] <= 32'b01000000000001101000000100010011;
ROM[246] <= 32'b00000000000000010000000110010011;
ROM[247] <= 32'b00000000000000010000001000010011;
ROM[248] <= 32'b00000000000000010000001010010011;
ROM[249] <= 32'b00000000000000010000001100010011;
ROM[250] <= 32'b00000000000000000000001110110111;
ROM[251] <= 32'b01000011010000111000001110010011;
ROM[252] <= 32'b00000000111000111000001110110011;
ROM[253] <= 32'b00000000011100010010000000100011;
ROM[254] <= 32'b00000000010000010000000100010011;
ROM[255] <= 32'b00000000001100010010000000100011;
ROM[256] <= 32'b00000000010000010000000100010011;
ROM[257] <= 32'b00000000010000010010000000100011;
ROM[258] <= 32'b00000000010000010000000100010011;
ROM[259] <= 32'b00000000010100010010000000100011;
ROM[260] <= 32'b00000000010000010000000100010011;
ROM[261] <= 32'b00000000011000010010000000100011;
ROM[262] <= 32'b00000000010000010000000100010011;
ROM[263] <= 32'b00000001010000000000001110010011;
ROM[264] <= 32'b00000000000000111000001110010011;
ROM[265] <= 32'b01000000011100010000001110110011;
ROM[266] <= 32'b00000000011100000000001000110011;
ROM[267] <= 32'b00000000001000000000000110110011;
ROM[268] <= 32'b00110001000000000000000011101111;
ROM[269] <= 32'b11111111110000010000000100010011;
ROM[270] <= 32'b00000000000000010010001110000011;
ROM[271] <= 32'b00111000100000000000000011101111;
ROM[272] <= 32'b00000000101000000000001110010011;
ROM[273] <= 32'b00000000011100010010000000100011;
ROM[274] <= 32'b00000000010000010000000100010011;
ROM[275] <= 32'b00000000000000000000001110110111;
ROM[276] <= 32'b01001001100000111000001110010011;
ROM[277] <= 32'b00000000111000111000001110110011;
ROM[278] <= 32'b00000000011100010010000000100011;
ROM[279] <= 32'b00000000010000010000000100010011;
ROM[280] <= 32'b00000000001100010010000000100011;
ROM[281] <= 32'b00000000010000010000000100010011;
ROM[282] <= 32'b00000000010000010010000000100011;
ROM[283] <= 32'b00000000010000010000000100010011;
ROM[284] <= 32'b00000000010100010010000000100011;
ROM[285] <= 32'b00000000010000010000000100010011;
ROM[286] <= 32'b00000000011000010010000000100011;
ROM[287] <= 32'b00000000010000010000000100010011;
ROM[288] <= 32'b00000001010000000000001110010011;
ROM[289] <= 32'b00000000010000111000001110010011;
ROM[290] <= 32'b01000000011100010000001110110011;
ROM[291] <= 32'b00000000011100000000001000110011;
ROM[292] <= 32'b00000000001000000000000110110011;
ROM[293] <= 32'b00000011110000000000000011101111;
ROM[294] <= 32'b00000001010000000000001110010011;
ROM[295] <= 32'b01000000011100011000001110110011;
ROM[296] <= 32'b00000000000000111010000010000011;
ROM[297] <= 32'b11111111110000010000000100010011;
ROM[298] <= 32'b00000000000000010010001110000011;
ROM[299] <= 32'b00000000011100100010000000100011;
ROM[300] <= 32'b00000000010000100000000100010011;
ROM[301] <= 32'b00000001010000000000001110010011;
ROM[302] <= 32'b01000000011100011000001110110011;
ROM[303] <= 32'b00000000010000111010000110000011;
ROM[304] <= 32'b00000000100000111010001000000011;
ROM[305] <= 32'b00000000110000111010001010000011;
ROM[306] <= 32'b00000001000000111010001100000011;
ROM[307] <= 32'b00000000000000001000000011100111;
ROM[308] <= 32'b00000000000000010010000000100011;
ROM[309] <= 32'b00000000010000010000000100010011;
ROM[310] <= 32'b00000000000000010010000000100011;
ROM[311] <= 32'b00000000010000010000000100010011;
ROM[312] <= 32'b00000000000000010010000000100011;
ROM[313] <= 32'b00000000010000010000000100010011;
ROM[314] <= 32'b00000000000000010010000000100011;
ROM[315] <= 32'b00000000010000010000000100010011;
ROM[316] <= 32'b00000000001000000000001110010011;
ROM[317] <= 32'b00000000011100010010000000100011;
ROM[318] <= 32'b00000000010000010000000100010011;
ROM[319] <= 32'b11111111110000010000000100010011;
ROM[320] <= 32'b00000000000000010010001110000011;
ROM[321] <= 32'b00000000011100011010011000100011;
ROM[322] <= 32'b00000000000000000000001110010011;
ROM[323] <= 32'b00000000011100010010000000100011;
ROM[324] <= 32'b00000000010000010000000100010011;
ROM[325] <= 32'b11111111110000010000000100010011;
ROM[326] <= 32'b00000000000000010010001110000011;
ROM[327] <= 32'b00000000011100011010000000100011;
ROM[328] <= 32'b00000000000100000000001110010011;
ROM[329] <= 32'b00000000011100010010000000100011;
ROM[330] <= 32'b00000000010000010000000100010011;
ROM[331] <= 32'b11111111110000010000000100010011;
ROM[332] <= 32'b00000000000000010010001110000011;
ROM[333] <= 32'b00000000011100011010001000100011;
ROM[334] <= 32'b00000000000000100010001110000011;
ROM[335] <= 32'b00000000011100010010000000100011;
ROM[336] <= 32'b00000000010000010000000100010011;
ROM[337] <= 32'b00000000000100000000001110010011;
ROM[338] <= 32'b00000000011100010010000000100011;
ROM[339] <= 32'b00000000010000010000000100010011;
ROM[340] <= 32'b11111111110000010000000100010011;
ROM[341] <= 32'b00000000000000010010001110000011;
ROM[342] <= 32'b11111111110000010000000100010011;
ROM[343] <= 32'b00000000000000010010010000000011;
ROM[344] <= 32'b00000000011101000010010010110011;
ROM[345] <= 32'b00000000100000111010010100110011;
ROM[346] <= 32'b00000000101001001000001110110011;
ROM[347] <= 32'b00000000000100111000001110010011;
ROM[348] <= 32'b00000000000100111111001110010011;
ROM[349] <= 32'b00000000011100010010000000100011;
ROM[350] <= 32'b00000000010000010000000100010011;
ROM[351] <= 32'b11111111110000010000000100010011;
ROM[352] <= 32'b00000000000000010010001110000011;
ROM[353] <= 32'b00000000000000111000101001100011;
ROM[354] <= 32'b00000000000000000000001110110111;
ROM[355] <= 32'b01011001110000111000001110010011;
ROM[356] <= 32'b00000000111000111000001110110011;
ROM[357] <= 32'b00000000000000111000000011100111;
ROM[358] <= 32'b00000100100000000000000011101111;
ROM[359] <= 32'b00000000000000000000001110010011;
ROM[360] <= 32'b00000000011100010010000000100011;
ROM[361] <= 32'b00000000010000010000000100010011;
ROM[362] <= 32'b00000001010000000000001110010011;
ROM[363] <= 32'b01000000011100011000001110110011;
ROM[364] <= 32'b00000000000000111010000010000011;
ROM[365] <= 32'b11111111110000010000000100010011;
ROM[366] <= 32'b00000000000000010010001110000011;
ROM[367] <= 32'b00000000011100100010000000100011;
ROM[368] <= 32'b00000000010000100000000100010011;
ROM[369] <= 32'b00000001010000000000001110010011;
ROM[370] <= 32'b01000000011100011000001110110011;
ROM[371] <= 32'b00000000010000111010000110000011;
ROM[372] <= 32'b00000000100000111010001000000011;
ROM[373] <= 32'b00000000110000111010001010000011;
ROM[374] <= 32'b00000001000000111010001100000011;
ROM[375] <= 32'b00000000000000001000000011100111;
ROM[376] <= 32'b00000000110000011010001110000011;
ROM[377] <= 32'b00000000011100010010000000100011;
ROM[378] <= 32'b00000000010000010000000100010011;
ROM[379] <= 32'b00000000000000100010001110000011;
ROM[380] <= 32'b00000000011100010010000000100011;
ROM[381] <= 32'b00000000010000010000000100010011;
ROM[382] <= 32'b11111111110000010000000100010011;
ROM[383] <= 32'b00000000000000010010001110000011;
ROM[384] <= 32'b11111111110000010000000100010011;
ROM[385] <= 32'b00000000000000010010010000000011;
ROM[386] <= 32'b00000000011101000010001110110011;
ROM[387] <= 32'b00000000011100010010000000100011;
ROM[388] <= 32'b00000000010000010000000100010011;
ROM[389] <= 32'b11111111110000010000000100010011;
ROM[390] <= 32'b00000000000000010010001110000011;
ROM[391] <= 32'b01000000011100000000001110110011;
ROM[392] <= 32'b00000000000100111000001110010011;
ROM[393] <= 32'b00000000011100010010000000100011;
ROM[394] <= 32'b00000000010000010000000100010011;
ROM[395] <= 32'b11111111110000010000000100010011;
ROM[396] <= 32'b00000000000000010010001110000011;
ROM[397] <= 32'b00000000000000111000101001100011;
ROM[398] <= 32'b00000000000000000000001110110111;
ROM[399] <= 32'b01101111110000111000001110010011;
ROM[400] <= 32'b00000000111000111000001110110011;
ROM[401] <= 32'b00000000000000111000000011100111;
ROM[402] <= 32'b00000000000000011010001110000011;
ROM[403] <= 32'b00000000011100010010000000100011;
ROM[404] <= 32'b00000000010000010000000100010011;
ROM[405] <= 32'b00000000010000011010001110000011;
ROM[406] <= 32'b00000000011100010010000000100011;
ROM[407] <= 32'b00000000010000010000000100010011;
ROM[408] <= 32'b11111111110000010000000100010011;
ROM[409] <= 32'b00000000000000010010001110000011;
ROM[410] <= 32'b11111111110000010000000100010011;
ROM[411] <= 32'b00000000000000010010010000000011;
ROM[412] <= 32'b00000000011101000000001110110011;
ROM[413] <= 32'b00000000011100010010000000100011;
ROM[414] <= 32'b00000000010000010000000100010011;
ROM[415] <= 32'b11111111110000010000000100010011;
ROM[416] <= 32'b00000000000000010010001110000011;
ROM[417] <= 32'b00000000011100011010010000100011;
ROM[418] <= 32'b00000000010000011010001110000011;
ROM[419] <= 32'b00000000011100010010000000100011;
ROM[420] <= 32'b00000000010000010000000100010011;
ROM[421] <= 32'b11111111110000010000000100010011;
ROM[422] <= 32'b00000000000000010010001110000011;
ROM[423] <= 32'b00000000011100011010000000100011;
ROM[424] <= 32'b00000000100000011010001110000011;
ROM[425] <= 32'b00000000011100010010000000100011;
ROM[426] <= 32'b00000000010000010000000100010011;
ROM[427] <= 32'b11111111110000010000000100010011;
ROM[428] <= 32'b00000000000000010010001110000011;
ROM[429] <= 32'b00000000011100011010001000100011;
ROM[430] <= 32'b00000000110000011010001110000011;
ROM[431] <= 32'b00000000011100010010000000100011;
ROM[432] <= 32'b00000000010000010000000100010011;
ROM[433] <= 32'b00000000000100000000001110010011;
ROM[434] <= 32'b00000000011100010010000000100011;
ROM[435] <= 32'b00000000010000010000000100010011;
ROM[436] <= 32'b11111111110000010000000100010011;
ROM[437] <= 32'b00000000000000010010001110000011;
ROM[438] <= 32'b11111111110000010000000100010011;
ROM[439] <= 32'b00000000000000010010010000000011;
ROM[440] <= 32'b00000000011101000000001110110011;
ROM[441] <= 32'b00000000011100010010000000100011;
ROM[442] <= 32'b00000000010000010000000100010011;
ROM[443] <= 32'b11111111110000010000000100010011;
ROM[444] <= 32'b00000000000000010010001110000011;
ROM[445] <= 32'b00000000011100011010011000100011;
ROM[446] <= 32'b11101110100111111111000011101111;
ROM[447] <= 32'b00000000010000011010001110000011;
ROM[448] <= 32'b00000000011100010010000000100011;
ROM[449] <= 32'b00000000010000010000000100010011;
ROM[450] <= 32'b00000001010000000000001110010011;
ROM[451] <= 32'b01000000011100011000001110110011;
ROM[452] <= 32'b00000000000000111010000010000011;
ROM[453] <= 32'b11111111110000010000000100010011;
ROM[454] <= 32'b00000000000000010010001110000011;
ROM[455] <= 32'b00000000011100100010000000100011;
ROM[456] <= 32'b00000000010000100000000100010011;
ROM[457] <= 32'b00000001010000000000001110010011;
ROM[458] <= 32'b01000000011100011000001110110011;
ROM[459] <= 32'b00000000010000111010000110000011;
ROM[460] <= 32'b00000000100000111010001000000011;
ROM[461] <= 32'b00000000110000111010001010000011;
ROM[462] <= 32'b00000001000000111010001100000011;
ROM[463] <= 32'b00000000000000001000000011100111;
ROM[464] <= 32'b00000000000000000000001110110111;
ROM[465] <= 32'b01111000110000111000001110010011;
ROM[466] <= 32'b00000000111000111000001110110011;
ROM[467] <= 32'b00000000011100010010000000100011;
ROM[468] <= 32'b00000000010000010000000100010011;
ROM[469] <= 32'b00000000001100010010000000100011;
ROM[470] <= 32'b00000000010000010000000100010011;
ROM[471] <= 32'b00000000010000010010000000100011;
ROM[472] <= 32'b00000000010000010000000100010011;
ROM[473] <= 32'b00000000010100010010000000100011;
ROM[474] <= 32'b00000000010000010000000100010011;
ROM[475] <= 32'b00000000011000010010000000100011;
ROM[476] <= 32'b00000000010000010000000100010011;
ROM[477] <= 32'b00000001010000000000001110010011;
ROM[478] <= 32'b00000000000000111000001110010011;
ROM[479] <= 32'b01000000011100010000001110110011;
ROM[480] <= 32'b00000000011100000000001000110011;
ROM[481] <= 32'b00000000001000000000000110110011;
ROM[482] <= 32'b11001011100111111111000011101111;
ROM[483] <= 32'b00000001010000000000001110010011;
ROM[484] <= 32'b01000000011100011000001110110011;
ROM[485] <= 32'b00000000000000111010000010000011;
ROM[486] <= 32'b11111111110000010000000100010011;
ROM[487] <= 32'b00000000000000010010001110000011;
ROM[488] <= 32'b00000000011100100010000000100011;
ROM[489] <= 32'b00000000010000100000000100010011;
ROM[490] <= 32'b00000001010000000000001110010011;
ROM[491] <= 32'b01000000011100011000001110110011;
ROM[492] <= 32'b00000000010000111010000110000011;
ROM[493] <= 32'b00000000100000111010001000000011;
ROM[494] <= 32'b00000000110000111010001010000011;
ROM[495] <= 32'b00000001000000111010001100000011;
ROM[496] <= 32'b00000000000000001000000011100111;


        end
    assign address = addr[16:2];
    assign Inst = ROM[address];
        
endmodule


						
						

// module ROM ( //Instruction Memory
//     input [15:0] address,
//     input clock,
//     input IRWrite,
//     output reg [31:0] IR
//     );
    
//     (* ram_style="block" *)
//     reg [31:0] ROM[16383:0];

//     initial
//         begin
//             $readmemb("os.mem", ROM, 0, 16383);
//             IR <= 32'd15;
//         end
    
//     always @(posedge clock)
//         begin
//             if( IRWrite )
//                 IR <= ROM[address];
//         end
        
// endmodule

						
						


						
						
